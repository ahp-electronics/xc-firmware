---------------------------------------------------------------------- 
@E-
-R8vFkRDC:FR8IMMO0Ps3E
8R
R--wOkM0MHF:FR8IOMRF0kMClsRFD8kCCRoMNCs0RFs
-
-R-

-CRtMHCsO
#R
R--I0H8ERR-MLklCFsRVFROkCM0sHRL0
#R
R--sCC#00bNRs-RC0#CR0bN0MCsRsVFROCNEHRL0
R
-#-R0D8_FOoH_OPC05FsI0H8EFR8IFM0R,j2RoC33jR"j"jjR-

-MR uNFDRb-RFsDNHR0$F VRhHRbM
R
-j-RR0NOHRPCDRFI
-
-RN4ROP0HCHREo
ER
R--.FRMRR h5FODON	RD$IN#MRCNCLD8
2R
R--BuDsFRDN-FRbDHNs0F$RV R)1R abRHM
-
-RNjROP0HCFRDI
R
-4-RR0NOHRPCEEHoR-

-RR.M)FR a1 RF5MR#sCCb0RHRM2
-
-Rup8FRDN-FRbDHNs0F$RVmRpqb7RH
MR
R--jORN0CHPRIDFR-

-RR4NHO0PECRHRoE
-
-RM.RFmRpq57RNNDI$O#RF0kMH2MoR-

-DRB	o 8CRR-NHO0PCCR8RoCFBVRp
iR
R--jNRVDMDHo8RCo
CR
R--4HRs#oHMRoC8C
R
-z-RbI7FMs7HRO-RF0kMRs8HCHO0F
MR
R--jFROkRM08MFIR-

-RR4OMFk0bRkR-

-
R
-u-RF#s0R-

-qR7a-qRR08NNMRHb#k0RsVFRM#$OFEsM#FkRNDF8
R
-T-RRO-RF0kMCFsRkk0b0
#R
R--p7mqRC-RMDNLC$R#MsOEFkMF#FRDNI8RERCMNHO0PRC,
-
-R#CDCMRCNCLDRkOFMM0HoFR5bF0HMRNDVOkM0MHF2
R
- -RhRR-CLMNDOCRD	FORCIEMORN0CHPRb5F0MHFNVDRk0MOH2FMR-

- R)1R a-#RN$EMOsFFMks#RC0#CRb5F0MHFNVDRk0MOH2FMR-

-pRBiRR-OODF	MRHbRk0
-
-RzBmaRR-OsNs$kRF00bkR-

-QRBhRR-OsNs$MRHbRk0
-
-R7zuhRR-E8NsICHs8FR0R''jR-

--R----------------------------------------------------------R--



DsHLNRs$HCCC;kR
#HCRC3CC#_08DHFoO4_4nNc3DRD;
Ck#RsIF	C3oMObN	CNo3DND;
R

M
C0$H0RW7mhaBh)#RHRo

CsMCHIO5HE80RH:RMo0CC:sR=;R.Rs

C0#CbRN0:FROkCM0ssIF8=R:RRj;-#-R0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2
R
 FMuD:NRR0HMCsoCRR:=4-;R-,Rj4R,.NHO0PDCRFRI,EEHo,FRMM
CR
sBDuNFDRH:RMo0CC:sR=;R4RR--j,,4.ORN0CHPRIDF,HREoRE,MCFMRp

8DuFNRR:HCM0oRCs:4=R;-R-R4j,,N.ROP0HCFRDIE,RH,oERMMFC
R
B D	8RoC:MRH0CCos=R:RR4;-j-R,s4RHM#HoV,RNHDDMCoR8RoC
b
z7MFI7RHs:MRH0CCos=R:R-jR-,Rj4FROkRM08MFI,bRkR2

;
R
b0Fs5a7qqRR:H#MR0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2
;R
:TRR0FkR8#0_oDFHPO_CFO0sH5I8-0E4FR8IFM0R;j2Rp

mRq7:MRHR8#0_oDFHRO;
h
 RH:RM0R#8F_Do;HOR)

 a1 :MRHR8#0_oDFHRO;
p
BiRR:H#MR0D8_FOoH;
R
BamzRF:Rk#0R0D8_FOoH;
R
BRQh:MRHR8#0_oDFHRO;
u
z7:hRRRHM#_08DHFoO
R
2
;R
8CMRW7mhaBh)
;R
ONsECH0Os0kCeRp_W7mhaBh)R_)F7VRmBWhhRa)H
#
ObFlFMMC0BRBzB_7uR
RRsbF0R5
RRRRRR7RRRRRRRRRRRRRRRRRRRRRRRRRRRRR:HRRMRRRR71a_tpmQ
B;RRRRR7R1RRRRRRRRRRRRRRRRRRRRRRRRRRRRRR:RHRMRRaR17m_pt;QB
RRRRpRRmRq7RRRRRRRRRRRRRRRRRRRRRRRRRRR:RRHMR1RRap7_mBtQ;R
RRRRRBRQhRRRRRRRRRRRRRRRRRRRRRRRRR:RRRMRHRRRR1_a7pQmtBR;
RRRRRR1jRRRRRRRRRRRRRRRRRRRRRRRRRRRR:FRRkR0RR71a_tpmQ
B;RRRRRmRBzRaRRRRRRRRRRRRRRRRRRRRRRRRRRR:RFRk0RaR17m_pt2QB;M
C8FROlMbFC;M0
F
OlMbFCRM07BwwA
)]RbRRF5s0
RRRRBRR RRRRRRRRRRRRRRRRRRRRRRRRRRRRRR:RRHMR1RRap7_mBtQ;R
RRRRR7RRRRRRRRRRRRRRRRRRRRRRRRRRRR:RRRMRHRRRR1_a7pQmtBR;
RRRRRiBpRRRRRRRRRRRRRRRRRRRRRRRRRRRR:HRRMRRRR71a_tpmQ
B;RRRRRRR)RRRRRRRRRRRRRRRRRRRRRRRRRRRRRR:RHRMRRaR17m_pt;QB
RRRRTRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR:R0FkR1RRap7_mBtQ2C;
MO8RFFlbM0CM;


ObFlFMMC0wR7w1BA]R
RRsbF0R5
RRRRRRB RRRRRRRRRRRRRRRRRRRRRRRRRRRR:HRRMRRRR71a_tpmQ
B;RRRRRRR7RRRRRRRRRRRRRRRRRRRRRRRRRRRRRR:RHRMRRaR17m_pt;QB
RRRRBRRpRiRRRRRRRRRRRRRRRRRRRRRRRRRRRR:RRHMR1RRap7_mBtQ;R
RRRRR1RRRRRRRRRRRRRRRRRRRRRRRRRRRR:RRRMRHRRRR1_a7pQmtBR;
RRRRRRTRRRRRRRRRRRRRRRRRRRRRRRRRRRRR:FRRkR0RR71a_tpmQ;B2
8CMRlOFbCFMM
0;RRRRRRRR#MHoNODRN$ssR#:R0D8_FOoH_OPC05FsR8IH04E-RI8FMR0Fj;R2
RRRRRRRRo#HMRNDTH_#oRR:#_08DHFoOC_POs0F5HRI8-0E4FR8IFM0R2jR;R
RRRRRRHR#oDMNR#1_H:oRR8#0_oDFHPO_CFO0sI5RHE80-84RF0IMFRRj2R;
RRRRR#RRHNoMDFRDo4HORRRR:0R#8D_kFOoHRR:=';4'
RRRRRRRRo#HMRNDDHFoORjRRRR:#_08koDFH:OR=jR''R;
RRRRR#RRHNoMDDRO	H_#oRRR:0R#8D_kFOoHRR:=';j'R-R-RFODOF	RVRV
RRRRR#RRHNoMDDROsH_#oRRR:0R#8D_kFOoHRR:=';j'R-R-RCODN8sRHL#ND
C8RRRRRRRR#MHoNCDRMH_#oRRRR#:R0k8_DHFoO=R:R''4;-RR-DROFRO	CLMND
C8RRRRRRRR#MHoNDDR8H_#oRRRR#:R0k8_DHFoO=R:R''j;-RR-FRDN88RHL#ND
C8RRRRRRRR#MHoNODRDC	_MH_#oRRRR#:R0k8_DHFoO=R:R''j;-RR-FRDN88RHL#ND
C8LHCoMR

RRRRRVRRNDHDH_MoO:D	RRHV5	BD C8oRj=R2CRoMNCs0RC
RRRRRRRRR	OD_o#HRR<=MRF0B;pi
RRRRRRRR8CMRMoCC0sNCR;
RRRRRsRRHM#HoD_O	H:RVBR5D8	 o=CRRR42oCCMsCN0
RRRRRRRRORRD#	_H<oR=pRBiR;
RRRRRCRRMo8RCsMCN;0C
RRRR
RRRRRRRRRRNHO0PDC_FOI_DRs:H5VRBuDsFRDN=2RjRMoCC0sNCR
RRRRRRRRRO_Ds#RHo<M=RF)0R a1 ;R
RRRRRRMRC8CRoMNCs0
C;RRRRRRRRNHO0PEC_H_oEO:DsRRHV5sBDuNFDR4=R2CRoMNCs0RC
RRRRRRRRRsOD_o#HRR<=)  1aR;
RRRRRCRRMo8RCsMCN;0C
RRRRRRRR_MFO:DsRRHV5sBDuNFDR.=R2CRoMNCs0RC
RRRRRRRRRsOD_o#HRR<=DHFoO
j;RRRRRRRRCRM8oCCMsCN0;S

S0NOH_PCD_FIDR8:H5VRpF8uD=NRRRj2oCCMsCN0
RRRRRRRRDRR8H_#o=R<R0MFRqpm7S;
SCRRMH_#o=R<R; h
RRRRRRRR8CMRMoCC0sNCR;
RRRRRNRROP0HCH_EoDE_8H:RVpR58DuFNRR=4o2RCsMCN
0CRRRRRRRRR8RD_o#HRR<=p7mq;S
SRMRC_o#HRR<= 
h;RRRRRRRRCRM8oCCMsCN0;R
RRRRRRFRM_:D8RRHV5up8FRDN=2R.RMoCC0sNCR
RRRRRRRRRD#8_H<oR=FRDojHO;S
SRMRC_o#HRR<= 
h;RRRRRRRRCRM8oCCMsCN0;S

S0NOH_PCD_FIO_D	CRM:H5VR FMuD=NRRRj2oCCMsCN0
RRRRRRRRORRDC	_MH_#o=R<R_CM#;Ho
RRRRRRRR8CMRMoCC0sNCR;
RRRRRNRROP0HCH_EoOE_DC	_MH:RV R5MDuFNRR=4o2RCsMCN
0CRRRRRRRRRDRO	M_C_o#HRR<=MRF0C#M_H
o;RRRRRRRRCRM8oCCMsCN0;R
RRRRRRFRM_	OD_:CMRRHV5u MFRDN=2R.RMoCC0sNCR
RRRRRRRRRO_D	C#M_H<oR=FRDojHO;R
RRRRRRMRC8CRoMNCs0
C;
R
RRRRRR4Rz:BRBzB_7umRu)vaRqRu51RjRRR=>R#1_Hjo52
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRmRBz=aR>ORRN$ss5,j2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRRRR=>R#T_Hjo52
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRR7R1R=RR>7RRq5aqjR2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRqpm7RRR=R>RD#8_HRo,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRBRRQRhR=R>RD#8_H;o2
S
SHoV_CRM:H5VRsCC#00bN5Rj2=jR''o2RCsMCN
0CSRRRRRRRR:z.Rw7wB]A)R)umaqRvuRR5RRRT=R>RTH_#o25j,RR
RRRSRRRRRRRRRRRRRRRRRRRRRRRRRRRRR=7R>1RR_o#H5,j2RR
RRRSRRRRRRRRRRRRRRRRRRRRRRRRRRpRBi>R=RDRO	H_#o
,RRSRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR)R=R>RO_Ds#,HoRR
RRRSRRRRRRRRRRRRRRRRRRRRRRRRRR RBR>R=RDRO	M_C_o#HR
2;SMSC8CRoMNCs0HCRVC_oM
;
SVSH_MoC4H:RVsR5C0#Cb5N0j=2RR''42CRoMNCs0SC
RRRRRRRRz:.NRw7wB]A1R)umaqRvuRR5RRRT=R>RTH_#o25j,RR
RRRSRRRRRRRRRRRRRRRRRRRRRRRRRRRRR=7R>1RR_o#H5,j2RR
RRRSRRRRRRRRRRRRRRRRRRRRRRRRRRpRBi>R=RDRO	H_#o
,RRSRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR1R=R>RO_Ds#,HoRR
RRRSRRRRRRRRRRRRRRRRRRRRRRRRRR RBR>R=RDRO	M_C_o#HR
2;SMSC8CRoMNCs0HCRVC_oM
4;
R
RRRRRR4Rp:FRVsRRHH4MRRR0FI0H8ER-4oCCMsCN0
RRRRRRRRRRRRRRRR_p4zR4:B_Bz7RBuuam)Ruvq5R1jRR=>R#1_HHo52
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRmRBzRaR=R>ROsNs$25H,RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR7=RR>TRR_o#H5,H2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR7R1R>R=RqR7aHq52
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRpRRmRq7=R>RD#8_HRo,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRhBQRR=>RsONsH$5-242;S
SS_HVoGCM:VRHRC5s#bC0NH052RR='2j'RMoCC0sNCR
RRRRRRRRRRRRRR4Rp_:z.Rw7wB]A)R)umaqRvuTR5R>R=R#T_HHo52
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR7R=1>R_o#H5,H2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRpRBi>R=R	OD_o#H,RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR)=RR>DROsH_#o
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRBR R=O>RDC	_MH_#o;R2
SSSCRM8oCCMsCN0R_HVoGCM;S
SS_HVo$CM:VRHRC5s#bC0NH052RR='24'RMoCC0sNCR
RRRRRRRRRRRRRR4Rp_:zWRw7wB]A1R)umaqRvuTR5R>R=R#T_HHo52
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR7R=1>R_o#H5,H2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRpRBi>R=R	OD_o#H,RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR1=RR>DROsH_#o
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRBR R=O>RDC	_MH_#o;R2
SSSCRM8oCCMsCN0R_HVo$CM;R

RRRRRCRRMo8RCsMCN;0C
RRRRRRRR<TR=_RT#;Ho
mSBz<aR=NROs5s$I0H8E2-4;
S
CRM8p7e_mBWhh_a))
;

