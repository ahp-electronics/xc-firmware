--
@ER--B$FbsEHo0OR52gR4g-cRRj.jd$R1MHbDO$H0ROQM
R--fN]C8:CsR#//$DMbH0OH$N/lb0DN.Uj4J4.b/blNb#Cs/DGHH/MGD/HLoCCMs/HOo_CMoCCMs.HO/lsN_bsI_Ps3E48yR-f
--

----RpB p)RXq.vdXR47-----H
DLssN$CRHC
C;kR#CHCCC38#0_oDFH4O_43ncN;DD
Ck#RCHCC03#8F_Do_HO#MHoCN83D
D;DsHLNRs$k#MHH
l;kR#Ck#MHHPl3ObFlFMMC0N#3D
D;
0CMHR0$Xv)qd4.X7#RH
bRRFRs05R
RRRRRRuR7mRRR:kRF00R#8D_kFOoH;RRRRRRRRR
RRRRRRuR1mRRR:kRF00R#8D_kFOoH;R

RRRRRqRRjRRRRH:RM0R#8D_kFOoH;R
RRRRRR4RqRRRR:MRHR8#0_FkDo;HO
RRRRRRRRRq.R:RRRRHM#_08koDFH
O;RRRRRRRRqRdRRRR:H#MR0k8_DHFoOR;
RRRRRqRRcRRRRH:RM0R#8D_kFOoH;R
RRRRRRRR7RRRR:MRHR8#0_FkDo;HO
RRRRRRRR)7uq:jRRRHM#_08koDFH
O;RRRRRRRR7qu)4RR:H#MR0k8_DHFoOR;
RRRRR7RRu.)qRH:RM0R#8D_kFOoH;R
RRRRRRuR7)Rqd:MRHR8#0_FkDo;HO
RRRRRRRR)7uq:cRRRHM#_08koDFH
O;RRRRRRRRWiBpRRR:H#MR0k8_DHFoOR;RRRRRRRR
RRRRRWRR RRRRH:RM0R#8D_kFOoH
RRRRRRR2R;R
8CMRqX)vXd.4
7;NEsOHO0C0CksRqX)vXd.4e7_RRFVXv)qd4.X7#RH
SRR#MHoNIDRCRj,I,C4Rj#F,FR#48,RFRj,8:F4R8#0_oDFH
O;LHCoM7
Su<mR=FR8jERIC5MR7qu)cRR='2j'R#CDCFR84S;
1Rum<#=RFIjRERCM5Rqc=jR''C2RDR#C#;F4
CSIj=R<RRW NRM850MFR2qc;I
SC<4R= RWR8NMR;qc
zRSjRR:)4qvn7X4RR
RRRRRRRRRRRRRRFRbsl0RN5bR7>R=RR7,q=jR>jRq,4RqRR=>qR4,q=.R>.Rq,dRqRR=>q
d,RSSS7qu)j>R=R)7uqRj,7qu)4>R=R)7uqR4,7qu).>R=R)7uqR.,7qu)d>R=R)7uqRd,
SSSW= R>CRIjW,RBRpi=W>RB,piRm7uRR=>8,FjRm1uRR=>#2Fj;S
Rz:4RRv)q44nX7RR
RRRRRRRRRRRRRbRRFRs0lRNb5=7R>,R7RRqj=q>Rjq,R4>R=R,q4RRq.=q>R.q,Rd>R=R,qd
SRSS)7uq=jR>uR7),qjR)7uq=4R>uR7),q4R)7uq=.R>uR7),q.R)7uq=dR>uR7),qdRS
SSRW =I>RCR4,WiBpRR=>WiBp,uR7m>R=R48F,uR1m>R=R4#F2C;
MX8R)dqv.7X4_
e;
----B-R RppXv)qn4cX7-R--
--DsHLNRs$HCCC;#
kCCRHC#C30D8_FOoH_n44cD3NDk;
#HCRC3CC#_08DHFoOH_#o8MC3DND;H
DLssN$MRkHl#H;#
kCMRkHl#H3FPOlMbFC#M03DND;C

M00H$)RXqcvnXR47HR#
RsbF0
R5RRRRRRRR7RumRRR:FRk0#_08koDFHRO;RRRRR
RRRRRRRRRR1RumRRR:FRk0#_08koDFH
O;
RRRRRRRRRqjR:RRRRHM#_08koDFH
O;RRRRRRRRqR4RRRR:H#MR0k8_DHFoOR;
RRRRRqRR.RRRRH:RM0R#8D_kFOoH;R
RRRRRRdRqRRRR:MRHR8#0_FkDo;HO
RRRRRRRRRqcR:RRRRHM#_08koDFH
O;RRRRRRRRqR6RRRR:H#MR0k8_DHFoOR;
RRRRR7RRRRRRRH:RM0R#8D_kFOoH;R
RRRRRRuR7)Rqj:MRHR8#0_FkDo;HO
RRRRRRRR)7uq:4RRRHM#_08koDFH
O;RRRRRRRR7qu).RR:H#MR0k8_DHFoOR;
RRRRR7RRud)qRH:RM0R#8D_kFOoH;R
RRRRRRuR7)Rqc:MRHR8#0_FkDo;HO
RRRRRRRR)7uq:6RRRHM#_08koDFH
O;RRRRRRRRWiBpRRR:H#MR0k8_DHFoOR;RRRRRRRR
RRRRRWRR RRRRH:RM0R#8D_kFOoH
RRRRRRR2R;R
8CMRqX)vXnc4
7;NEsOHO0C0CksRqX)vXnc4e7_RRFVXv)qn4cX7#RH
SRR#MHoNIDRCRj,I,C4R.IC,CRId#,RFRj,#,F4R.#F,FR#d8,RFRj,8,F4R.8F,FR8d#:R0D8_FOoH;C
Lo
HMSm7uRR<=Rj8FRCIEM7R5u6)qR'=RjN'RM78Ruc)qR'=RjR'2CCD#RS
S8RF4IMECRu57)Rq6=jR''MRN8uR7)Rqc=4R''C2RDR#C
8SSFI.RERCM5)7uq=6RR''4R8NMR)7uq=cRR''j2DRC#
CRSFS8dS;
1Rum<R=R#RFjIMECR65qR'=RjN'RMq8RcRR='2j'R#CDCSR
S4#FRCIEMqR56RR='Rj'NRM8q=cRR''42DRC#
CRSFS#.ERIC5MRq=6RR''4R8NMRRqc=jR''C2RDR#C
#SSF
d;SjICRR<=WN RM58RMRF0qR62NRM850MFR2qc;I
SC<4R= RWR8NMRF5M06Rq2MRN8cRq;I
SC<.R= RWR8NMRRq6NRM850MFR2qc;I
SC<dR= RWR8NMRRq6NRM8q
c;RjSzR):Rqnv4XR47
RRRRRRRRRRRRRRRRsbF0NRlb7R5RR=>7q,Rj>R=R,qjRRq4=q>R4q,R.>R=R,q.RRqd=q>RdR,
S7SSuj)qRR=>7qu)j7,Ru4)qRR=>7qu)47,Ru.)qRR=>7qu).7,Rud)qRR=>7qu)d
,RSWSS >R=RjIC,BRWp=iR>BRWpRi,7Rum=8>RFRj,1Rum=#>RF;j2
zRS4RR:)4qvn7X4RR
RRRRRRRRRRRRRRFRbsl0RN5bR7>R=RR7,q=jR>jRq,4RqRR=>qR4,q=.R>.Rq,dRqRR=>q
d,RSSS7qu)j>R=R)7uqRj,7qu)4>R=R)7uqR4,7qu).>R=R)7uqR.,7qu)d>R=R)7uqRd,
SSSW= R>CRI4W,RBRpi=W>RB,piRm7uRR=>8,F4Rm1uRR=>#2F4;S
Rz:.RRv)q44nX7RR
RRRRRRRRRRRRRbRRFRs0lRNb5=7R>,R7RRqj=q>Rjq,R4>R=R,q4RRq.=q>R.q,Rd>R=R,qd
SRSS)7uq=jR>uR7),qjR)7uq=4R>uR7),q4R)7uq=.R>uR7),q.R)7uq=dR>uR7),qdRS
SSRW =I>RCR.,WiBpRR=>WiBp,uR7m>R=R.8F,uR1m>R=R.#F2R;
SRzd:qR)vX4n4
7RRRRRRRRRRRRRRRRRb0FsRblNRR57=7>R,jRqRR=>qRj,q=4R>4Rq,.RqRR=>qR.,q=dR>dRq,S
RSuS7)Rqj=7>Ruj)q,uR7)Rq4=7>Ru4)q,uR7)Rq.=7>Ru.)q,uR7)Rqd=7>Rud)q,SR
S SWRR=>I,CdRpWBi>R=RpWBi7,Ru=mR>FR8d1,Ru=mR>FR#d
2;CRM8Xv)qn4cX7;_e
-
-

---1-RHDlbCqR)vHRI0#ERHDMoC7Rq71) 1FRVsFRL0sERCRN8NRM8I0sHC-
-RsaNoRC0:HRXDGHM

--
LDHs$NsRCHCCk;
#HCRC3CC#_08DHFoO4_4nNc3D
D;kR#CHCCC38#0_oDFH#O_HCoM8D3NDD;
HNLssk$RMHH#lk;
#kCRMHH#lO3PFFlbM0CM#D3NDC;
M00H$qR)vW_)uR_)HS#
oCCMsRHO5R
SRVRRNDlH$RR:#H0sM:oR=MR"F"MC;S
SI0H8ERR:HCM0oRCs:4=R;SR
S8N8s8IH0:ERR0HMCsoCRR:=nR;RRRRRR-R-RoLHRFCMkRoEVRFs80CbES
S80CbERR:HCM0oRCs:c=RUS;
SFs8ks0_C:oRRFLFDMCNRR:=V#NDCR;RRRRR-E-RNF#Rkk0b0CRsoS
SIk8F0C_soRR:LDFFCRNM:V=RNCD#;-SS-NRE#kRF00bkRosC
8SSHsM_C:oRRFLFDMCNRR:=V#NDCR;RRRRRR-R-R#ENR08NNMRHbRk0s
CoSNSs8_8ssRCo:FRLFNDCM=R:RDVN#RC;RRRRRR--ERN#s8CNR8N8s#C#RosC
ISSNs88_osCRL:RFCFDNRMR:V=RNCD#RRRRR-R-R#ENRHIs0NCR8C8s#s#RCSo
S
2;SsbF0
R5S_S)7amz:kRF00R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj;S
SWm_7z:aRR0FkR8#0_oDFHPO_CFO0sH5I8-0E4FR8IFM0R;j2
)SSq)77RH:RM0R#8F_Do_HOP0COFNs58I8sHE80-84RF0IMF2Rj;S
S7RQhRH:RM0R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj;S
SW7q7)RR:H#MR0D8_FOoH_OPC05FsNs88I0H8ER-48MFI0jFR2S;
SRW RH:RM0R#8F_Do;HORRRRR-RR-sRIHR0CCLMNDVCRFssRNSl
SiBpRH:RM0R#8F_Do;HORRRRR-RR-DROFRO	VRFss,NlR8N8s8,RHSM
Sm)_BRpi:MRHR8#0_oDFHRO;RRRRR-R-R0FbRFODOV	RFssR_k8F0S
SWB_mp:iRRRHM#_08DHFoO-RR-0FbRsVFR8I_F
k0S;S2
8CMR0CMHR0$)_qv)_Wu)
;
---
-HRwsR#0HDlbCMlC0HN0FlMRkR#0LOCRNCDD8sRNO
Ej-N-
sHOE00COkRsCLODF	N_slVRFRv)q_u)W_H)R#F
OlMbFCRM0Xv)qd4.X7RRRb0FsRR5
RRRRR7RRuRmRRF:Rk#0R0k8_DHFoOR;RRRRRRRR
RRRRR1RRuRmRRF:Rk#0R0k8_DHFoO
;
RRRRRRRRqRjRRRR:H#MR0k8_DHFoOR;
RRRRRqRR4RRRRH:RM0R#8D_kFOoH;R
RRRRRR.RqRRRR:MRHR8#0_FkDo;HO
RRRRRRRRRqdR:RRRRHM#_08koDFH
O;RRRRRRRRqRcRRRR:H#MR0k8_DHFoOR;
RRRRR7RRRRRRRH:RM0R#8D_kFOoH;R
RRRRRRuR7)Rqj:MRHR8#0_FkDo;HO
RRRRRRRR)7uq:4RRRHM#_08koDFH
O;RRRRRRRR7qu).RR:H#MR0k8_DHFoOR;
RRRRR7RRud)qRH:RM0R#8D_kFOoH;R
RRRRRRuR7)Rqc:MRHR8#0_FkDo;HO
RRRRRRRRpWBi:RRRRHM#_08koDFHRO;RRRRR
RRRRRRRRRRWR RRRR:H#MR0k8_DHFoOR
RRRRRRR2;RM
C8FROlMbFC;M0
lOFbCFMMX0R)nqvc7X4RbRRFRs05R
RRRRRRuR7mRRR:kRF00R#8D_kFOoH;RRRRRRRRR
RRRRRRuR1mRRR:kRF00R#8D_kFOoH;R

RRRRRqRRjRRRRH:RM0R#8D_kFOoH;R
RRRRRR4RqRRRR:MRHR8#0_FkDo;HO
RRRRRRRRRq.R:RRRRHM#_08koDFH
O;RRRRRRRRqRdRRRR:H#MR0k8_DHFoOR;
RRRRRqRRcRRRRH:RM0R#8D_kFOoH;R
RRRRRR6RqRRRR:MRHR8#0_FkDo;HO
RRRRRRRRR7RR:RRRRHM#_08koDFH
O;RRRRRRRR7qu)jRR:H#MR0k8_DHFoOR;
RRRRR7RRu4)qRH:RM0R#8D_kFOoH;R
RRRRRRuR7)Rq.:MRHR8#0_FkDo;HO
RRRRRRRR)7uq:dRRRHM#_08koDFH
O;RRRRRRRR7qu)cRR:H#MR0k8_DHFoOR;
RRRRR7RRu6)qRH:RM0R#8D_kFOoH;R
RRRRRRBRWpRiR:MRHR8#0_FkDo;HORRRRRRRR
RRRRRRRRRW R:RRRRHM#_08koDFHRO
RRRRR;R2RCR
MO8RFFlbM0CM;k
VMHO0FVMRk_MOH0MH5:LRRFLFDMCN2CRs0MksRs#0HRMoHL#
CMoH
HRRVLR52ER0CRM
RsRRCs0kM"5"2R;
R#CDCR
RRCRs0Mks5F"BkRD8MRF0HDlbCMlC0DRAFRO	)3qvRRQ#0RECs8CNR8N8s#C#RosCHC#0sRC8kM#HoER0CNR#lOCRD	FORRN#0REC)?qv"
2;RMRC8VRH;M
C8kRVMHO_M;H0
MVkOF0HMCRo0M_C8C_8b50E#CHxRH:RMo0CC;sRRb8C0:ERR0HMCsoC2CRs0MksR0HMCsoCR
H#PHNsNCLDRMlH_x#HCRR:HCM0oRCs:j=R;C
Lo
HMRHRlMH_#x:CR=CR8b;0E
HRRV#R5HRxC<CR8b20ERC0EMR
RRHRlMH_#x:CR=HR#x
C;RMRC8VRH;R
RskC0slMRH#M_H;xC
8CMR0oC_8CM_b8C0
E;Ns00H0LkCCRoMNCs0_FssFCbs:0RRs#0H;Mo
0N0skHL0oCRCsMCNs0F_bsCFRs0FLVRD	FO_lsNRN:RsHOE00COkRsCHV#Rk_MOH0MH58sN8ss_C;o2
R--LHCoMDRLFRO	sRNlHDlbCMlC0HN0F#MRHNoMD0#
$RbCH_M0NNss$#RHRsNsN5$RjFR0RR62FHVRMo0CC
s;O#FM00NMR8IH0NE_s$sNRH:RMN0_s$sNRR:=5R4,.c,R,,RgR,4UR2dn;F
OMN#0M80RCEb0_sNsN:$RR0HM_sNsN:$R=4R5ncdU,4RUgR.,cnjg,jR.cRU,4cj.,4R6.
2;O#FM00NMRP8Hd:.RR0HMCsoCRR:=58IH04E-2n/d;F
OMN#0M80RHnP4RH:RMo0CC:sR=IR5HE80-/424
U;O#FM00NMRP8HURR:HCM0oRCs:5=RI0H8E2-4/
g;O#FM00NMRP8HcRR:HCM0oRCs:5=RI0H8E2-4/
c;O#FM00NMRP8H.RR:HCM0oRCs:5=RI0H8E2-4/
.;O#FM00NMRP8H4RR:HCM0oRCs:5=RI0H8E2-4/
4;
MOF#M0N0FRLFRD4:FRLFNDCM=R:RH58P>4RR;j2
MOF#M0N0FRLFRD.:FRLFNDCM=R:RH58P>.RR;j2
MOF#M0N0FRLFRDc:FRLFNDCM=R:RH58P>cRR;j2
MOF#M0N0FRLFRDU:FRLFNDCM=R:RH58P>URR;j2
MOF#M0N0FRLFnD4RL:RFCFDN:MR=8R5HnP4Rj>R2O;
F0M#NRM0LDFFd:.RRFLFDMCNRR:=5P8Hd>.RR;j2
F
OMN#0M80RHnP4dRUc:MRH0CCos=R:RC58b-0E442/ncdU;F
OMN#0M80RH4PUg:.RR0HMCsoCRR:=5b8C04E-24/Ug
.;O#FM00NMRP8HcnjgRH:RMo0CC:sR=8R5CEb0-/42cnjg;F
OMN#0M80RHjP.c:URR0HMCsoCRR:=5b8C04E-2j/.c
U;O#FM00NMRP8H4cj.RH:RMo0CC:sR=8R5CEb0-/424cj.;F
OMN#0M80RH4P6.RR:HCM0oRCs:5=R80CbE2-4/.64;O

F0M#NRM0LDFF6R4.:FRLFNDCM=R:RH58P.64Rj>R2O;
F0M#NRM0LDFF4cj.RL:RFCFDN:MR=8R5HjP4.>cRR;j2
MOF#M0N0FRLFjD.c:URRFLFDMCNRR:=5P8H.UjcRj>R2O;
F0M#NRM0LDFFcnjgRL:RFCFDN:MR=8R5HjPcg>nRR;j2
MOF#M0N0FRLF4DUg:.RRFLFDMCNRR:=5P8HU.4gRj>R2O;
F0M#NRM0LDFF4UndcRR:LDFFCRNM:5=R84HPncdURj>R2
;
O#FM00NMRl#k_8IH0:ERR0HMCsoCRR:=Apmm 'qhb5F#LDFF4+2RRmAmph q'#bF5FLFDR.2+mRAmqp hF'b#F5LF2DcRA+Rm mpqbh'FL#5FUFD2RR+Apmm 'qhb5F#LDFF4;n2
MOF#M0N0kR#lC_8bR0E:MRH0CCos=R:R-6RRm5Amqp hF'b#F5LF4D6.+2RRmAmph q'#bF5FLFD.4jc+2RRmAmph q'#bF5FLFDc.jU+2RRmAmph q'#bF5FLFDgcjn+2RRmAmph q'#bF5FLFDgU4.;22
F
OMN#0MI0R_FOEH_OCI0H8ERR:HCM0oRCs:I=RHE80_sNsN#$5kIl_HE802O;
F0M#NRM0IE_OFCHO_b8C0:ERR0HMCsoCRR:=80CbEs_Ns5N$#_klI0H8E
2;O#FM00NMRO8_EOFHCH_I8R0E:MRH0CCos=R:R8IH0NE_s$sN5l#k_b8C0;E2
MOF#M0N0_R8OHEFO8C_CEb0RH:RMo0CC:sR=CR8b_0ENNss$k5#lC_8b20E;O

F0M#NRM0IH_I8_0EM_klODCD#RR:HCM0oRCs:5=RI0H8E2-4/OI_EOFHCH_I8R0E+;R4
MOF#M0N0_RI80CbEk_MlC_ODRD#:MRH0CCos=R:RC58b-0E4I2/_FOEH_OC80CbERR+4
;
O#FM00NMRI8_HE80_lMk_DOCD:#RR0HMCsoCRR:=58IH04E-2_/8OHEFOIC_HE80R4+R;F
OMN#0M80R_b8C0ME_kOl_C#DDRH:RMo0CC:sR=8R5CEb0-/428E_OFCHO_b8C0+ERR
4;
MOF#M0N0_RI#CHxRH:RMo0CC:sR=_RII0H8Ek_MlC_ODRD#*_RI80CbEk_MlC_OD;D#
MOF#M0N0_R8#CHxRH:RMo0CC:sR=_R8I0H8Ek_MlC_ODRD#*_R880CbEk_MlC_OD;D#
F
OMN#0ML0RF_FD8RR:LDFFCRNM:5=R8H_#x-CRR#I_HRxC<j=R2O;
F0M#NRM0LDFF_:IRRFLFDMCNRR:=M5F0LDFF_;82
F
OMN#0MO0REOFHCH_I8R0E:MRH0CCos=R:Rm5Amqp hF'b#F5LF8D_2RR*8E_OFCHO_8IH0RE2+AR5m mpqbh'FL#5F_FDI*2RROI_EOFHCH_I820E;F
OMN#0MO0REOFHCC_8bR0E:MRH0CCos=R:Rm5Amqp hF'b#F5LF8D_2RR*8E_OFCHO_b8C0RE2+AR5m mpqbh'FL#5F_FDI*2RROI_EOFHCC_8b20E;F
OMN#0MI0RHE80_lMk_DOCD:#RR0HMCsoCRR:=5mAmph q'#bF5FLFD2_8RI*5HE80-/428E_OFCHO_8IH0RE2+AR5m mpqbh'FL#5F_FDI*2RRH5I8-0E4I2/_FOEH_OCI0H8E+2RR
4;O#FM00NMRb8C0ME_kOl_C#DDRH:RMo0CC:sR=AR5m mpqbh'FL#5F_FD8*2R5b8C04E-2_/8OHEFO8C_CEb02RR+5mAmph q'#bF5FLFD2_IR5*R80CbE2-4/OI_EOFHCC_8b20ER4+R;$
0bFCRkL0_k_#40C$bRRH#NNss$8R5CEb0_lMk_DOCD4#-RI8FMR0FjI,RHE80_lMk_DOCD4#-RI8FMR0FjF2RV0R#8F_Do;HO
o#HMRNDs0Fk_#Lk4RR:F_k0L4k#_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFR8s_FRk05bHMk00RFsR0H0-#N#0C2H
#oDMNRkIF0k_L#:4RR0Fk_#Lk4$_0b
C;0C$bR0Fk_#Lk.$_0bHCR#sRNsRN$5b8C0ME_kOl_C#DD-84RF0IMF,RjRI.*HE80_lMk_DOCD4#+RI8FMR0FjF2RV0R#8F_Do;HO
o#HMRNDs0Fk_#Lk.RR:F_k0L.k#_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFR8s_FRk05bHMk00RFsR0H0-#N#0C2H
#oDMNRkIF0k_L#:.RR0Fk_#Lk.$_0b
C;0C$bR0Fk_#Lkc$_0bHCR#sRNsRN$5b8C0ME_kOl_C#DD-84RF0IMF,RjRIc*HE80_lMk_DOCDd#+RI8FMR0FjF2RV0R#8F_Do;HO
o#HMRNDs0Fk_#LkcRR:F_k0Lck#_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFR8s_FRk05bHMk00RFsR0H0-#N#0C2H
#oDMNRkIF0k_L#:cRR0Fk_#Lkc$_0b
C;0C$bR0Fk_#LkU$_0bHCR#sRNsRN$5b8C0ME_kOl_C#DD-84RF0IMF,RjRIU*HE80_lMk_DOCD(#+RI8FMR0FjF2RV0R#8F_Do;HO
o#HMRNDs0Fk_#LkURR:F_k0LUk#_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFR8s_FRk05bHMk00RFsR0H0-#N#0C2H
#oDMNRkIF0k_L#:URR0Fk_#LkU$_0b
C;0C$bRsbNH_0$LUk#_b0$C#RHRsNsN5$R80CbEk_MlC_OD-D#4FR8IFM0RRj,I0H8Ek_MlC_OD-D#4FR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNRNsbs$H0_#LkURR:bHNs0L$_k_#U0C$b;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RV_Rs80FkRM5HbRk000FRs#H-0CN0##2
HNoMDbRIN0sH$k_L#:URRsbNH_0$LUk#_b0$C0;
$RbCF_k0L4k#n$_0bHCR#sRNsRN$5b8C0ME_kOl_C#DD-84RF0IMF,RjR*4nI0H8Ek_MlC_OD+D#486RF0IMF2RjRRFV#_08DHFoO#;
HNoMDFRskL0_kn#4RF:RkL0_kn#4_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$FsVR_k8F0HR5M0bkRR0F0-sH#00NC
#2#MHoNIDRF_k0L4k#nRR:F_k0L4k#n$_0b
C;0C$bRsbNH_0$L4k#n$_0bHCR#sRNsRN$5b8C0ME_kOl_C#DD-84RF0IMF,RjRI.*HE80_lMk_DOCD4#+RI8FMR0FjF2RV0R#8F_Do;HO
o#HMRNDssbNH_0$L4k#nRR:bHNs0L$_kn#4_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFR8s_FRk05bHMk00RFsR0H0-#N#0C2H
#oDMNRNIbs$H0_#Lk4:nRRsbNH_0$L4k#n$_0b
C;0C$bR0Fk_#Lkd0._$RbCHN#Rs$sNRC58b_0EM_klODCD#R-48MFI0jFR,.Rd*8IH0ME_kOl_C#DD+Rd48MFI0jFR2VRFR8#0_oDFH
O;#MHoNsDRF_k0Ldk#.RR:F_k0Ldk#.$_0bRC;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFVsF_8k50RHkMb0FR0RH0s-N#002C#
o#HMRNDI0Fk_#Lkd:.RR0Fk_#Lkd0._$;bC
b0$CNRbs$H0_#Lkd0._$RbCHN#Rs$sNRC58b_0EM_klODCD#R-48MFI0jFR,*RcI0H8Ek_MlC_OD+D#dFR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNRNsbs$H0_#Lkd:.RRsbNH_0$Ldk#.$_0bRC;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RV_Rs80FkRM5HbRk000FRs#H-0CN0##2
HNoMDbRIN0sH$k_L#Rd.:NRbs$H0_#Lkd0._$;bC
o#HMRNDs0Fk_RCM:0R#8F_Do_HOP0COF8s5CEb0_lMk_DOCD4#-RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-C-RMDNLCV#RF0sRs#H-0CN0#H
#oDMNRkIF0M_CR#:R0D8_FOoH_OPC05Fs80CbEk_MlC_OD-D#4FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--CLMNDRC#VRFs0-sH#00NC##
HNoMDsRI0M_CR#:R0D8_FOoH_OPC05Fs80CbEk_MlC_OD-D#4FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--I0sHCMRCNCLD#FRVsNRCOsERFFIRVqR)vCROD
D##MHoNHDRMC_soRR:#_08DHFoOC_POs0F58IH0dE+6FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-#RkC08RFCRso0H#C7sRQ
hR#MHoNsDRF_k0sRCo:0R#8F_Do_HOP0COFIs5HE80+Rd68MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-k-R#RC80sFRC#oH0RCs7amz
o#HMRNDI0Fk_osCR#:R0D8_FOoH_OPC05FsI0H8E6+dRI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--k8#CRR0FsHCo#s0CRz7maH
#oDMNRksF0C_so:4RR8#0_oDFHPO_CFO0sH5I8-0E4FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--k8#CRR0FOFEF#LCRCC0IC7MRQNhRMF8Rkk0b0VRFRFADO)	Rq#v
HNoMDNRs8C_soRR:#_08DHFoOC_POs0F58N8s8IH04E-RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RCk#8FR0RosCHC#0sqR)7
7)#MHoNIDRNs8_C:oRR8#0_oDFHPO_CFO0s85N8HsI8-0E4FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-#RkC08RFCRso0H#CWsRq)77
o#HMRNDD_FIs8N8sRR:#_08DHFoOC_POs0F5R4d8MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--s8N8sHRL0H#RM0bkRR0F)RqvODCD#cR5R0LH#CRsJskHC
82#MHoNDDRFII_Ns88R#:R0D8_FOoH_OPC05Fs48dRF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-I-RNs88R0LH#MRHbRk00)FRqOvRC#DDRR5cL#H0RJsCkCHs8#2
HNoMDqR)7_7)0Rlb:0R#8F_Do_HOP0COFNs58I8sHE80-84RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-k-R#RC80bFRHDbCHRMC)7q7)H
#oDMNR7Wq70)_l:bRR8#0_oDFHPO_CFO0s85N8HsI8-0E4FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-#RkC08RFHRbbHCDMWCRq)77
o#HMRND7_Qh0Rlb:0R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RCk#8FR0RbbHCMDHCQR7hH
#oDMNR_W 0Rlb:0R#8F_Do;HORRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-#RkC08RFHRbbHCDMWCR -
-R8CMRFLDOs	RNHlRlCbDl0CMNF0HMHR#oDMN#-
-RoLCH#MRCODC0NRsllRHblDCCNM00MHFRo#HM#ND
MVkOF0HMCRo0k_Mlc_n5b8C0RE:HCM0o2CsR0sCkRsMHCM0oRCsHP#
NNsHLRDCPRND:MRH0CCos=R:R
j;LHCoMR
RPRND:8=RCEb0/;nc
HRRV5R580CbEFRl8cRn2RR>cRU20MEC
RRRRDPNRR:=PRND+;R4
CRRMH8RVR;
R0sCkRsMP;ND
8CMR0oC_lMk_;nc
MVkOF0HMCRo0C_DVP0FCds_.C58bR0E:MRH0CCoss2RCs0kMMRH0CCos#RH
oLCHRM
R0sCk5sM80CbEFRl8cRn2C;
Mo8RCD0_CFV0P_Csd
.;VOkM0MHFR0oC_VDC0CFPsC58bR0E:MRH0CCosl;RN:GRR0HMCsoC2CRs0MksR0HMCsoCR
H#PHNsNCLDRDPNRH:RMo0CC:sR=;Rj
oLCHRM
RRHV5b8C0-ERRGlNRR>=j02RE
CMRRRRPRND:8=RCEb0Rl-RN
G;RDRC#RC
RPRRN:DR=CR8b;0E
CRRMH8RVR;
R0sCk5sMP2ND;M
C8CRo0C_DVP0FC
s;VOkM0MHFR0oC_lMk_5d.80CbERR:HCM0o2CsR0sCkRsMHCM0oRCsHP#
NNsHLRDCPRND:MRH0CCos=R:R
j;LHCoMR
RH5VR80CbE=R<RRcUNRM880CbERR>4Rn20MEC
RRRRNRPD=R:R
4;RMRC8VRH;R
RskC0sPMRN
D;CRM8o_C0M_kld
.;VOkM0MHFR0oC_lMk_54n80CbERR:HCM0o2CsR0sCkRsMHCM0oRCsHP#
NNsHLRDCPRND:MRH0CCos=R:R
j;LHCoMR
RH5VR80CbE=R<RR4nNRM880CbERR>j02RE
CMRRRRRDPNRR:=4R;
R8CMR;HV
sRRCs0kMNRPDC;
Mo8RCM0_k4l_nO;
F0M#NRM0M_klODCD_Rnc:MRH0CCos=R:R0oC_lMk_5nc80CbE
2;O#FM00NMRVDC0CFPs._dRH:RMo0CC:sR=CRo0C_DVP0FCds_.C58b20E;F
OMN#0MM0RkOl_C_DDd:.RR0HMCsoCRR:=o_C0M_kldD.5CFV0P_Csd;.2
MOF#M0N0CRDVP0FC4s_nRR:HCM0oRCs:o=RCD0_CFV0P5CsD0CVFsPC_,d.R2d.;F
OMN#0MM0RkOl_C_DD4:nRR0HMCsoCRR:=o_C0M_kl4Dn5CFV0P_Cs4;n2
$
0bFCRkL0_k0#_$_bCnRc#HN#Rs$sNRk5MlC_ODnD_cFR8IFM0RRj,I0H8ER-48MFI0jFR2VRFR8#0_oDFH
O;0C$bR0Fk_#Lk_b0$C._d##RHRsNsN5$RM_klODCD_Rd.8MFI0jFR,HRI8-0E4FR8IFM0RRj2F#VR0D8_FOoH;$
0bFCRkL0_k0#_$_bC4Rn#HN#Rs$sNRk5MlC_OD4D_nFR8IFM0RRj,I0H8ER-48MFI0jFR2VRFR8#0_oDFH
O;#MHoNsDRF_k0L_k#nRc#:kRF0k_L#$_0bnC_cR#;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RVFR8k50RHkMb0FR0RH0s-N#002C#
o#HMRNDI0Fk_#Lk_#ncRF:RkL0_k0#_$_bCn;c#RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$F8VRFRk05bHMk00RFsR0H0-#N#0C2H
#oDMNRksF0k_L#._d#RR:F_k0L_k#0C$b_#d.;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFV80FkRM5HbRk000FRs#H-0CN0##2
HNoMDFRIkL0_kd#_.:#RR0Fk_#Lk_b0$C._d##;
HNoMDFRskL0_k4#_n:#RR0Fk_#Lk_b0$Cn_4#R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFRk8F0HR5M0bkRR0F0-sH#00NC
#2#MHoNIDRF_k0L_k#4Rn#:kRF0k_L#$_0b4C_n
#;#MHoNsDRF_k0C#M_R#:R0D8_FOoH_OPC05FsM_klODCD_Rnc8MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-MRCNCLD#FRVssR0H0-#N#0C
o#HMRNDI0Fk__CM#RR:#_08DHFoOC_POs0F5lMk_DOCDc_nRI8FMR0Fj
2;#MHoNsDRF_k0CdM_.RR:#_08DHFoO#;
HNoMDFRIkC0_M._dR#:R0D8_FOoH;H
#oDMNRksF0M_C_R4n:0R#8F_Do;HO
o#HMRNDI0Fk__CM4:nRR8#0_oDFH
O;#MHoNIDRsC0_MR_#:0R#8F_Do_HOP0COFMs5kOl_C_DDn8cRF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RHIs0CCRMDNLCV#RFCsRNROEsRFIF)VRqOvRC#DD
o#HMRNDI_s0CdM_.RR:#_08DHFoO#;
HNoMDsRI0M_C_R4n:0R#8F_Do;HO
o#HMRNDHsM_C#o_R#:R0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--k8#CRR0FsHCo#s0CRh7QRH
#oDMNRksF0C_soR_#:0R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-#RkC08RFCRso0H#C7sRm
za#MHoNIDRF_k0s_Co#RR:#_08DHFoOC_POs0F58IH04E-RI8FMR0FjR2;R#R
HNoMDNRs8C_soR_#:0R#8F_Do_HOP0COFNs58I8sHE80-84RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-k-R#RC80sFRC#oH0RCsq)77
o#HMRNDI_N8s_Co#RR:#_08DHFoOC_POs0F58N8s8IH04E-RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RCk#8FR0RosCHC#0s7Rq7#)
HNoMDFRDIN_s8_8s#RR:#_08DHFoOC_POs0F586RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-N-R8R8sL#H0RbHMk00RFqR)vCRODRD#5LcRHR0#skCJH8sC2H
#oDMNRIDF_8IN8#s_R#:R0D8_FOoH_OPC05Fs6FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-8RN8LsRHR0#HkMb0FR0Rv)qRDOCD5#RcHRL0s#RCHJks2C8
R--CRM8#CCDOs0RNHlRlCbDl0CMNF0HMHR#oDMN#0
N0LsHkR0C\N3slV_FV0#C\RR:#H0sM
o;
oLCHRM
Rdzc:VRHRN5s8_8ss2CoRMoCC0sNC-R-RMoCC0sNCDRLFRO	s
NlRRRR-Q-RV8RN8HsI8R0E<EROFCHO_8IH0NER#o#HMjR''FR0RkkM#RC8L#H0
RRRRRzjRH:RVNR58I8sHE80R4=R2CRoMNCs0SC
RRRRD_FIs8N8s=R<Rj"jjjjjjjjjj"jjRs&RNs8_Cjo52S;
RRRRD_FII8N8s=R<Rj"jjjjjjjjjj"jjRI&RNs8_Cjo52S;
CRM8oCCMsCN0R;zj
RRRRRz4RH:RVNR58I8sHE80R.=R2CRoMNCs0SC
SIDF_8sN8<sR=jR"jjjjjjjjj"jjRs&RNs8_C4o5RI8FMR0Fj
2;SRRRRIDF_8IN8<sR=jR"jjjjjjjjj"jjRI&RNs8_C4o5RI8FMR0Fj
2;S8CMRMoCC0sNC4Rz;R
RR.RzRRR:H5VRNs88I0H8ERR=do2RCsMCN
0CSFSDIN_s8R8s<"=Rjjjjjjjjj"jjRs&RNs8_C.o5RI8FMR0Fj
2;SRRRRIDF_8IN8<sR=jR"jjjjjjjjjRj"&NRI8C_soR5.8MFI0jFR2S;
CRM8oCCMsCN0R;z.
RRRRRzdRH:RVNR58I8sHE80Rc=R2CRoMNCs0SC
SIDF_8sN8<sR=jR"jjjjjjjjj&"RR8sN_osC58dRF0IMF2Rj;R
SRDRRFII_Ns88RR<="jjjjjjjj"jjRI&RNs8_Cdo5RI8FMR0Fj
2;S8CMRMoCC0sNCdRz;R
RRcRzRRR:H5VRNs88I0H8ERR=6o2RCsMCN
0CSRRRRIDF_8sN8<sR=jR"jjjjjjjj"RR&s_N8s5CocFR8IFM0R;j2
RSRRFRDIN_I8R8s<"=Rjjjjjjjjj&"RR8IN_osC58cRF0IMF2Rj;C
SMo8RCsMCNR0Cz
c;RRRRzR6R:VRHR85N8HsI8R0E=2RnRMoCC0sNCR
SRDRRFsI_Ns88RR<="jjjjjjjj&"RR8sN_osC586RF0IMF2Rj;S
SD_FII8N8s=R<Rj"jjjjjjRj"&NRI8C_soR568MFI0jFR2S;
CRM8oCCMsCN0R;z6
RRRRRznRH:RVNR58I8sHE80R(=R2CRoMNCs0SC
RRRRD_FIs8N8s=R<Rj"jjjjjj&"RR8sN_osC58nRF0IMF2Rj;S
SD_FII8N8s=R<Rj"jjjjjj&"RR8IN_osC58nRF0IMF2Rj;C
SMo8RCsMCNR0Cz
n;RRRRzR(R:VRHR85N8HsI8R0E=2RURMoCC0sNCR
SRDRRFsI_Ns88RR<="jjjj"jjRs&RNs8_C(o5RI8FMR0Fj
2;SFSDIN_I8R8s<"=RjjjjjRj"&NRI8C_soR5(8MFI0jFR2S;
CRM8oCCMsCN0R;z(
RRRRRzURH:RVNR58I8sHE80Rg=R2CRoMNCs0SC
RRRRD_FIs8N8s=R<Rj"jj"jjRs&RNs8_CUo5RI8FMR0Fj
2;SFSDIN_I8R8s<"=Rjjjjj&"RR8IN_osC58URF0IMF2Rj;C
SMo8RCsMCNR0Cz
U;RRRRzRgR:VRHR85N8HsI8R0E=jR42CRoMNCs0SC
RRRRD_FIs8N8s=R<Rj"jjRj"&NRs8C_soR5g8MFI0jFR2S;
SIDF_8IN8<sR=jR"j"jjRI&RNs8_Cgo5RI8FMR0Fj
2;S8CMRMoCC0sNCgRz;R
RR4Rzj:RRRRHV58N8s8IH0=ERR244RMoCC0sNCR
SRDRRFsI_Ns88RR<="jjj"RR&s_N8s5Co48jRF0IMF2Rj;S
SD_FII8N8s=R<Rj"jj&"RR8IN_osC5R4j8MFI0jFR2S;
CRM8oCCMsCN0Rjz4;R
RR4Rz4:RRRRHV58N8s8IH0=ERR24.RMoCC0sNCR
SRDRRFsI_Ns88RR<=""jjRs&RNs8_C4o54FR8IFM0R;j2
DSSFII_Ns88RR<=""jjRI&RNs8_C4o54FR8IFM0R;j2
MSC8CRoMNCs0zCR4
4;RRRRzR4.RH:RVNR58I8sHE80R4=Rdo2RCsMCN
0CSRRRRIDF_8sN8<sR=jR''RR&s_N8s5Co48.RF0IMF2Rj;S
SD_FII8N8s=R<R''jRI&RNs8_C4o5.FR8IFM0R;j2
MSC8CRoMNCs0zCR4
.;RRRRzR4dRH:RVNR58I8sHE80R4>Rdo2RCsMCN
0CSRRRRIDF_8sN8<sR=NRs8C_sod54RI8FMR0Fj
2;SRRRRIDF_8IN8<sR=NRI8C_sod54RI8FMR0Fj
2;S8CMRMoCC0sNC4Rzd
;
RRRR-Q-RV8R5HsM_CRo2sHCo#s0CRh7QRHk#MBoRpRi
RzRR4RcR:VRHRH58MC_soo2RCsMCN
0CRRRRRRRRbOsFCR##5iBp,QR7hL2RCMoH
RRRRRRRRRRRRRHV5iBpR'=R4N'RMB8RpCi'P0CM2ER0CRM
RRRRRRRRRRRRRHRRMC_so=R<Rj5"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jjR7&RQ;h2
RRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMRFbsO#C#;C
SMo8RCsMCNR0Cz;4c
RRRR6z4RRR:H5VRMRF08_HMs2CoRMoCC0sNCR
RRRRRRRRRRMRH_osCRR<=5j"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjRj"&QR7h
2;S8CMRMoCC0sNC4Rz6
;
RRRR-Q-RVsR580Fk_osC2CRso0H#C)sR_z7ma#RkHRMo)B_mpRi
RzRR48nsFRk0RH:RVsR580Fk_osC2CRoMNCs0RC
RRRRRbRRsCFO#5#R)B_mpRi,s0Fk_osC2CRLo
HMRRRRRRRRRRRRH5VR)B_mp=iRR''4R8NMRm)_B'piCMPC002RE
CMRRRRRRRRRRRRRRRR)m_7z<aR=FRsks0_C;o4
RRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMRFbsO#C#;R
RRRRRRMRC8CRoMNCs0zCR48nsF;k0
RRRR(z4sk8F0:RRRRHV50MFRFs8ks0_CRo2oCCMsCN0
RRRRRRRRRRRR7)_mRza<s=RF_k0s4Co;C
SMo8RCsMCNR0Czs4(80Fk;S

zI4n80FkRRR:H5VRIk8F0C_soo2RCsMCN
0CRRRRRRRRbOsFCR##5mW_B,piRkIF0C_soL2RCMoH
RRRRRRRRRRRRRHV5mW_BRpi=4R''MRN8_RWmiBp'CCPMR020MEC
RRRRRRRRRRRRRRRR7W_mRza<I=RF_k0s5CoI0H8ER-48MFI0jFR2R;
RRRRRRRRRCRRMH8RVR;
RRRRRCRRMb8RsCFO#
#;RRRRRRRRCRM8oCCMsCN0Rnz4Ik8F0R;
RzRR48(IFRk0RH:RVMR5FI0R80Fk_osC2CRoMNCs0RC
RRRRRRRRRWRR_z7ma=R<RkIF0C_soH5I8-0E4FR8IFM0R;j2
MSC8CRoMNCs0zCR48(IF;k0
R
RR-R-RRQV58sN8ss_CRo2sHCo#s0CR7)q7k)R#oHMRpmBiR
RR4RznRsR:VRHRN5s8_8ss2CoRMoCC0sNC-
-RRRRRRRRbOsFCR##5pmBi),Rq)772CRLo
HM-R-RRRRRRRRRRVRHRB5mp=iRR''4R8NMRpmBiP'CC2M0RC0EM-
-RRRRRRRRRRRRRRRRs_N8sRCo<)=Rq)7758N8s8IH04E-RI8FMR0Fj
2;-R-RRRRRRRRRRMRC8VRH;-
-RRRRRRRRCRM8bOsFC;##
S--CRM8oCCMsCN0Rnz4s-;
-RRRR(z4sRR:H5VRMRF0s8N8sC_soo2RCsMCN
0CRRRRRRRRRRRRs_N8sRCo<)=Rq)77;C
SMo8RCsMCNR0Czs4n;S

-Q-RVIR5Ns88_osC2CRso0H#CWsRq)77RHk#MWoR_pmBiR
RR4RznRIR:VRHRN5I8_8ss2CoRMoCC0sNCR
RRRRRRsRbF#OC#BR5pRi,W7q7)L2RCMoH
RRRRRRRRRRRRRHV5iBpR'=R4N'RMB8RpCi'P0CM2ER0CRM
RRRRRRRRRRRRRIRRNs8_C<oR=qRW757)Ns88I0H8ER-48MFI0jFR2R;
RRRRRRRRRCRRMH8RVR;
RRRRRCRRMb8RsCFO#
#;S8CMRMoCC0sNC4Rzn
I;RRRRzI4(RH:RVMR5FI0RNs88_osC2CRoMNCs0RC
RRRRRRRRRIRRNs8_C<oR=qRW7;7)
MSC8CRoMNCs0zCR4;(I
R
RR-R-R0 GsDNRFOoHRsVFRN7kDFRbsO0RN
#CSCzsoRR:bOsFC5##B2piRoLCHSM
RVRHRp5Bie'  RhaNRM8BRpi=4R''02RE
CMSRRR7_Qh0Rlb<7=RQ
h;SRRR)7q7)l_0b=R<R7)q7
);SRRRW7q7)l_0b=R<R7Wq7
);SRRRW0 _l<bR= RW;R
SR8CMR;HV
MSC8sRbF#OC#
;
SR--Q)VRCRN8qs88CR##=sRWHR0Cqs88C,##RbL$NR##7RQh0FFRkk0b0VRHRRW HC#RMDNLCS8
zGlkRb:RsCFO#W#5 l_0b),Rq)77_b0l,qRW7_7)0,lbRh7Q_b0l,FRsks0_C
o2SLRRCMoH
RSRRVRHRq5W7_7)0Rlb=qR)7_7)0RlbNRM8W0 _l=bRR''42ER0CSM
SsRRF_k0s4CoRR<=7_Qh0;lb
CSSD
#CSRSRs0Fk_osC4=R<RksF0C_soH5I8-0E4FR8IFM0R;j2
CSSMH8RVS;
CRM8bOsFC;##
RSRRRR
R-RR-CRtMNCs00CRE)CRqOvRC#DDR8NMRD#CCRO0DHFoOFRVsqR)vnA4__141S4
zR4U:VRHRE5OFCHO_8IH0=ERRR42oCCMsCN0
RRRR4SzgRR:VRFsHMRHRC58b_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
-S-RRQV58N8s8IH0>ERR24cRCMC8FR0RCOsNR0CI0sHCMRCNCLDR8NMR0FkbRk0CLMND#CRCODC0FRDo
HORRRRRRRRSjz.RH:RVNR58I8sHE80R4>Rco2RCsMCN
0CSR--VRHGVRFsODNDRU4dUR(,#CCDOF0RVsR0HN#00MCRFL0RCoHMRosCHC#0s
C8SSSSs0Fk_5CMH<2R=4R''ERIC5MR)7q7)l_0b85N8HsI8-0E4FR8IFM0R24cRH=R2DRC#'CRj
';SSSSI0Fk_5CMH<2R=4R''ERIC5MRI_N8s5CoNs88I0H8ER-48MFI04FRc=2RRRH2CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R ERIC5MRI_N8s5CoNs88I0H8ER-48MFI04FRc=2RRRH2CCD#R''j;R
RRRRRRCRSMo8RCsMCNR0Cz;.j
-S-RRQV58N8s8IH0<ER=cR42FRMRHIs0CCRMDNLCsRFR0FkbRk0CLMND#CRCODC0FRDoRHOM8CCCR8
SRRRR.Sz4RR:H5VRNs88I0H8E=R<R24cRMoCC0sNCS
SSFSskC0_M25HRR<=';4'
SSSSkIF0M_C5RH2<'=R4
';RRRRRRRRRRRRRRRRI_s0CHM52=R<R;W 
RRRRRRRRMSC8CRoMNCs0zCR.
4;SR--tCCMsCN0RC0ERv)qRDOCDN#RM08Rs#H-0CN0#R
RRRRRRzRS.:.RRsVFRH[RMIR5HE80_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNCR
RRRRRRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqA)vn_4dXUc4:7RRLDNCHDR#WR""R;
RRRRRRRRRRRRRLRRCMoH
RRRRRRRRRRRR)SAq4v_ncdUXR47:qR)vnA4__141S4
RRRRRRRRRRRRb0FsRblNRQ57q25jRR=>HsM_C[o52q,R7q7)RR=>D_FII8N8sd54RI8FMR0FjR2,7RQA=">RjR",q)77A>R=RIDF_8sN84s5dFR8IFM0R,j2
SSSSq hRR=>',4'R)11q>R=R''j, RWq>R=R0Is_5CMHR2,BqpiRR=>B,piRA hRR=>',4'R)11A>R=R''j, RWA>R=R''j,pRBi=AR>pRBiS,
SRSRRmR7q25jRR=>I0Fk_#Lk4,5H[R2,75mAj=2R>FRskL0_k5#4H2,[2
;
RRRRRRRRRRRRRRRRs0Fk_osC5R[2<s=RF_k0L4k#5[H,2ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';SSSSI0Fk_osC5R[2<I=RF_k0L4k#5KH,2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRS8CMRMoCC0sNC.Rz.R;
RRRRS8CMRMoCC0sNC4RzgR;
RCRRMo8RCsMCNR0Cz;4URRRR
RRRR
RRRRRR-t-RCsMCNR0C0REC)RqvODCD#MRN8CR#D0CORoDFHVORF)sRq4vAn._1_
1.Sdz.RH:RVOR5EOFHCH_I8R0E=2R.RMoCC0sNCR
RRzRS.:cRRsVFRHHRM8R5CEb0_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNC-
S-VRQR85N8HsI8R0E>dR42CRMC08RFsROCCN0RHIs0CCRMDNLCMRN8kRF00bkRNCMLRDC#CCDOD0RFOoH
RRRRRRRR.Sz6RR:H5VRNs88I0H8ERR>4Rd2oCCMsCN0
-S-RGVHRsVFRDONDdR4U,U(RD#CCRO0F0VRs0H#NR0CMRF0LMCHoCRso0H#C8sC
RRRRRRRRRRRRRRRRksF0M_C5RH2<'=R4I'RERCM57)q70)_lNb58I8sHE80-84RF0IMFdR42RR=HC2RDR#C';j'
SSSSkIF0M_C5RH2<'=R4I'RERCM58IN_osC58N8s8IH04E-RI8FMR0F4Rd2=2RHR#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=WI RERCM58IN_osC58N8s8IH04E-RI8FMR0F4Rd2=2RHR#CDCjR''R;
RRRRRSRRCRM8oCCMsCN0R6z.;-
S-VRQR85N8HsI8R0E<4=RdM2RFsRIHR0CCLMNDFCRskRF00bkRNCMLRDC#CCDOD0RFOoHRCMC8
C8RRSRRzRS.:nRRRHV58N8s8IH0<ER=dR42CRoMNCs0SC
RRRRRRRRRRRRs0Fk_5CMH<2R=4R''S;
SISSF_k0CHM52=R<R''4;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R R;
RRRRRSRRCRM8oCCMsCN0Rnz.;-
S-CRtMNCs00CRE)CRqOvRC#DDR8NMRH0s-N#00
C#RRRRRRRRS(z.RV:RF[sRRRHM58IH0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CRRRRRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FAVR)_qvU.4gXR.7:NRDLRCDH"#RW
";RRRRRRRRRRRRRRRRLHCoMR
RRRRRRRRRRARS)_qvU.4gXR.7:qR)vnA4__1.1S.
RRRRRRRRRRRRb0FsRblNRQ57q>R=R_HMs5Co.+*[4FR8IFM0R[.*2q,R7q7)RR=>D_FII8N8s.54RI8FMR0FjR2,7RQA=">Rj,j"R7q7)=AR>FRDIN_s858s48.RF0IMF2Rj,S
SSRRRRq hRR=>',4'R)11q>R=R''j, RWq>R=R0Is_5CMHR2,BqpiRR=>B,piRA hRR=>',4'R)11A>R=R''j, RWA>R=R''j,pRBi=AR>pRBiS,
SRSRRmR7q254RR=>I0Fk_#Lk.,5H.+*[4R2,75mqj=2R>FRIkL0_k5#.H*,.[R2,75mA4=2R>FRskL0_k5#.H*,.[2+4,mR7A25jRR=>s0Fk_#Lk.,5HR[.*2
2;RRRRRRRRRRRRRRRRs0Fk_osC5[.*2=R<RksF0k_L#H.5,[.*2ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRs0Fk_osC5[.*+R42<s=RF_k0L.k#5.H,*4[+2ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';SSSSI0Fk_osC5[.*2=R<RkIF0k_L#H.5,[.*2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRI0Fk_osC5[.*+R42<I=RF_k0L.k#5.H,*4[+2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';
RRRRRRRRMSC8CRoMNCs0zCR.
(;RRRRRMSC8CRoMNCs0zCR.
c;RRRRCRM8oCCMsCN0Rdz.;
RR
RSRR-R-RMtCC0sNCER0CqR)vCRODRD#NRM8#CCDOD0RFOoHRsVFRv)qA_4n11c_cz
S.:URRRHV5FOEH_OCI0H8ERR=co2RCsMCN
0CRRRRSgz.RV:RFHsRRRHM5b8C0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CSR--Q5VRNs88I0H8ERR>4R.2M8CCRR0FONsC0ICRsCH0RNCMLRDCNRM8Fbk0kC0RMDNLCCR#D0CORoDFHRO
RRRRRSRRzRdj:VRHR85N8HsI8R0E>.R42CRoMNCs0SC
-V-RHVGRFOsRNRDD4UdU(#,RCODC0VRFRH0s#00NCFRM0CRLHRMosHCo#s0CCR8
RRRRRRRRRRRRRsRRF_k0CHM52=R<R''4RCIEM)R5q)77_b0l58N8s8IH04E-RI8FMR0F4R.2=2RHR#CDCjR''S;
SISSF_k0CHM52=R<R''4RCIEMIR5Ns8_CNo58I8sHE80-84RF0IMF.R42RR-HC2RDR#C';j'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RWRCIEMIR5Ns8_CNo58I8sHE80-84RF0IMF.R42RR=HC2RDR#C';j'
RRRRRRRRMSC8CRoMNCs0zCRd
j;SR--Q5VRNs88I0H8E=R<R24.RRMFI0sHCMRCNCLDRRFsFbk0kC0RMDNLCCR#D0CORoDFHMORCCC88S
RRRRRS4zdRH:RVNR58I8sHE80RR<=4R.2oCCMsCN0
SSSSksF0M_C5RH2<'=R4
';SSSSI0Fk_5CMH<2R=4R''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=W
 ;RRRRRRRRS8CMRMoCC0sNCdRz4S;
-t-RCsMCNR0C0REC)RqvODCD#MRN8sR0H0-#N#0C
RRRRRRRRdSz.RR:VRFs[MRHRH5I8_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
RRRRRRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVAv)q_gcjn7XcRD:RNDLCRRH#";W"
RRRRRRRRRRRRRRRRoLCHRM
RRRRRRRRRSRRAv)q_gcjn7XcR):Rq4vAnc_1_
1cSRRRRRRRRRRRRsbF0NRlb7R5Q=qR>MRH_osC5[c*+8dRF0IMF*Rc[R2,q)77q>R=RIDF_8IN84s54FR8IFM0R,j2RA7QRR=>"jjjjR",q)77A>R=RIDF_8sN84s54FR8IFM0R,j2
SSSSq hRR=>',4'R)11q>R=R''j, RWq>R=R0Is_5CMHR2,BqpiRR=>B,piRA hRR=>',4'R)11A>R=R''j, RWA>R=R''j,pRBi=AR>pRBiS,
S7SSmdq52>R=RkIF0k_L#Hc5,*Rc[2+d,SR
S7SSm.q52>R=RkIF0k_L#Hc5,[c*+,.2RS
SSmS7q254RR=>I0Fk_#Lkc,5Hc+*[4R2,
SSSSq7m5Rj2=I>RF_k0Lck#5RH,c2*[,S
SSmS7A25dRR=>s0Fk_#Lkc,5HR[c*+,d2RS
SSmS7A25.RR=>s0Fk_#Lkc,5Hc+*[.R2,
SSSSA7m5R42=s>RF_k0Lck#5cH,*4[+2
,RSSSS75mAj=2R>FRskL0_k5#cHc,R*2[2;S
SSFSsks0_Cco5*R[2<s=RF_k0Lck#5cH,*R[2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRsks0_Cco5*4[+2=R<RksF0k_L#Hc5,[c*+R42IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRsks0_Cco5*.[+2=R<RksF0k_L#Hc5,[c*+R.2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRsks0_Cco5*d[+2=R<RksF0k_L#Hc5,[c*+Rd2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRIks0_Cco5*R[2<I=RF_k0Lck#5cH,*R[2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRIks0_Cco5*4[+2=R<RkIF0k_L#Hc5,[c*+R42IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRIks0_Cco5*.[+2=R<RkIF0k_L#Hc5,[c*+R.2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRIks0_Cco5*d[+2=R<RkIF0k_L#Hc5,[c*+Rd2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R

RRRRRSRRCRM8oCCMsCN0R.zd;R
RRSRRCRM8oCCMsCN0Rgz.;R
RRMRC8CRoMNCs0zCR.
U;
RSRR-R-RMtCC0sNCER0CqR)vCRODRD#NRM8#CCDOD0RFOoHRsVFRv)qA_4n11g_gz
Sd:dRRRHV5FOEH_OCI0H8ERR=go2RCsMCN
0CRRRRSczdRV:RFHsRRRHM5b8C0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CSR--Q5VRNs88I0H8ERR>4R42M8CCRR0FONsC0ICRsCH0RNCMLRDCNRM8Fbk0kC0RMDNLCCR#D0CORoDFHRO
RRRRRSRRzRd6:VRHR85N8HsI8R0E>4R42CRoMNCs0SC
-V-RHVGRFOsRNRDD4UdU(#,RCODC0VRFRH0s#00NCFRM0CRLHRMosHCo#s0CCR8
RRRRRRRRRRRRRsRRF_k0CHM52=R<R''4RCIEM)R5q)77_b0l58N8s8IH04E-RI8FMR0F4R42=2RHR#CDCjR''S;
SISSF_k0CHM52=R<R''4RCIEMIR5Ns8_CNo58I8sHE80-84RF0IMF4R42RR=HC2RDR#C';j'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RWRCIEMIR5Ns8_CNo58I8sHE80-84RF0IMF4R42RR=HC2RDR#C';j'
RRRRRRRRMSC8CRoMNCs0zCRd
6;SR--Q5VRNs88I0H8E=R<R244RRMFI0sHCMRCNCLDRRFsFbk0kC0RMDNLCCR#D0CORoDFHMORCCC88S
RRRRRSnzdRH:RVNR58I8sHE80RR<=4R42oCCMsCN0
RSRRRRRRRRRRFRskC0_M25HRR<=';4'
SSSSkIF0M_C5RH2<'=R4
';RRRRRRRRRRRRRRRRI_s0CHM52=R<R;W 
RRRRRRRRMSC8CRoMNCs0zCRd
n;SR--tCCMsCN0RC0ERv)qRDOCDN#RM08Rs#H-0CN0#R
RRRRRRzRSd:(RRsVFRH[RMIR5HE80_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNCR
RRRRRRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqA)vj_.cUUX7RR:DCNLD#RHR""W;R
RRRRRRRRRRRRRRCRLo
HMRRRRRRRRRRRRSqA)vj_.cUUX7RR:)Aqv41n_gg_1
RRRRRRRRRRRRRRRRbRRFRs0lRNb5q7QRR=>HsM_Cgo5*([+RI8FMR0Fg2*[,7Rq7R)q=D>RFII_Ns885R4j8MFI0jFR27,RQ=AR>jR"jjjjj"jj,7Rq7R)A=D>RFsI_Ns885R4j8MFI0jFR2R,
RRRRRRRRRRRRRRRRRRRRRRRRR RRh=qR>4R''1,R1R)q='>RjR',WR q=I>RsC0_M25H,pRBi=qR>pRBi ,Rh=AR>4R''1,R1R)A='>RjR',WR A='>RjR',BApiRR=>B,piRR
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7q25(RR=>I0Fk_#LkU,5HU+*[(R2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRq7m5Rn2=I>RF_k0LUk#5UH,*n[+2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mq6=2R>FRIkL0_k5#UH*,U[2+6,RR
RRRRRRRRRRRRRRRRRRRRRRRRR7RRmcq52>R=RkIF0k_L#HU5,[U*+,c2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7q25dRR=>I0Fk_#LkU,5HU+*[dR2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRq7m5R.2=I>RF_k0LUk#5UH,*.[+2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mq4=2R>FRIkL0_k5#UH*,U[2+4,RR
RRRRRRRRRRRRRRRRRRRRRRRRR7RRmjq52>R=RkIF0k_L#HU5,[U*2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mA(=2R>FRskL0_k5#UH*,U[2+(,RR
RRRRRRRRRRRRRRRRRRRRRRRRR7RRmnA52>R=RksF0k_L#HU5,[U*+,n2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7A256RR=>s0Fk_#LkU,5HU+*[6R2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRA7m5Rc2=s>RF_k0LUk#5UH,*c[+2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mAd=2R>FRskL0_k5#UH*,U[2+d,RR
RRRRRRRRRRRRRRRRRRRRRRRRR7RRm.A52>R=RksF0k_L#HU5,[U*+,.2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7A254RR=>s0Fk_#LkU,5HU+*[4R2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRA7m5Rj2=s>RF_k0LUk#5UH,*,[2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRQR7ujq52>R=R_HMs5Cog+*[UR2,7AQuRR=>",j"
RRRRRRRRRRRRRRRRRRRRRRRRRRRRu7mq25jRR=>IsbNH_0$LUk#5[H,27,Rm5uAj=2R>bRsN0sH$k_L#HU5,2[2;R
RRRRRRRRRRRRRRFRsks0_Cgo5*R[2<s=RF_k0LUk#5UH,*R[2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRsks0_Cgo5*4[+2=R<RksF0k_L#HU5,[U*+R42IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRsks0_Cgo5*.[+2=R<RksF0k_L#HU5,[U*+R.2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRsks0_Cgo5*d[+2=R<RksF0k_L#HU5,[U*+Rd2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRsks0_Cgo5*c[+2=R<RksF0k_L#HU5,[U*+Rc2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRsks0_Cgo5*6[+2=R<RksF0k_L#HU5,[U*+R62IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRsks0_Cgo5*n[+2=R<RksF0k_L#HU5,[U*+Rn2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRsks0_Cgo5*([+2=R<RksF0k_L#HU5,[U*+R(2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRsks0_Cgo5*U[+2=R<RNsbs$H0_#LkU,5H[I2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRkIF0C_so*5g[<2R=FRIkL0_k5#UH*,U[I2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRkIF0C_so*5g[2+4RR<=I0Fk_#LkU,5HU+*[4I2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRkIF0C_so*5g[2+.RR<=I0Fk_#LkU,5HU+*[.I2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRkIF0C_so*5g[2+dRR<=I0Fk_#LkU,5HU+*[dI2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRkIF0C_so*5g[2+cRR<=I0Fk_#LkU,5HU+*[cI2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRkIF0C_so*5g[2+6RR<=I0Fk_#LkU,5HU+*[6I2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRkIF0C_so*5g[2+nRR<=I0Fk_#LkU,5HU+*[nI2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRkIF0C_so*5g[2+(RR<=I0Fk_#LkU,5HU+*[(I2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRkIF0C_so*5g[2+URR<=IsbNH_0$LUk#5[H,2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRS8CMRMoCC0sNCdRz(R;
RRRRS8CMRMoCC0sNCdRzcR;
RCRRMo8RCsMCNR0Cz;dd
R
SR-RR-CRtMNCs00CRE)CRqOvRC#DDR8NMRD#CCRO0DHFoOFRVsqR)vnA4_U14_U14
dSzURR:H5VROHEFOIC_HE80R4=RUo2RCsMCN
0CRRRRSgzdRV:RFHsRRRHM5b8C0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CSR--Q5VRNs88I0H8ERR>4Rj2M8CCRR0FONsC0ICRsCH0RNCMLRDCNRM8Fbk0kC0RMDNLCCR#D0CORoDFHRO
RRRRRSRRzRcj:VRHR85N8HsI8R0E>jR42CRoMNCs0SC
-V-RHVGRFOsRNRDD4UdU(#,RCODC0VRFRH0s#00NCFRM0CRLHRMosHCo#s0CCR8
RRRRRRRRRRRRRsRRF_k0CHM52=R<R''4RCIEM)R5q)77_b0l58N8s8IH04E-RI8FMR0F4Rj2=2RHR#CDCjR''S;
SISSF_k0CHM52=R<R''4RCIEMIR5Ns8_CNo58I8sHE80-84RF0IMFjR42RR=HRR2CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R ERIC5MRI_N8s5CoNs88I0H8ER-48MFI04FRj=2RRRH2CCD#R''j;R
RRRRRRCRSMo8RCsMCNR0Cz;cj
-S-RRQV58N8s8IH0<ER=jR42FRMRHIs0CCRMDNLCsRFR0FkbRk0CLMND#CRCODC0FRDoRHOM8CCCR8
SRRRRcSz4RR:H5VRNs88I0H8E=R<R24jRMoCC0sNCR
SRRRRRRRRRsRRF_k0CHM52=R<R''4;S
SSFSIkC0_M25HRR<=';4'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RW;R
RRRRRRCRSMo8RCsMCNR0Cz;c4
-S-RMtCC0sNCER0CqR)vCRODRD#NRM80-sH#00NCR#
RRRRRSRRzRc.:FRVsRR[H5MRI0H8Ek_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0RC
RRRRRRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)RAq4v_jX.c4Rn7:NRDLRCDH"#RW
";RRRRRRRRRRRRRRRRLHCoMR
RRRRRRRRRRARS)_qv4cj.X74nR):Rq4vAn4_1U4_1UR
RRRRRRRRRRRRRRRRRb0FsRblNRQ57q>R=R_HMs5Co4[U*+R468MFI04FRU2*[,7Rq7R)q=D>RFII_Ns8858gRF0IMF2Rj,QR7A>R=Rj"jjjjjjjjjjjjjj,j"R7q7)=AR>FRDIN_s858sgFR8IFM0R,j2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRq hRR=>',4'R)11q>R=R''j, RWq>R=R0Is_5CMHR2,BqpiRR=>B,piRA hRR=>',4'R)11A>R=R''j, RWA>R=R''j,pRBi=AR>pRBi
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mq4R62=I>RF_k0L4k#n,5H4[n*+246,RR
RRRRRRRRRRRRRRRRRRRRRRRRR7RRm4q5c=2R>FRIkL0_kn#454H,n+*[4,c2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7qd542>R=RkIF0k_L#54nHn,4*4[+dR2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRq7m524.RR=>I0Fk_#Lk4Hn5,*4n[.+42
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mq4R42=I>RF_k0L4k#n,5H4[n*+244,RR
RRRRRRRRRRRRRRRRRRRRRRRRR7RRm4q5j=2R>FRIkL0_kn#454H,n+*[4,j2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7q25gRR=>I0Fk_#Lk4Hn5,*4n[2+g,RR
RRRRRRRRRRRRRRRRRRRRRRRRR7RRmUq52>R=RkIF0k_L#54nHn,4*U[+2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mq(=2R>FRIkL0_kn#454H,n+*[(R2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRq7m5Rn2=I>RF_k0L4k#n,5H4[n*+,n2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7q256RR=>I0Fk_#Lk4Hn5,*4n[2+6,RR
RRRRRRRRRRRRRRRRRRRRRRRRR7RRmcq52>R=RkIF0k_L#54nHn,4*c[+2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mqd=2R>FRIkL0_kn#454H,n+*[dR2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRq7m5R.2=I>RF_k0L4k#n,5H4[n*+,.2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7q254RR=>I0Fk_#Lk4Hn5,*4n[2+4,RR
RRRRRRRRRRRRRRRRRRRRRRRRR7RRmjq52>R=RkIF0k_L#54nHn,4*,[2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7A6542>R=RksF0k_L#54nHn,4*4[+6R2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRA7m524cRR=>s0Fk_#Lk4Hn5,*4n[c+42
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mA4Rd2=s>RF_k0L4k#n,5H4[n*+24d,RR
RRRRRRRRRRRRRRRRRRRRRRRRR7RRm4A5.=2R>FRskL0_kn#454H,n+*[4,.2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7A4542>R=RksF0k_L#54nHn,4*4[+4R2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRA7m524jRR=>s0Fk_#Lk4Hn5,*4n[j+42
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mAg=2R>FRskL0_kn#454H,n+*[gR2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRA7m5RU2=s>RF_k0L4k#n,5H4[n*+,U2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7A25(RR=>s0Fk_#Lk4Hn5,*4n[2+(,RR
RRRRRRRRRRRRRRRRRRRRRRRRR7RRmnA52>R=RksF0k_L#54nHn,4*n[+2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mA6=2R>FRskL0_kn#454H,n+*[6R2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRA7m5Rc2=s>RF_k0L4k#n,5H4[n*+,c2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7A25dRR=>s0Fk_#Lk4Hn5,*4n[2+d,RR
RRRRRRRRRRRRRRRRRRRRRRRRR7RRm.A52>R=RksF0k_L#54nHn,4*.[+2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mA4=2R>FRskL0_kn#454H,n+*[4R2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRA7m5Rj2=s>RF_k0L4k#n,5H4[n*2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRR7qQuRR=>HsM_C4o5U+*[48(RF0IMFUR4*4[+nR2,7AQuRR=>""jj,R
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7u4q52>R=RNIbs$H0_#Lk4Hn5,[.*+,42Ru7mq25jRR=>IsbNH_0$L4k#n,5H.2*[,R
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7u4A52>R=RNsbs$H0_#Lk4Hn5,[.*+,42Ru7mA25jRR=>ssbNH_0$L4k#n,5H.2*[2R;
RRRRRRRRRRRRRsRRF_k0s5Co4[U*2=R<RksF0k_L#54nHn,4*R[2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRsks0_C4o5U+*[4<2R=FRskL0_kn#454H,n+*[4I2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRksF0C_soU54*.[+2=R<RksF0k_L#54nHn,4*.[+2ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRs0Fk_osC5*4U[2+dRR<=s0Fk_#Lk4Hn5,*4n[2+dRCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRsRRF_k0s5Co4[U*+Rc2<s=RF_k0L4k#n,5H4[n*+Rc2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRsks0_C4o5U+*[6<2R=FRskL0_kn#454H,n+*[6I2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRksF0C_soU54*n[+2=R<RksF0k_L#54nHn,4*n[+2ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRs0Fk_osC5*4U[2+(RR<=s0Fk_#Lk4Hn5,*4n[2+(RCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRsRRF_k0s5Co4[U*+RU2<s=RF_k0L4k#n,5H4[n*+RU2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRsks0_C4o5U+*[g<2R=FRskL0_kn#454H,n+*[gI2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRksF0C_soU54*4[+j<2R=FRskL0_kn#454H,n+*[4Rj2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRsks0_C4o5U+*[4R42<s=RF_k0L4k#n,5H4[n*+244RCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRsRRF_k0s5Co4[U*+24.RR<=s0Fk_#Lk4Hn5,*4n[.+42ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRs0Fk_osC5*4U[d+42=R<RksF0k_L#54nHn,4*4[+dI2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRksF0C_soU54*4[+c<2R=FRskL0_kn#454H,n+*[4Rc2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRsks0_C4o5U+*[4R62<s=RF_k0L4k#n,5H4[n*+246RCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRsRRF_k0s5Co4[U*+24nRR<=ssbNH_0$L4k#n,5H.2*[RCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRsRRF_k0s5Co4[U*+24(RR<=ssbNH_0$L4k#n,5H.+*[4I2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
R
RRRRRRRRRRRRRRFRIks0_C4o5U2*[RR<=I0Fk_#Lk4Hn5,*4n[I2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRkIF0C_soU54*4[+2=R<RkIF0k_L#54nHn,4*4[+2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRI0Fk_osC5*4U[2+.RR<=I0Fk_#Lk4Hn5,*4n[2+.RCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRIRRF_k0s5Co4[U*+Rd2<I=RF_k0L4k#n,5H4[n*+Rd2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRIks0_C4o5U+*[c<2R=FRIkL0_kn#454H,n+*[cI2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRkIF0C_soU54*6[+2=R<RkIF0k_L#54nHn,4*6[+2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRI0Fk_osC5*4U[2+nRR<=I0Fk_#Lk4Hn5,*4n[2+nRCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRIRRF_k0s5Co4[U*+R(2<I=RF_k0L4k#n,5H4[n*+R(2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRIks0_C4o5U+*[U<2R=FRIkL0_kn#454H,n+*[UI2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRkIF0C_soU54*g[+2=R<RkIF0k_L#54nHn,4*g[+2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRI0Fk_osC5*4U[j+42=R<RkIF0k_L#54nHn,4*4[+jI2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRkIF0C_soU54*4[+4<2R=FRIkL0_kn#454H,n+*[4R42IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRIks0_C4o5U+*[4R.2<I=RF_k0L4k#n,5H4[n*+24.RCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRIRRF_k0s5Co4[U*+24dRR<=I0Fk_#Lk4Hn5,*4n[d+42ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRI0Fk_osC5*4U[c+42=R<RkIF0k_L#54nHn,4*4[+cI2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRkIF0C_soU54*4[+6<2R=FRIkL0_kn#454H,n+*[4R62IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRIks0_C4o5U+*[4Rn2<I=RbHNs0L$_kn#45.H,*R[2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRIks0_C4o5U+*[4R(2<I=RbHNs0L$_kn#45.H,*4[+2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';
RRRRRRRRMSC8CRoMNCs0zCRc
.;RRRRRMSC8CRoMNCs0zCRd
g;RRRRCRM8oCCMsCN0RUzd;S

RRRR-t-RCsMCNR0C0REC)RqvODCD#MRN8CR#D0CORoDFHVORF)sRq4vAnd_1nd_1nz
SdRUN:VRHRE5OFCHO_8IH0=ERR2dnRMoCC0sNCR
SRzRRdRgN:FRVsRRHH5MR80CbEk_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0SC
-Q-RVNR58I8sHE80Rg>R2CRMC08RFsROCCN0RHIs0CCRMDNLCMRN8kRF00bkRNCMLRDC#CCDOD0RFOoH
SSSzNcjRH:RVNR58I8sHE80Rg>R2CRoMNCs0SC
-V-RHVGRFOsRNRDD4UdU(#,RCODC0VRFRH0s#00NCFRM0CRLHRMosHCo#s0CCS8
SsSSF_k0CHM52=R<R''4RCIEM)R5q)77_b0l58N8s8IH04E-RI8FMR0Fg=2RRRH2CCD#R''j;S
SSFSIkC0_M25HRR<='R4'IMECRN5I8C_so85N8HsI8-0E4FR8IFM0RRg2=RRH2DRC#'CRj
';SSSSI_s0CHM52=R<RRW IMECRN5I8C_so85N8HsI8-0E4FR8IFM0RRg2=2RHR#CDCjR''S;
SMSC8CRoMNCs0zCRc;jN
-S-RRQV58N8s8IH0<ER=2RgRRMFI0sHCMRCNCLDRRFsFbk0kC0RMDNLCCR#D0CORoDFHMORCCC88S
SS4zcNRR:H5VRNs88I0H8E=R<RRg2oCCMsCN0
SSSSksF0M_C5RH2<'=R4
';SSSSI0Fk_5CMH<2R=4R''S;
SISSsC0_M25HRR<=W
 ;SCSSMo8RCsMCNR0CzNc4;-
S-CRtMNCs00CRE)CRqOvRC#DDR8NMRH0s-N#00
C#SzSScR.N:FRVsRR[H5MRI0H8Ek_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0RC
RRRRRRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)RAq6v_4d.X.:7RRLDNCHDR#WR""R;
RRRRRRRRRRRRRLRRCMoH
RRRRRRRRRRRRRRRRARR)_qv6X4.dR.7:qR)vnA4_n1d_n1d
RRRRRRRRRRRRRRRRRRRRsbF0NRlb7R5Q=qR>MRH_osC5*dn[4+dRI8FMR0Fd[n*2q,R7q7)RR=>D_FII8N8sR5U8MFI0jFR27,RQ=AR>jR"jjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj,7Rq7R)A=D>RFsI_Ns8858URF0IMF2Rj,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR Rhq='>R4R',1q1)RR=>',j'RqW RR=>I_s0CHM52B,RpRiq=B>RpRi, RhA='>R4R',1A1)RR=>',j'RAW RR=>',j'RiBpA>R=RiBp,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mqdR42=I>RF_k0Ldk#.,5Hd[.*+2d4,RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRq7m52djRR=>I0Fk_#LkdH.5,*d.[j+d2R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRq7m52.gRR=>I0Fk_#LkdH.5,*d.[g+.2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7qU5.2>R=RkIF0k_L#5d.H.,d*.[+UR2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRm.q5(=2R>FRIkL0_k.#d5dH,.+*[.,(2
RRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRm.q5n=2R>FRIkL0_k.#d5dH,.+*[.,n2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mq.R62=I>RF_k0Ldk#.,5Hd[.*+2.6,RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRq7m52.cRR=>I0Fk_#LkdH.5,*d.[c+.2R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRq7m52.dRR=>I0Fk_#LkdH.5,*d.[d+.2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7q.5.2>R=RkIF0k_L#5d.H.,d*.[+.R2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRm.q54=2R>FRIkL0_k.#d5dH,.+*[.,42
RRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRm.q5j=2R>FRIkL0_k.#d5dH,.+*[.,j2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mq4Rg2=I>RF_k0Ldk#.,5Hd[.*+24g,RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRq7m524URR=>I0Fk_#LkdH.5,*d.[U+42R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRq7m524(RR=>I0Fk_#LkdH.5,*d.[(+42
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7qn542>R=RkIF0k_L#5d.H.,d*4[+nR2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRm4q56=2R>FRIkL0_k.#d5dH,.+*[4,62
RRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRm4q5c=2R>FRIkL0_k.#d5dH,.+*[4,c2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mq4Rd2=I>RF_k0Ldk#.,5Hd[.*+24d,RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRq7m524.RR=>I0Fk_#LkdH.5,*d.[.+42R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRq7m5244RR=>I0Fk_#LkdH.5,*d.[4+42
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7qj542>R=RkIF0k_L#5d.H.,d*4[+jR2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRmgq52>R=RkIF0k_L#5d.H.,d*g[+2R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRq7m5RU2=I>RF_k0Ldk#.,5Hd[.*+,U2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mq(=2R>FRIkL0_k.#d5dH,.+*[(R2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRmnq52>R=RkIF0k_L#5d.H.,d*n[+2R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRq7m5R62=I>RF_k0Ldk#.,5Hd[.*+,62RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mqc=2R>FRIkL0_k.#d5dH,.+*[cR2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRmdq52>R=RkIF0k_L#5d.H.,d*d[+2R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRq7m5R.2=I>RF_k0Ldk#.,5Hd[.*+,.2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mq4=2R>FRIkL0_k.#d5dH,.+*[4R2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRmjq52>R=RkIF0k_L#5d.H.,d*,[2
RRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRmdA54=2R>FRskL0_k.#d5dH,.+*[d,42RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mAdRj2=s>RF_k0Ldk#.,5Hd[.*+2dj,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mA.Rg2=s>RF_k0Ldk#.,5Hd[.*+2.g,RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRA7m52.URR=>s0Fk_#LkdH.5,*d.[U+.2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7A(5.2>R=RksF0k_L#5d.H.,d*.[+(
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7An5.2>R=RksF0k_L#5d.H.,d*.[+nR2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRm.A56=2R>FRskL0_k.#d5dH,.+*[.,62RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mA.Rc2=s>RF_k0Ldk#.,5Hd[.*+2.c,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mA.Rd2=s>RF_k0Ldk#.,5Hd[.*+2.d,RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRA7m52..RR=>s0Fk_#LkdH.5,*d.[.+.2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7A45.2>R=RksF0k_L#5d.H.,d*.[+4
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7Aj5.2>R=RksF0k_L#5d.H.,d*.[+jR2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRm4A5g=2R>FRskL0_k.#d5dH,.+*[4,g2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mA4RU2=s>RF_k0Ldk#.,5Hd[.*+24U,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mA4R(2=s>RF_k0Ldk#.,5Hd[.*+24(,RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRA7m524nRR=>s0Fk_#LkdH.5,*d.[n+42
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7A6542>R=RksF0k_L#5d.H.,d*4[+6
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7Ac542>R=RksF0k_L#5d.H.,d*4[+cR2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRm4A5d=2R>FRskL0_k.#d5dH,.+*[4,d2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mA4R.2=s>RF_k0Ldk#.,5Hd[.*+24.,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mA4R42=s>RF_k0Ldk#.,5Hd[.*+244,RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRA7m524jRR=>s0Fk_#LkdH.5,*d.[j+42
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7A25gRR=>s0Fk_#LkdH.5,*d.[2+g,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mAU=2R>FRskL0_k.#d5dH,.+*[UR2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRm(A52>R=RksF0k_L#5d.H.,d*([+2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7A25nRR=>s0Fk_#LkdH.5,*d.[2+n,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mA6=2R>FRskL0_k.#d5dH,.+*[6R2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRmcA52>R=RksF0k_L#5d.H.,d*c[+2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7A25dRR=>s0Fk_#LkdH.5,*d.[2+d,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mA.=2R>FRskL0_k.#d5dH,.+*[.R2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRm4A52>R=RksF0k_L#5d.H.,d*4[+2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7A25jRR=>s0Fk_#LkdH.5,*d.[
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRQR7u=qR>MRH_osC5*dn[6+dRI8FMR0Fd[n*+2d.,QR7u=AR>jR"j"jj,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR7qmu5Rd2=I>RbHNs0L$_k.#d5cH,*d[+27,Rm5uq.=2R>bRIN0sH$k_L#5d.H*,c[2+.,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR7qmu5R42=I>RbHNs0L$_k.#d5cH,*4[+27,Rm5uqj=2R>bRIN0sH$k_L#5d.H*,c[
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7udA52>R=RNsbs$H0_#LkdH.5,[c*+,d2Ru7mA25.RR=>ssbNH_0$Ldk#.,5Hc+*[.
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7u4A52>R=RNsbs$H0_#LkdH.5,[c*+,42Ru7mA25jRR=>ssbNH_0$Ldk#.,5Hc2*[2R;
RRRRRRRRRRRRRRRRRksF0C_son5d*R[2<s=RF_k0Ldk#.,5Hd[.*2ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRsks0_Cdo5n+*[4<2R=FRskL0_k.#d5dH,.+*[4I2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRsRRF_k0s5Cod[n*+R.2<s=RF_k0Ldk#.,5Hd[.*+R.2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRs0Fk_osC5*dn[2+dRR<=s0Fk_#LkdH.5,*d.[2+dRCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRksF0C_son5d*c[+2=R<RksF0k_L#5d.H.,d*c[+2ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRsks0_Cdo5n+*[6<2R=FRskL0_k.#d5dH,.+*[6I2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRsRRF_k0s5Cod[n*+Rn2<s=RF_k0Ldk#.,5Hd[.*+Rn2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRs0Fk_osC5*dn[2+(RR<=s0Fk_#LkdH.5,*d.[2+(RCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRksF0C_son5d*U[+2=R<RksF0k_L#5d.H.,d*U[+2ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRsks0_Cdo5n+*[g<2R=FRskL0_k.#d5dH,.+*[gI2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRsRRF_k0s5Cod[n*+24jRR<=s0Fk_#LkdH.5,*d.[j+42ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRsks0_Cdo5n+*[4R42<s=RF_k0Ldk#.,5Hd[.*+244RCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRksF0C_son5d*4[+.<2R=FRskL0_k.#d5dH,.+*[4R.2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRs0Fk_osC5*dn[d+42=R<RksF0k_L#5d.H.,d*4[+dI2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRsRRF_k0s5Cod[n*+24cRR<=s0Fk_#LkdH.5,*d.[c+42ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRsks0_Cdo5n+*[4R62<s=RF_k0Ldk#.,5Hd[.*+246RCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRksF0C_son5d*4[+n<2R=FRskL0_k.#d5dH,.+*[4Rn2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRs0Fk_osC5*dn[(+42=R<RksF0k_L#5d.H.,d*4[+(I2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRsRRF_k0s5Cod[n*+24URR<=s0Fk_#LkdH.5,*d.[U+42ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRsks0_Cdo5n+*[4Rg2<s=RF_k0Ldk#.,5Hd[.*+24gRCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRksF0C_son5d*.[+j<2R=FRskL0_k.#d5dH,.+*[.Rj2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRs0Fk_osC5*dn[4+.2=R<RksF0k_L#5d.H.,d*.[+4I2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRsRRF_k0s5Cod[n*+2..RR<=s0Fk_#LkdH.5,*d.[.+.2ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRsks0_Cdo5n+*[.Rd2<s=RF_k0Ldk#.,5Hd[.*+2.dRCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRksF0C_son5d*.[+c<2R=FRskL0_k.#d5dH,.+*[.Rc2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRs0Fk_osC5*dn[6+.2=R<RksF0k_L#5d.H.,d*.[+6I2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRsRRF_k0s5Cod[n*+2.nRR<=s0Fk_#LkdH.5,*d.[n+.2ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRsks0_Cdo5n+*[.R(2<s=RF_k0Ldk#.,5Hd[.*+2.(RCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRksF0C_son5d*.[+U<2R=FRskL0_k.#d5dH,.+*[.RU2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRs0Fk_osC5*dn[g+.2=R<RksF0k_L#5d.H.,d*.[+gI2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRsRRF_k0s5Cod[n*+2djRR<=s0Fk_#LkdH.5,*d.[j+d2ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRsks0_Cdo5n+*[dR42<s=RF_k0Ldk#.,5Hd[.*+2d4RCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRksF0C_son5d*d[+.<2R=bRsN0sH$k_L#5d.H*,c[I2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRsRRF_k0s5Cod[n*+2ddRR<=ssbNH_0$Ldk#.,5Hc+*[4I2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRsRRF_k0s5Cod[n*+2dcRR<=ssbNH_0$Ldk#.,5Hc+*[.I2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRsRRF_k0s5Cod[n*+2d6RR<=ssbNH_0$Ldk#.,5Hc+*[dI2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR
RRRRRRRRRRRRRRRRRRRFRIks0_Cdo5n2*[RR<=I0Fk_#LkdH.5,*d.[I2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRIRRF_k0s5Cod[n*+R42<I=RF_k0Ldk#.,5Hd[.*+R42IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRI0Fk_osC5*dn[2+.RR<=I0Fk_#LkdH.5,*d.[2+.RCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRkIF0C_son5d*d[+2=R<RkIF0k_L#5d.H.,d*d[+2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRIks0_Cdo5n+*[c<2R=FRIkL0_k.#d5dH,.+*[cI2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRIRRF_k0s5Cod[n*+R62<I=RF_k0Ldk#.,5Hd[.*+R62IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRI0Fk_osC5*dn[2+nRR<=I0Fk_#LkdH.5,*d.[2+nRCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRkIF0C_son5d*([+2=R<RkIF0k_L#5d.H.,d*([+2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRIks0_Cdo5n+*[U<2R=FRIkL0_k.#d5dH,.+*[UI2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRIRRF_k0s5Cod[n*+Rg2<I=RF_k0Ldk#.,5Hd[.*+Rg2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRI0Fk_osC5*dn[j+42=R<RkIF0k_L#5d.H.,d*4[+jI2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRIRRF_k0s5Cod[n*+244RR<=I0Fk_#LkdH.5,*d.[4+42ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRIks0_Cdo5n+*[4R.2<I=RF_k0Ldk#.,5Hd[.*+24.RCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRkIF0C_son5d*4[+d<2R=FRIkL0_k.#d5dH,.+*[4Rd2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRI0Fk_osC5*dn[c+42=R<RkIF0k_L#5d.H.,d*4[+cI2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRIRRF_k0s5Cod[n*+246RR<=I0Fk_#LkdH.5,*d.[6+42ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRIks0_Cdo5n+*[4Rn2<I=RF_k0Ldk#.,5Hd[.*+24nRCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRkIF0C_son5d*4[+(<2R=FRIkL0_k.#d5dH,.+*[4R(2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRI0Fk_osC5*dn[U+42=R<RkIF0k_L#5d.H.,d*4[+UI2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRIRRF_k0s5Cod[n*+24gRR<=I0Fk_#LkdH.5,*d.[g+42ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRIks0_Cdo5n+*[.Rj2<I=RF_k0Ldk#.,5Hd[.*+2.jRCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRkIF0C_son5d*.[+4<2R=FRIkL0_k.#d5dH,.+*[.R42IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRI0Fk_osC5*dn[.+.2=R<RkIF0k_L#5d.H.,d*.[+.I2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRIRRF_k0s5Cod[n*+2.dRR<=I0Fk_#LkdH.5,*d.[d+.2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRIks0_Cdo5n+*[.Rc2<I=RF_k0Ldk#.,5Hd[.*+2.cRCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRkIF0C_son5d*.[+6<2R=FRIkL0_k.#d5dH,.+*[.R62IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRI0Fk_osC5*dn[n+.2=R<RkIF0k_L#5d.H.,d*.[+nI2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRIRRF_k0s5Cod[n*+2.(RR<=I0Fk_#LkdH.5,*d.[(+.2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRIks0_Cdo5n+*[.RU2<I=RF_k0Ldk#.,5Hd[.*+2.URCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRkIF0C_son5d*.[+g<2R=FRIkL0_k.#d5dH,.+*[.Rg2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRI0Fk_osC5*dn[j+d2=R<RkIF0k_L#5d.H.,d*d[+jI2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRIRRF_k0s5Cod[n*+2d4RR<=I0Fk_#LkdH.5,*d.[4+d2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRIks0_Cdo5n+*[dR.2<I=RbHNs0L$_k.#d5cH,*R[2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRI0Fk_osC5*dn[d+d2=R<RNIbs$H0_#LkdH.5,[c*+R42IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRI0Fk_osC5*dn[c+d2=R<RNIbs$H0_#LkdH.5,[c*+R.2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRI0Fk_osC5*dn[6+d2=R<RNIbs$H0_#LkdH.5,[c*+Rd2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;S

SMSC8CRoMNCs0zCRc;.N
CSSMo8RCsMCNR0CzNdg;C
SMo8RCsMCNR0CzNdU;R
RCRM8oCCMsCN0Rdzc;R

RczcRH:RVMR5Fs0RNs88_osC2CRoMNCs0-CR-CRoMNCs0#CRCODC0NRslR
RR-R-RRQVNs88I0H8ERR<6#RN#MHoR''jRR0Fk#MkCL8RH
0#RRRRzRjR:VRHR85N8HsI8R0E=2R4RMoCC0sNCR
RRRRRRFRDIN_s8_8s#=R<Rj"jj"jjRs&RNs8_C#o_5;j2
RRRRRRRRIDF_8IN8#s_RR<="jjjjRj"&NRI8C_so5_#j
2;RRRRCRM8oCCMsCN0R;zj
RRRRRz4RH:RVNR58I8sHE80R.=R2CRoMNCs0RC
RRRRRDRRFsI_Ns88_<#R=jR"j"jjRs&RNs8_C#o_584RF0IMF2Rj;R
RRRRRRFRDIN_I8_8s#=R<Rj"jjRj"&NRI8C_so5_#4FR8IFM0R;j2
RRRR8CMRMoCC0sNC4Rz;R
RR.RzRRR:H5VRNs88I0H8ERR=do2RCsMCN
0CRRRRRRRRD_FIs8N8sR_#<"=Rj"jjRs&RNs8_C#o_58.RF0IMF2Rj;R
RRRRRRFRDIN_I8_8s#=R<Rj"jj&"RR8IN_osC_.#5RI8FMR0Fj
2;RRRRCRM8oCCMsCN0R;z.
RRRRRzdRH:RVNR58I8sHE80Rc=R2CRoMNCs0RC
RRRRRDRRFsI_Ns88_<#R=jR"j&"RR8sN_osC_d#5RI8FMR0Fj
2;RRRRRRRRD_FII8N8sR_#<"=RjRj"&NRI8C_so5_#dFR8IFM0R;j2
RRRR8CMRMoCC0sNCdRz;z
ScRS:H5VRNs88I0H8ERR=6o2RCsMCN
0CSFSDIN_s8_8s#=R<R''jRs&RNs8_C#o_58cRF0IMF2Rj;S
SD_FII8N8sR_#<'=Rj&'RR8IN_osC_c#5RI8FMR0Fj
2;S8CMRMoCC0sNCcRz;R
RR6RzRRR:H5VRNs88I0H8ERR>6o2RCsMCN
0CRRRRRRRRD_FIs8N8sR_#<s=RNs8_C#o_586RF0IMF2Rj;R
RRRRRRFRDIN_I8_8s#=R<R8IN_osC_6#5RI8FMR0Fj
2;RRRRCRM8oCCMsCN0R;z6
R
RR-R-RRQV5M8H_osC2CRso0H#C7sRQkhR#oHMRiBp
RRRRRznRH:RV8R5HsM_CRo2oCCMsCN0
RRRRRRRRFbsO#C#Rp5Bi7,RQRh2LHCoMR
RRRRRRRRRRVRHRp5BiRR='R4'NRM8B'piCMPC002RE
CMRRRRRRRRRRRRRRRRHsM_C#o_RR<=7;Qh
RRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMRFbsO#C#;R
RRMRC8CRoMNCs0zCRnR;
RzRR(:RRRRHV50MFRM8H_osC2CRoMNCs0RC
RRRRRRRRRHRRMC_soR_#<7=RQ
h;RRRRCRM8oCCMsCN0R;z(
R
RR-R-RRQV5Fs8ks0_CRo2sHCo#s0CRz7ma#RkHRMomiBp
RRRRszURRR:H5VRsk8F0C_soo2RCsMCN
0CRRRRRRRRbOsFCR##5m)_B,piRksF0C_so2_#RoLCHRM
RRRRRRRRRHRRV)R5_pmBiRR='R4'NRM8)B_mpCi'P0CM2ER0CRM
RRRRRRRRRRRRR)RR_z7ma=R<RksF0C_so;_#
RRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMRFbsO#C#;R
RRMRC8CRoMNCs0zCRU
s;RRRRzRgsRH:RVMR5Fs0R80Fk_osC2CRoMNCs0RC
RRRRRRRRR)RR_z7ma=R<RksF0C_so;_#
RRRR8CMRMoCC0sNCgRzs
;
SIzURRR:H5VRIk8F0C_soo2RCsMCN
0CRRRRRRRRbOsFCR##5mW_B,piRkIF0C_so2_#RoLCHRM
RRRRRRRRRHRRVWR5_pmBiRR='R4'NRM8WB_mpCi'P0CM2ER0CRM
RRRRRRRRRRRRRWRR_z7ma=R<RkIF0C_so;_#
RRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMRFbsO#C#;R
RRMRC8CRoMNCs0zCRU
I;RRRRzRgIRH:RVMR5FI0R80Fk_osC2CRoMNCs0RC
RRRRRRRRRWRR_z7ma=R<RkIF0C_so;_#
RRRR8CMRMoCC0sNCgRzI
;
RRRR-Q-RVsR5Ns88_osC2CRso0H#CqsR7R7)kM#HopRBiR
RR4Rzj:RRRRHV58sN8ss_CRo2oCCMsCN0
RRRRRRRRFbsO#C#R_5)miBp,qR)727)RoLCHRM
RRRRRRRRRHRRV)R5_pmBiRR='R4'NRM8)B_mpCi'P0CM2ER0CRM
RRRRRRRRRRRRRsRRNs8_C#o_RR<=)7q7)85N8HsI8-0E4FR8IFM0R;j2
RRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMRFbsO#C#;R
RRMRC8CRoMNCs0zCR4
j;RRRRzR44:VRHRF5M0NRs8_8ss2CoRMoCC0sNCR
RRRRRRRRRRNRs8C_soR_#<)=Rq)77;R
RRMRC8CRoMNCs0zCR4
4;
RRRRR--Q5VRI8N8sC_sos2RC#oH0RCsq)77RHk#MBoRpRi
RzRR4R.R:VRHRN5I8_8ss2CoRMoCC0sNCR
RRRRRRsRbF#OC#BR5pRi,W7q7)L2RCMoH
RRRRRRRRRRRRRHV5iBpR'=R4N'RMB8RpCi'P0CM2ER0CRM
RRRRRRRRRRRRRIRRNs8_C#o_RR<=W7q7)85N8HsI8-0E4FR8IFM0R;j2
RRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMRFbsO#C#;R
RRMRC8CRoMNCs0zCR4
.;RRRRzR4d:VRHRF5M0NRI8_8ss2CoRMoCC0sNCR
RRRRRRRRRRNRI8C_soR_#<W=Rq)77;R
RRMRC8CRoMNCs0zCR4
d;RRRRRRRR
RRRRR--tCCMsCN0RC0ERv)qRDOCDN#RM#8RCODC0FRDo
HORRRRzR4c:FRVsRRHH5MRM_klODCD_Rnc-2R4RI8FMR0FjCRoMNCs0RC
R-RR-VRQR85N8HsI8R0E>2R6RCMC8FR0RCOsNR0CI0sHCMRCNCLDR8NMR0FkbRk0CLMND#CRCODC0FRDo
HORRRRRRRRzR46:VRHR85N8HsI8R0E>2RnRMoCC0sNCR
RRRRRRRRRRRRRRFRskC0_M5_#H<2R=4R''ERIC5MRs_N8s_Co#85N8HsI8-0E4FR8IFM0RRn2=2RHR#CDCjR''S;
SISSF_k0C#M_5RH2<'=R4I'RERCM58IN_osC_N#58I8sHE80-84RF0IMF2RnRH=R2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0C#M_5RH2<W=R ERIC5MRI_N8s_Co#85N8HsI8-0E4FR8IFM0RRn2=2RHR#CDCjR''R;
RRRRRCRRMo8RCsMCNR0Cz;46
RRRRR--Q5VRNs88I0H8E=R<RR62MIFRsCH0RNCMLRDCFFsRkk0b0MRCNCLDRD#CCRO0DHFoOCRMC88C
RRRRRRRRnz4RH:RVNR58I8sHE80RR<=no2RCsMCN
0CRRRRRRRRRRRRRRRRs0Fk__CM#25HRR<=';4'
SSSSkIF0M_C_H#52=R<R''4;R
RRRRRRRRRRRRRRsRI0M_C_H#52=R<R;W 
RRRRRRRR8CMRMoCC0sNC4RznR;
R-RR-CRtMNCs00CRE)CRqOvRC#DDR8NMRH0s-N#00
C#RRRRRRRRzR4(:FRVsRR[H5MRI0H8ERR-482RF0IMFRRjoCCMsCN0
RRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVzv)qn:cRRLDNCHDR#1R"7Ra"&MRH0CCosl'HN5oCI0H8E&2RR""7RH&RMo0CCHs'lCNo5nH*c&2RR""WRH&RMo0CCHs'lCNo5R[2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50E54H+2c*n,CR8b20E2RR&"RX"&MRH0CCosl'HN5oC[2+4;R
RRRRRRRRRRCRLo
HMRRRRRRRRRRRRzv)qn:cRRqX)vXnc4
7RRRRRRRRRRRRRRRRRb0FsRblNRR57=H>RMC_so5_#[R2,q=jR>FRDIN_I8_8s#25j,4RqRR=>D_FII8N8s5_#4R2,q=.R>FRDIN_I8_8s#25.,R
RRRRRRRRRRRRRRRRRRRRRRRRRq=dR>FRDIN_I8_8s#25d,cRqRR=>D_FII8N8s5_#cR2,q=6R>FRDIN_I8_8s#256,SR
SSSSS7RRuj)qRR=>D_FIs8N8s5_#jR2,7qu)4>R=RIDF_8sN8#s_5,42R)7uq=.R>FRDIN_s8_8s#25.,S
SSSSSRuR7)Rqd=D>RFsI_Ns88_d#527,Ruc)qRR=>D_FIs8N8s5_#cR2,7qu)6>R=RIDF_8sN8#s_5,62RS
SSSSSR RWRR=>I_s0C#M_5,H2RpWBi>R=RiBp,uR7m>R=RksF0k_L#c_n#,5H[R2,1Rum=I>RF_k0L_k#n5c#H2,[2R;
RRRRRRRRRRRRRsRRF_k0s_Co#25[RR<=s0Fk_#Lk_#nc5[H,2ERIC5MRs0Fk__CM#25HR'=R4R'2CCD#R''Z;S
SSFSIks0_C#o_5R[2<I=RF_k0L_k#n5c#H2,[RCIEMIR5F_k0C#M_5RH2=4R''C2RDR#C';Z'
RRRRRRRR8CMRMoCC0sNC4Rz(R;
RRRRCRM8oCCMsCN0Rcz4;RRRRRRRRRRRRR
RRRRR
RRRRR--tCCMsCN0RdNR.FRIs88RCRCb)RqvODCDRRHVNsbbFHbsNR0CRRRRRRRRRRRRRRR
RzRR4:URRRHV5lMk_DOCD._dR4=R2CRoMNCs0RC
R-RR-VRQR85N8HsI8R0E>2R(RCMC8FR0RCOsNR0CI0sHCMRCNCLDR8NMR0FkbRk0CLMND#CRCODC0FRDo
HORRRRRRRRzN4gRH:RVNR58I8sHE80Rn>R2CRoMNCs0RC
RRRRRRRRRRRRRsRRF_k0CdM_.=R<R''4RCIEM5R5s_N8s_Co#85N8HsI8-0E4FR8IFM0RRn2=kRMlC_ODnD_cN2RM58Rs_N8s_Co#256R'=Rj2'2R#CDCjR''S;
SISSF_k0CdM_.=R<R''4RCIEM5R5I_N8s_Co#85N8HsI8-0E4FR8IFM0RRn2=kRMlC_ODnD_cN2RM58RI_N8s_Co#256R'=Rj2'2R#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_M._dRR<=WI RERCM5N5I8C_so5_#Ns88I0H8ER-48MFI0nFR2RR=M_klODCD_2ncR8NMRN5I8C_so5_#6=2RR''j2C2RDR#C';j'
RRRRRRRR8CMRMoCC0sNC4Rzg
N;RRRRRRRRzL4gRH:RVNR58I8sHE80Rn=RR8NMRlMk_DOCDc_nRj=R2CRoMNCs0RC
RRRRRRRRRRRRRsRRF_k0CdM_.=R<R''4RCIEM5R5s_N8s_Co#256R'=Rj2'2R#CDCjR''S;
SISSF_k0CdM_.=R<R''4RCIEM5R5I_N8s_Co#256R'=Rj2'2R#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_M._dRR<=WI RERCM5N5I8C_so5_#6=2RR''j2C2RDR#C';j'
RRRRRRRR8CMRMoCC0sNC4RzgRL;R-RR-VRQR85N8HsI8R0E<6=R2FRMRHIs0CCRMDNLCsRFR0FkbRk0CLMND#CRCODC0FRDoRHOM8CCCR8
RRRRRzRR.:jRRRHV58N8s8IH0<ER=2R6RMoCC0sNCR
RRRRRRRRRRRRRRFRskC0_M._dRR<=';4'
SSSSkIF0M_C_Rd.<'=R4
';RRRRRRRRRRRRRRRRI_s0CdM_.=R<R;W 
RRRRRRRR8CMRMoCC0sNC.RzjR;
R-RR-CRtMNCs00CRE)CRqOvRCRDDNRM80-sH#00NCR
RRRRRR.Rz4RR:VRFs[MRHRH5I8R0E-2R4RI8FMR0FjCRoMNCs0RC
RRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)Rzq.vdRD:RNDLCRRH#"a17"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloMC5kOl_C_DDnnc*c&2RR""WRH&RMo0CCHs'lCNo5R[2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50EM_klODCD_*ncn+cRR,d.Rb8C02E2R"&RX&"RR0HMCsoC'NHlo[C5+;42
RRRRRRRRRRRRoLCHRM
RRRRRRRRRzRR)dqv.RR:Xv)qd4.X7RR
RRRRRRRRRRRRRbRRFRs0lRNb5=7R>MRH_osC_[#52q,Rj>R=RIDF_8IN8#s_5,j2RRq4=D>RFII_Ns88_4#52q,R.>R=RIDF_8IN8#s_5,.2
RRRRRRRRRRRRRRRRRRRRRRRRqRRd>R=RIDF_8IN8#s_5,d2RRqc=D>RFII_Ns88_c#52
,RSSSSSRSR7qu)j>R=RIDF_8sN8#s_5,j2R)7uq=4R>FRDIN_s8_8s#254,uR7)Rq.=D>RFsI_Ns88_.#52S,
SSSSS7RRud)qRR=>D_FIs8N8s5_#dR2,7qu)c>R=RIDF_8sN8#s_5,c2RS
SSSSSR RWRR=>I_s0CdM_.W,RBRpi=B>RpRi,7Rum=s>RF_k0L_k#d5.#M_klODCD_,d.[R2,1Rum=I>RF_k0L_k#d5.#M_klODCD_,d.[;22
RRRRRRRRRRRRRRRRksF0C_so5_#[<2R=FRskL0_kd#_.M#5kOl_C_DDd[.,2ERIC5MRs0Fk__CMd=.RR''42DRC#'CRZ
';SSSSI0Fk_osC_[#52=R<RkIF0k_L#._d#k5MlC_ODdD_.2,[RCIEMIR5F_k0CdM_.RR='24'R#CDCZR''R;
RRRRRRRRCRM8oCCMsCN0R4z.;R
RRCRRMo8RCsMCNR0Cz;4URRRRRRRRR
R
RRRR-t-RCsMCNR0CNnR4RsIF8CR8C)bRqOvRCRDDHNVRbFbsbNsH0RCRRRRRRRRRRRRRRR
RR.Rz.RR:H5VRM_klODCD_R4n=2R4RMoCC0sNCR
RR-R-RRQV58N8s8IH0>ERRR62M8CCRR0FONsC0ICRsCH0RNCMLRDCNRM8Fbk0kC0RMDNLCCR#D0CORoDFHRO
RRRRRzRR.RdN:VRHR85N8HsI8R0E>RRnNRM8M_klODCD_Rd.=2R4RMoCC0sNCR
RRRRRRRRRRRRRRFRskC0_Mn_4RR<='R4'IMECRs55Ns8_C#o_58N8s8IH04E-RI8FMR0Fn=2RRlMk_DOCDc_n2MRN8sR5Ns8_C#o_5R62=4R''N2RM58Rs_N8s_Co#25cR'=Rj2'2R#CDCjR''S;
SISSF_k0C4M_n=R<R''4RCIEM5R5I_N8s_Co#85N8HsI8-0E4FR8IFM0RRn2=kRMlC_ODnD_cN2RM58RI_N8s_Co#256R'=R4R'2NRM858IN_osC_c#52RR='2j'2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0C4M_n=R<RRW IMECRI55Ns8_C#o_58N8s8IH04E-RI8FMR0Fn=2RRlMk_DOCDc_n2MRN8IR5Ns8_C#o_5R62=4R''N2RM58RI_N8s_Co#25cR'=Rj2'2R#CDCjR''R;
RRRRRCRRMo8RCsMCNR0CzN.d;R
RRRRRR.Rzd:LRRRHV58N8s8IH0>ERRNnRMM8RkOl_C_DDd/.R=2R4RMoCC0sNCR
RRRRRRRRRRRRRRFRskC0_Mn_4RR<='R4'IMECRs55Ns8_C#o_58N8s8IH04E-RI8FMR0Fn=2RRlMk_DOCDc_n2MRN8sR5Ns8_C#o_5R62=jR''N2RM58Rs_N8s_Co#25cR'=Rj2'2R#CDCjR''S;
SISSF_k0C4M_n=R<R''4RCIEM5R5I_N8s_Co#85N8HsI8-0E4FR8IFM0RRn2=kRMlC_ODnD_cN2RM58RI_N8s_Co#256R'=RjR'2NRM858IN_osC_c#52RR='2j'2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0C4M_n=R<RRW IMECRI55Ns8_C#o_58N8s8IH04E-RI8FMR0Fn=2RRlMk_DOCDc_n2MRN8IR5Ns8_C#o_5R62=jR''N2RM58RI_N8s_Co#25cR'=Rj2'2R#CDCjR''R;
RRRRRCRRMo8RCsMCNR0CzL.d;R
RRRRRR.Rzd:ORRRHV58N8s8IH0=ERRNnRMM8RkOl_C_DDd=.RRR42oCCMsCN0
RRRRRRRRRRRRRRRRksF0M_C_R4n<'=R4I'RERCM5N5s8C_so5_#6=2RR''42MRN8sR5Ns8_C#o_5Rc2=jR''R22CCD#R''j;S
SSFSIkC0_Mn_4RR<='R4'IMECRI55Ns8_C#o_5R62=4R''N2RM58RI_N8s_Co#25cR'=Rj2'2R#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_Mn_4RR<=WI RERCM5N5I8C_so5_#6=2RR''42MRN8IR5Ns8_C#o_5Rc2=jR''R22CCD#R''j;R
RRRRRRMRC8CRoMNCs0zCR.;dO
RRRRRRRRdz.8RR:H5VRNs88I0H8ERR=6MRN8kRMlC_ODdD_.=R/RR42oCCMsCN0
RRRRRRRRRRRRRRRRksF0M_C_R4n<'=R4I'RERCM5N5s8C_so5_#Ns88I0H8ER-48MFI0cFR2RR=M_klODCD_2d.2DRC#'CRj
';SSSSI0Fk__CM4<nR=4R''ERIC5MR58IN_osC_N#58I8sHE80-84RF0IMF2RcRM=RkOl_C_DDd2.2R#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_Mn_4RR<=WI RERCM5N5I8C_so5_#Ns88I0H8ER-48MFI0cFR2RR=M_klODCD_2d.2DRC#'CRj
';RRRRRRRRCRM8oCCMsCN0Rdz.8R;RR-R-RRQV58N8s8IH0<ER=2R6RRMFI0sHCMRCNCLDRRFsFbk0kC0RMDNLCCR#D0CORoDFHMORCCC88R
RRRRRR.RzcRR:H5VRNs88I0H8E=R<RRc2oCCMsCN0
RRRRRRRRRRRRRRRRksF0M_C_R4n<'=R4
';SSSSI0Fk__CM4<nR=4R''R;
RRRRRRRRRRRRRIRRsC0_Mn_4RR<=W
 ;RRRRRRRRCRM8oCCMsCN0Rcz.;R
RR-R-RMtCC0sNCER0CqR)vCRODNDRM08Rs#H-0CN0
RRRRRRRR6z.RV:RF[sRRRHM58IH0-ERRR428MFI0jFRRMoCC0sNCR
RRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqz)vR4n:NRDLRCDH"#R1"7aRH&RMo0CCHs'lCNo58IH0RE2&7R""RR&HCM0o'CsHolNCk5MlC_ODnD_cc*nRM+RkOl_C_DDdd.*.&2RR""WRH&RMo0CCHs'lCNo5R[2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50EM_klODCD_*ncn+cRRlMk_DOCD._d*Rd.+nR4,CR8b20E2RR&"RX"&MRH0CCosl'HN5oC[2+4;R
RRRRRRRRRRCRLo
HMRRRRRRRRRRRRzv)q4:nRRv)q44nX7RR
RRRRRRRRRRRRRbRRFRs0lRNb5=7R>MRH_osC_[#52q,Rj>R=RIDF_8IN8#s_5,j2RRq4=D>RFII_Ns88_4#52q,R.>R=RIDF_8IN8#s_5,.2
RRRRRRRRRRRRRRRRRRRRRRRRqRRd>R=RIDF_8IN8#s_5,d2R)7uq=jR>FRDIN_s8_8s#25j,uR7)Rq4=D>RFsI_Ns88_4#527,Ru.)qRR=>D_FIs8N8s5_#.
2,SSSSSRSR7qu)d>R=RIDF_8sN8#s_5,d2RRW =I>RsC0_Mn_4,BRWp=iR>pRBi7,Ru=mR>FRskL0_k4#_nM#5kOl_C_DD4[n,21,Ru=mR>FRIkL0_k4#_nM#5kOl_C_DD4[n,2
2;RRRRRRRRRRRRRRRRs0Fk_osC_[#52=R<RksF0k_L#n_4#k5MlC_OD4D_n2,[RCIEMsR5F_k0C4M_nRR='24'R#CDCZR''S;
SISSF_k0s_Co#25[RR<=I0Fk_#Lk_#4n5lMk_DOCDn_4,R[2IMECRF5IkC0_Mn_4R'=R4R'2CCD#R''Z;R
RRRRRRMRC8CRoMNCs0zCR.
6;RRRRCRM8oCCMsCN0R.z.;RRRRR
RCRM8oCCMsCN0Rczc;M
C8sRNO0EHCkO0sLCRD	FO_lsN;-

---------------------M--FI_s_COEO-	----------------------
-
NEsOHO0C0CksR_MFsOI_E	CORRFV)_qv)_Wu)#RH
lOFbCFMMX0R)dqv.7X4RbRRFRs05R
RRRRRRuR7mRRR:kRF00R#8D_kFOoH;RRRRRRRRR
RRRRRRuR1mRRR:kRF00R#8D_kFOoH;R

RRRRRqRRjRRRRH:RM0R#8D_kFOoH;R
RRRRRR4RqRRRR:MRHR8#0_FkDo;HO
RRRRRRRRRq.R:RRRRHM#_08koDFH
O;RRRRRRRRqRdRRRR:H#MR0k8_DHFoOR;
RRRRRqRRcRRRRH:RM0R#8D_kFOoH;R
RRRRRRRR7RRRR:MRHR8#0_FkDo;HO
RRRRRRRR)7uq:jRRRHM#_08koDFH
O;RRRRRRRR7qu)4RR:H#MR0k8_DHFoOR;
RRRRR7RRu.)qRH:RM0R#8D_kFOoH;R
RRRRRRuR7)Rqd:MRHR8#0_FkDo;HO
RRRRRRRR)7uq:cRRRHM#_08koDFH
O;RRRRRRRRWiBpRRR:H#MR0k8_DHFoOR;RRRRRRRR
RRRRRWRR RRRRH:RM0R#8D_kFOoH
RRRRRRR2R;R
8CMRlOFbCFMM
0;ObFlFMMC0)RXqcvnXR47RFRbs50R
RRRRRRRRm7uR:RRR0FkR8#0_FkDo;HORRRRRRRR
RRRRRRRRm1uR:RRR0FkR8#0_FkDo;HO
R
RRRRRRjRqRRRR:MRHR8#0_FkDo;HO
RRRRRRRRRq4R:RRRRHM#_08koDFH
O;RRRRRRRRqR.RRRR:H#MR0k8_DHFoOR;
RRRRRqRRdRRRRH:RM0R#8D_kFOoH;R
RRRRRRcRqRRRR:MRHR8#0_FkDo;HO
RRRRRRRRRq6R:RRRRHM#_08koDFH
O;RRRRRRRR7RRRRRR:H#MR0k8_DHFoOR;
RRRRR7RRuj)qRH:RM0R#8D_kFOoH;R
RRRRRRuR7)Rq4:MRHR8#0_FkDo;HO
RRRRRRRR)7uq:.RRRHM#_08koDFH
O;RRRRRRRR7qu)dRR:H#MR0k8_DHFoOR;
RRRRR7RRuc)qRH:RM0R#8D_kFOoH;R
RRRRRRuR7)Rq6:MRHR8#0_FkDo;HO
RRRRRRRRpWBi:RRRRHM#_08koDFHRO;RRRRR
RRRRRRRRRRWR RRRR:H#MR0k8_DHFoOR
RRRRRRR2;RM
C8FROlMbFC;M0
MVkOF0HMkRVMHO_M5H0LRR:LDFFC2NMR0sCkRsM#H0sMHoR#C
Lo
HMRVRHR25LRC0EMR
RRCRs0Mks52"";R
RCCD#
RRRR0sCk5sM"kBFDM8RFH0RlCbDl0CMRFADO)	RqRv3Q0#REsCRCRN8Ns88CR##sHCo#s0CCk8R#oHMRC0ERl#NCDROFRO	N0#RE)CRq"v?2R;
R8CMR;HV
8CMRMVkOM_HH
0;VOkM0MHFR0oC_8CM_b8C0#E5HRxC:MRH0CCosRR;80CbERR:HCM0o2CsR0sCkRsMHCM0oRCsHP#
NNsHLRDCl_HM#CHxRH:RMo0CC:sR=;Rj
oLCHRM
RMlH_x#HC=R:Rb8C0
E;RVRHRH5#x<CRRb8C0RE20MEC
RRRRMlH_x#HC=R:Rx#HCR;
R8CMR;HV
sRRCs0kMHRlMH_#x
C;CRM8o_C0C_M880CbEN;
0H0sLCk0RMoCC0sNFss_CsbF0RR:#H0sM
o;Ns00H0LkCCRoMNCs0_FssFCbsF0RVFRM__sIOOEC	RR:NEsOHO0C0CksRRH#VOkM_HHM0N5s8_8ss2Co;-
-RoLCHLMRD	FORlsNRbHlDCClM00NHRFM#MHoN
D#0C$bR0HM_sNsNH$R#sRNsRN$50jRF2R6RRFVHCM0o;Cs
MOF#M0N0HRI8_0ENNss$RR:H_M0NNss$=R:R,54RR.,cg,R,UR4,nRd2O;
F0M#NRM080CbEs_NsRN$:MRH0s_NsRN$:5=R4UndcU,R4,g.Rgcjn.,Rj,cUR.4jc6,R4;.2
MOF#M0N0HR8PRd.:MRH0CCos=R:RH5I8-0E4d2/nO;
F0M#NRM084HPnRR:HCM0oRCs:5=RI0H8E2-4/;4U
MOF#M0N0HR8P:URR0HMCsoCRR:=58IH04E-2;/g
MOF#M0N0HR8P:cRR0HMCsoCRR:=58IH04E-2;/c
MOF#M0N0HR8P:.RR0HMCsoCRR:=58IH04E-2;/.
MOF#M0N0HR8P:4RR0HMCsoCRR:=58IH04E-2;/4
F
OMN#0ML0RF4FDRL:RFCFDN:MR=8R5HRP4>2Rj;F
OMN#0ML0RF.FDRL:RFCFDN:MR=8R5HRP.>2Rj;F
OMN#0ML0RFcFDRL:RFCFDN:MR=8R5HRPc>2Rj;F
OMN#0ML0RFUFDRL:RFCFDN:MR=8R5HRPU>2Rj;F
OMN#0ML0RF4FDnRR:LDFFCRNM:5=R84HPnRR>j
2;O#FM00NMRFLFDRd.:FRLFNDCM=R:RH58PRd.>2Rj;O

F0M#NRM084HPncdURH:RMo0CC:sR=8R5CEb0-/424UndcO;
F0M#NRM08UHP4Rg.:MRH0CCos=R:RC58b-0E4U2/4;g.
MOF#M0N0HR8PgcjnRR:HCM0oRCs:5=R80CbE2-4/gcjnO;
F0M#NRM08.HPjRcU:MRH0CCos=R:RC58b-0E4.2/j;cU
MOF#M0N0HR8P.4jcRR:HCM0oRCs:5=R80CbE2-4/.4jcO;
F0M#NRM086HP4:.RR0HMCsoCRR:=5b8C04E-24/6.
;
O#FM00NMRFLFD.64RL:RFCFDN:MR=8R5H4P6.RR>j
2;O#FM00NMRFLFD.4jcRR:LDFFCRNM:5=R84HPjR.c>2Rj;F
OMN#0ML0RF.FDjRcU:FRLFNDCM=R:RH58Pc.jURR>j
2;O#FM00NMRFLFDgcjnRR:LDFFCRNM:5=R8cHPjRgn>2Rj;F
OMN#0ML0RFUFD4Rg.:FRLFNDCM=R:RH58PgU4.RR>j
2;O#FM00NMRFLFDd4nU:cRRFLFDMCNRR:=5P8H4UndcRR>j
2;
MOF#M0N0kR#lH_I8R0E:MRH0CCos=R:RmAmph q'#bF5FLFDR42+mRAmqp hF'b#F5LF2D.RA+Rm mpqbh'FL#5FcFD2RR+Apmm 'qhb5F#LDFFU+2RRmAmph q'#bF5FLFD24n;F
OMN#0M#0Rk8l_CEb0RH:RMo0CC:sR=RR6-AR5m mpqbh'FL#5F6FD4R.2+mRAmqp hF'b#F5LFjD4.Rc2+mRAmqp hF'b#F5LFjD.cRU2+mRAmqp hF'b#F5LFjDcgRn2+mRAmqp hF'b#F5LF4DUg2.2;O

F0M#NRM0IE_OFCHO_8IH0:ERR0HMCsoCRR:=I0H8Es_Ns5N$#_klI0H8E
2;O#FM00NMROI_EOFHCC_8bR0E:MRH0CCos=R:Rb8C0NE_s$sN5l#k_8IH0;E2
MOF#M0N0_R8OHEFOIC_HE80RH:RMo0CC:sR=HRI8_0ENNss$k5#lC_8b20E;F
OMN#0M80R_FOEH_OC80CbERR:HCM0oRCs:8=RCEb0_sNsN#$5k8l_CEb02
;
O#FM00NMRII_HE80_lMk_DOCD:#RR0HMCsoCRR:=58IH04E-2_/IOHEFOIC_HE80R4+R;F
OMN#0MI0R_b8C0ME_kOl_C#DDRH:RMo0CC:sR=8R5CEb0-/42IE_OFCHO_b8C0+ERR
4;
MOF#M0N0_R8I0H8Ek_MlC_ODRD#:MRH0CCos=R:RH5I8-0E482/_FOEH_OCI0H8ERR+4O;
F0M#NRM08C_8b_0EM_klODCD#RR:HCM0oRCs:5=R80CbE2-4/O8_EOFHCC_8bR0E+;R4
F
OMN#0MI0R_x#HCRR:HCM0oRCs:I=R_8IH0ME_kOl_C#DDRI*R_b8C0ME_kOl_C#DD;F
OMN#0M80R_x#HCRR:HCM0oRCs:8=R_8IH0ME_kOl_C#DDR8*R_b8C0ME_kOl_C#DD;O

F0M#NRM0LDFF_:8RRFLFDMCNRR:=5#8_HRxC-_RI#CHxRR<=j
2;O#FM00NMRFLFDR_I:FRLFNDCM=R:R0MF5FLFD2_8;O

F0M#NRM0OHEFOIC_HE80RH:RMo0CC:sR=AR5m mpqbh'FL#5F_FD8*2RRO8_EOFHCH_I820ER5+RApmm 'qhb5F#LDFF_RI2*_RIOHEFOIC_HE802O;
F0M#NRM0OHEFO8C_CEb0RH:RMo0CC:sR=AR5m mpqbh'FL#5F_FD8*2RRO8_EOFHCC_8b20ER5+RApmm 'qhb5F#LDFF_RI2*_RIOHEFO8C_CEb02O;
F0M#NRM0I0H8Ek_MlC_ODRD#:MRH0CCos=R:Rm5Amqp hF'b#F5LF8D_25R*I0H8E2-4/O8_EOFHCH_I820ER5+RApmm 'qhb5F#LDFF_RI2*IR5HE80-/42IE_OFCHO_8IH0RE2+;R4
MOF#M0N0CR8b_0EM_klODCD#RR:HCM0oRCs:5=RApmm 'qhb5F#LDFF_R82*C58b-0E482/_FOEH_OC80CbE+2RRm5Amqp hF'b#F5LFID_2RR*5b8C04E-2_/IOHEFO8C_CEb02RR+40;
$RbCF_k0L4k#_b0$C#RHRsNsN5$R80CbEk_MlC_OD-D#4FR8IFM0RRj,I0H8Ek_MlC_OD-D#4FR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNRksF0k_L#:4RR0Fk_#Lk4$_0bRC;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RV_Rs80FkRM5HbRk000FRs#H-0CN0##2
HNoMDFRIkL0_kR#4:kRF0k_L#04_$;bC
b0$CkRF0k_L#0._$RbCHN#Rs$sNRC58b_0EM_klODCD#R-48MFI0jFR,*R.I0H8Ek_MlC_OD+D#4FR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNRksF0k_L#:.RR0Fk_#Lk.$_0bRC;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RV_Rs80FkRM5HbRk000FRs#H-0CN0##2
HNoMDFRIkL0_kR#.:kRF0k_L#0._$;bC
b0$CkRF0k_L#0c_$RbCHN#Rs$sNRC58b_0EM_klODCD#R-48MFI0jFR,*RcI0H8Ek_MlC_OD+D#dFR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNRksF0k_L#:cRR0Fk_#Lkc$_0bRC;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RV_Rs80FkRM5HbRk000FRs#H-0CN0##2
HNoMDFRIkL0_kR#c:kRF0k_L#0c_$;bC
b0$CkRF0k_L#0U_$RbCHN#Rs$sNRC58b_0EM_klODCD#R-48MFI0jFR,*RUI0H8Ek_MlC_OD+D#(FR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNRksF0k_L#:URR0Fk_#LkU$_0bRC;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RV_Rs80FkRM5HbRk000FRs#H-0CN0##2
HNoMDFRIkL0_kR#U:kRF0k_L#0U_$;bC
b0$CNRbs$H0_#LkU$_0bHCR#sRNsRN$5b8C0ME_kOl_C#DD-84RF0IMF,RjR8IH0ME_kOl_C#DD-84RF0IMF2RjRRFV#_08DHFoO#;
HNoMDbRsN0sH$k_L#:URRsbNH_0$LUk#_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$FsVR_k8F0HR5M0bkRR0F0-sH#00NC
#2#MHoNIDRbHNs0L$_kR#U:NRbs$H0_#LkU$_0b
C;0C$bR0Fk_#Lk40n_$RbCHN#Rs$sNRC58b_0EM_klODCD#R-48MFI0jFR,nR4*8IH0ME_kOl_C#DD+R468MFI0jFR2VRFR8#0_oDFH
O;#MHoNsDRF_k0L4k#nRR:F_k0L4k#n$_0bRC;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RV_Rs80FkRM5HbRk000FRs#H-0CN0##2
HNoMDFRIkL0_kn#4RF:RkL0_kn#4_b0$C0;
$RbCbHNs0L$_kn#4_b0$C#RHRsNsN5$R80CbEk_MlC_OD-D#4FR8IFM0RRj,.H*I8_0EM_klODCD#R+48MFI0jFR2VRFR8#0_oDFH
O;#MHoNsDRbHNs0L$_kn#4Rb:RN0sH$k_L#_4n0C$b;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFVsF_8k50RHkMb0FR0RH0s-N#002C#
o#HMRNDIsbNH_0$L4k#nRR:bHNs0L$_kn#4_b0$C0;
$RbCF_k0Ldk#.$_0bHCR#sRNsRN$5b8C0ME_kOl_C#DD-84RF0IMF,RjR*d.I0H8Ek_MlC_OD+D#d84RF0IMF2RjRRFV#_08DHFoO#;
HNoMDFRskL0_k.#dRF:RkL0_k.#d_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFR8s_FRk05bHMk00RFsR0H0-#N#0C2H
#oDMNRkIF0k_L#Rd.:kRF0k_L#_d.0C$b;$
0bbCRN0sH$k_L#_d.0C$bRRH#NNss$8R5CEb0_lMk_DOCD4#-RI8FMR0Fjc,R*8IH0ME_kOl_C#DD+8dRF0IMF2RjRRFV#_08DHFoO#;
HNoMDbRsN0sH$k_L#Rd.:NRbs$H0_#Lkd0._$;bCRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$FsVR_k8F0HR5M0bkRR0F0-sH#00NC
#2#MHoNIDRbHNs0L$_k.#dRb:RN0sH$k_L#_d.0C$b;H
#oDMNRksF0M_CR#:R0D8_FOoH_OPC05Fs80CbEk_MlC_OD-D#4FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--CLMNDRC#VRFs0-sH#00NC##
HNoMDFRIkC0_MRR:#_08DHFoOC_POs0F5b8C0ME_kOl_C#DD-84RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RNCML#DCRsVFRH0s-N#00
C##MHoNIDRsC0_MRR:#_08DHFoOC_POs0F5b8C0ME_kOl_C#DD-84RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RHIs0CCRMDNLCV#RFCsRNROEsRFIF)VRqOvRC#DD
o#HMRNDHsM_C:oRR8#0_oDFHPO_CFO0sH5I8+0Ed86RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-k-R#RC80sFRC#oH0RCs7RQh
o#HMRNDs0Fk_osCR#:R0D8_FOoH_OPC05FsI0H8E6+dRI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--k8#CRR0FsHCo#s0CRz7maH
#oDMNRkIF0C_soRR:#_08DHFoOC_POs0F58IH0dE+6FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RCk#8FR0RosCHC#0smR7z#a
HNoMDFRsks0_CRo4:0R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RCk#8FR0RFOEFR#CLIC0CRCM7RQhNRM8Fbk0kF0RVDRAFRO	)
qv#MHoNsDRNs8_C:oRR8#0_oDFHPO_CFO0s85N8HsI8-0E4FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-#RkC08RFCRso0H#C)sRq)77
o#HMRNDI_N8sRCo:0R#8F_Do_HOP0COFNs58I8sHE80-84RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-k-R#RC80sFRC#oH0RCsW7q7)H
#oDMNRIDF_8sN8:sRR8#0_oDFHPO_CFO0sd54RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-R8sN8LsRHR0#HkMb0FR0Rv)qRDOCD5#RcHRL0s#RCHJks2C8
o#HMRNDD_FII8N8sRR:#_08DHFoOC_POs0F5R4d8MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--I8N8sHRL0H#RM0bkRR0F)RqvODCD#cR5R0LH#CRsJskHC
82#MHoN)DRq)77_b0lR#:R0D8_FOoH_OPC05FsNs88I0H8ER-48MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--k8#CRR0FbCHbDCHMR7)q7#)
HNoMDqRW7_7)0Rlb:0R#8F_Do_HOP0COFNs58I8sHE80-84RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-k-R#RC80bFRHDbCHRMCW7q7)H
#oDMNRh7Q_b0lR#:R0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-#RkC08RFHRbbHCDM7CRQ#h
HNoMD RW_b0lR#:R0D8_FOoH;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-k-R#RC80bFRHDbCHRMCW# 
HNoMD_RsNs88_osCR#:R0D8_FOoH_OPC05FsNs88I0H8ER-48MFI0jFR2-;
-MRC8DRLFRO	sRNlHDlbCMlC0HN0F#MRHNoMD-#
-CRLoRHM#CCDOs0RNHlRlCbDl0CMNF0HMHR#oDMN#k
VMHO0FoMRCM0_knl_cC58b:0ER0HMCsoC2CRs0MksR0HMCsoCR
H#PHNsNCLDRDPNRH:RMo0CC:sR=;Rj
oLCHRM
RDPNRR:=80CbEc/n;R
RH5VR5b8C0lERFn8Rc>2RR2cURC0EMR
RRNRPD=R:RDPNR4+R;R
RCRM8H
V;RCRs0MksRDPN;M
C8CRo0k_Mlc_n;k
VMHO0FoMRCD0_CFV0P_Csd8.5CEb0RH:RMo0CCRs2skC0sHMRMo0CCHsR#C
Lo
HMRCRs0Mks5b8C0lERFn8Rc
2;CRM8o_C0D0CVFsPC_;d.
MVkOF0HMCRo0C_DVP0FC8s5CEb0RH:RMo0CCRs;lRNG:MRH0CCoss2RCs0kMMRH0CCos#RH
sPNHDNLCNRPDRR:HCM0oRCs:j=R;C
Lo
HMRVRHRC58bR0E-NRlG=R>RRj20MEC
RRRRDPNRR:=80CbERR-l;NG
CRRD
#CRRRRPRND:8=RCEb0;R
RCRM8H
V;RCRs0Mks5DPN2C;
Mo8RCD0_CFV0P;Cs
MVkOF0HMCRo0k_Ml._d5b8C0:ERR0HMCsoC2CRs0MksR0HMCsoCR
H#PHNsNCLDRDPNRH:RMo0CC:sR=;Rj
oLCHRM
RRHV5b8C0<ER=URcR8NMRb8C0>ERR24nRC0EMR
RRPRRN:DR=;R4
CRRMH8RVR;
R0sCkRsMP;ND
8CMR0oC_lMk_;d.
MVkOF0HMCRo0k_Mln_45b8C0:ERR0HMCsoC2CRs0MksR0HMCsoCR
H#PHNsNCLDRDPNRH:RMo0CC:sR=;Rj
oLCHRM
RRHV5b8C0<ER=nR4R8NMRb8C0>ERRRj20MEC
RRRRNRPD=R:R
4;RMRC8VRH;R
RskC0sPMRN
D;CRM8o_C0M_kl4
n;O#FM00NMRlMk_DOCDc_nRH:RMo0CC:sR=CRo0k_Mlc_n5b8C0;E2
MOF#M0N0CRDVP0FCds_.RR:HCM0oRCs:o=RCD0_CFV0P_Csd8.5CEb02O;
F0M#NRM0M_klODCD_Rd.:MRH0CCos=R:R0oC_lMk_5d.D0CVFsPC_2d.;F
OMN#0MD0RCFV0P_Cs4:nRR0HMCsoCRR:=o_C0D0CVFsPC5VDC0CFPs._d,.Rd2O;
F0M#NRM0M_klODCD_R4n:MRH0CCos=R:R0oC_lMk_54nD0CVFsPC_24n;0

$RbCF_k0L_k#0C$b_#ncRRH#NNss$MR5kOl_C_DDn8cRF0IMF,RjR8IH04E-RI8FMR0FjF2RV0R#8F_Do;HO
b0$CkRF0k_L#$_0bdC_.H#R#sRNsRN$5lMk_DOCD._dRI8FMR0FjI,RHE80-84RF0IMF2RjRRFV#_08DHFoO0;
$RbCF_k0L_k#0C$b_#4nRRH#NNss$MR5kOl_C_DD48nRF0IMF,RjR8IH04E-RI8FMR0FjF2RV0R#8F_Do;HO
o#HMRNDs0Fk_#Lk_#ncRF:RkL0_k0#_$_bCn;c#RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$F8VRFRk05bHMk00RFsR0H0-#N#0C2H
#oDMNRkIF0k_L#c_n#RR:F_k0L_k#0C$b_#nc;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFV80FkRM5HbRk000FRs#H-0CN0##2
HNoMDFRskL0_kd#_.:#RR0Fk_#Lk_b0$C._d#R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFRk8F0HR5M0bkRR0F0-sH#00NC
#2#MHoNIDRF_k0L_k#dR.#:kRF0k_L#$_0bdC_.
#;#MHoNsDRF_k0L_k#4Rn#:kRF0k_L#$_0b4C_nR#;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RVFR8k50RHkMb0FR0RH0s-N#002C#
o#HMRNDI0Fk_#Lk_#4nRF:RkL0_k0#_$_bC4;n#
o#HMRNDs0Fk__CM#RR:#_08DHFoOC_POs0F5lMk_DOCDc_nRI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-C-RMDNLCV#RF0sRs#H-0CN0#H
#oDMNRkIF0M_C_:#RR8#0_oDFHPO_CFO0sk5MlC_ODnD_cFR8IFM0R;j2
o#HMRNDs0Fk__CMd:.RR8#0_oDFH
O;#MHoNIDRF_k0CdM_.RR:#_08DHFoO#;
HNoMDFRskC0_Mn_4R#:R0D8_FOoH;H
#oDMNRkIF0M_C_R4n:0R#8F_Do;HO
o#HMRNDI_s0C#M_R#:R0D8_FOoH_OPC05FsM_klODCD_Rnc8MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-sRIHR0CCLMNDRC#VRFsCENORIsFRRFV)RqvODCD#H
#oDMNR0Is__CMd:.RR8#0_oDFH
O;#MHoNIDRsC0_Mn_4R#:R0D8_FOoH;H
#oDMNR_HMs_Co#RR:#_08DHFoOC_POs0F58IH04E-RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RCk#8FR0RosCHC#0sQR7h#R
HNoMDFRsks0_C#o_R#:R0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-k-R#RC80sFRC#oH0RCs7amz
o#HMRNDI0Fk_osC_:#RR8#0_oDFHPO_CFO0sH5I8-0E4FR8IFM0R;j2R
RR#MHoNsDRNs8_C#o_R#:R0D8_FOoH_OPC05FsNs88I0H8ER-48MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--k8#CRR0FsHCo#s0CR7q7)H
#oDMNR8IN_osC_:#RR8#0_oDFHPO_CFO0s85N8HsI8-0E4FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-#RkC08RFCRso0H#CqsR7
7)#MHoNDDRFsI_Ns88_:#RR8#0_oDFHPO_CFO0sR568MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--Ns88R0LH#MRHbRk00)FRqOvRC#DDRR5cL#H0RJsCkCHs8#2
HNoMDFRDIN_I8_8s#RR:#_08DHFoOC_POs0F586RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-N-R8R8sL#H0RbHMk00RFqR)vCRODRD#5LcRHR0#skCJH8sC2-
-R8CMRD#CCRO0sRNlHDlbCMlC0HN0F#MRHNoMDN#
0H0sLCk0Rs\3NFl_VCV#0:\RRs#0H;Mo
C
Lo
HMRcRzdH:RVsR5Ns88_osC2CRoMNCs0-CR-CRoMNCs0LCRD	FORlsN
RRRRR--QNVR8I8sHE80RO<REOFHCH_I8R0ENH##o'MRj0'RFMRkk8#CR0LH#R
RRjRzRRR:H5VRNs88I0H8ERR=4o2RCsMCN
0CSRRRRIDF_8sN8<sR=jR"jjjjjjjjjjjj"RR&s_N8s5Coj
2;SRRRRIDF_8IN8<sR=jR"jjjjjjjjjjjj"RR&I_N8s5Coj
2;S8CMRMoCC0sNCjRz;R
RR4RzRRR:H5VRNs88I0H8ERR=.o2RCsMCN
0CSFSDIN_s8R8s<"=Rjjjjjjjjjjjj"RR&s_N8s5Co4FR8IFM0R;j2
RSRRFRDIN_I8R8s<"=Rjjjjjjjjjjjj"RR&I_N8s5Co4FR8IFM0R;j2
MSC8CRoMNCs0zCR4R;
RzRR.:RRRRHV58N8s8IH0=ERRRd2oCCMsCN0
DSSFsI_Ns88RR<="jjjjjjjjjjj"RR&s_N8s5Co.FR8IFM0R;j2
RSRRFRDIN_I8R8s<"=Rjjjjjjjjj"jjRI&RNs8_C.o5RI8FMR0Fj
2;S8CMRMoCC0sNC.Rz;R
RRdRzRRR:H5VRNs88I0H8ERR=co2RCsMCN
0CSFSDIN_s8R8s<"=RjjjjjjjjjRj"&NRs8C_soR5d8MFI0jFR2S;
RRRRD_FII8N8s=R<Rj"jjjjjjjjj"RR&I_N8s5CodFR8IFM0R;j2
MSC8CRoMNCs0zCRdR;
RzRRc:RRRRHV58N8s8IH0=ERRR62oCCMsCN0
RSRRFRDIN_s8R8s<"=Rjjjjjjjjj&"RR8sN_osC58cRF0IMF2Rj;R
SRDRRFII_Ns88RR<="jjjjjjjjRj"&NRI8C_soR5c8MFI0jFR2S;
CRM8oCCMsCN0R;zc
RRRRRz6RH:RVNR58I8sHE80Rn=R2CRoMNCs0SC
RRRRD_FIs8N8s=R<Rj"jjjjjjRj"&NRs8C_soR568MFI0jFR2S;
SIDF_8IN8<sR=jR"jjjjj"jjRI&RNs8_C6o5RI8FMR0Fj
2;S8CMRMoCC0sNC6Rz;R
RRnRzRRR:H5VRNs88I0H8ERR=(o2RCsMCN
0CSRRRRIDF_8sN8<sR=jR"jjjjjRj"&NRs8C_soR5n8MFI0jFR2S;
SIDF_8IN8<sR=jR"jjjjjRj"&NRI8C_soR5n8MFI0jFR2S;
CRM8oCCMsCN0R;zn
RRRRRz(RH:RVNR58I8sHE80RU=R2CRoMNCs0SC
RRRRD_FIs8N8s=R<Rj"jjjjj"RR&s_N8s5Co(FR8IFM0R;j2
DSSFII_Ns88RR<="jjjj"jjRI&RNs8_C(o5RI8FMR0Fj
2;S8CMRMoCC0sNC(Rz;R
RRURzRRR:H5VRNs88I0H8ERR=go2RCsMCN
0CSRRRRIDF_8sN8<sR=jR"jjjj"RR&s_N8s5CoUFR8IFM0R;j2
DSSFII_Ns88RR<="jjjjRj"&NRI8C_soR5U8MFI0jFR2S;
CRM8oCCMsCN0R;zU
RRRRRzgRH:RVNR58I8sHE80R4=Rjo2RCsMCN
0CSRRRRIDF_8sN8<sR=jR"j"jjRs&RNs8_Cgo5RI8FMR0Fj
2;SFSDIN_I8R8s<"=Rjjjj"RR&I_N8s5CogFR8IFM0R;j2
MSC8CRoMNCs0zCRgR;
RzRR4RjR:VRHR85N8HsI8R0E=4R42CRoMNCs0SC
RRRRD_FIs8N8s=R<Rj"jj&"RR8sN_osC5R4j8MFI0jFR2S;
SIDF_8IN8<sR=jR"jRj"&NRI8C_soj54RI8FMR0Fj
2;S8CMRMoCC0sNC4RzjR;
RzRR4R4R:VRHR85N8HsI8R0E=.R42CRoMNCs0SC
RRRRD_FIs8N8s=R<Rj"j"RR&s_N8s5Co484RF0IMF2Rj;S
SD_FII8N8s=R<Rj"j"RR&I_N8s5Co484RF0IMF2Rj;C
SMo8RCsMCNR0Cz;44
RRRR.z4RRR:H5VRNs88I0H8ERR=4Rd2oCCMsCN0
RSRRFRDIN_s8R8s<'=Rj&'RR8sN_osC5R4.8MFI0jFR2S;
SIDF_8IN8<sR=jR''RR&I_N8s5Co48.RF0IMF2Rj;C
SMo8RCsMCNR0Cz;4.
RRRRdz4RRR:H5VRNs88I0H8ERR>4Rd2oCCMsCN0
RSRRFRDIN_s8R8s<s=RNs8_C4o5dFR8IFM0R;j2
RSRRFRDIN_I8R8s<I=RNs8_C4o5dFR8IFM0R;j2
MSC8CRoMNCs0zCR4
d;
RRRRR--Q5VR8_HMs2CoRosCHC#0sQR7h#RkHRMoB
piRRRRzR4cRH:RV8R5HsM_CRo2oCCMsCN0
RRRRRRRRFbsO#C#Rp5Bi7,RQRh2LHCoMR
RRRRRRRRRRVRHRp5BiRR='R4'NRM8B'piCMPC002RE
CMRRRRRRRRRRRRRRRRHsM_C<oR="R5jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"RR&72Qh;R
RRRRRRRRRRMRC8VRH;R
RRRRRRMRC8sRbF#OC#S;
CRM8oCCMsCN0Rcz4;R
RR4Rz6:RRRRHV50MFRM8H_osC2CRoMNCs0RC
RRRRRRRRRHRRMC_so=R<Rj5"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jjR7&RQ;h2
MSC8CRoMNCs0zCR4
6;
RRRRR--Q5VRsk8F0C_sos2RC#oH0RCs)m_7zkaR#oHMRm)_B
piRRRRzs4n80FkRRR:H5VRsk8F0C_soo2RCsMCN
0CRRRRRRRRbOsFCR##5m)_B,piRksF0C_soR42LHCoMR
RRRRRRRRRRVRHR_5)miBpR'=R4N'RM)8R_pmBiP'CC2M0RC0EMR
RRRRRRRRRRRRRR_R)7amzRR<=s0Fk_osC4R;
RRRRRRRRRCRRMH8RVR;
RRRRRCRRMb8RsCFO#
#;RRRRRRRRCRM8oCCMsCN0Rnz4sk8F0R;
RzRR48(sFRk0RH:RVMR5Fs0R80Fk_osC2CRoMNCs0RC
RRRRRRRRR)RR_z7ma=R<RksF0C_so
4;S8CMRMoCC0sNC4Rz(Fs8k
0;
4SznFI8kR0R:VRHR85IF_k0s2CoRMoCC0sNCR
RRRRRRsRbF#OC#WR5_pmBiI,RF_k0s2CoRoLCHRM
RRRRRRRRRHRRVWR5_pmBiRR='R4'NRM8WB_mpCi'P0CM2ER0CRM
RRRRRRRRRRRRRWRR_z7ma=R<RkIF0C_soH5I8-0E4FR8IFM0R;j2
RRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMRFbsO#C#;R
RRRRRRMRC8CRoMNCs0zCR48nIF;k0
RRRR(z4Ik8F0:RRRRHV50MFRFI8ks0_CRo2oCCMsCN0
RRRRRRRRRRRR7W_mRza<I=RF_k0s5CoI0H8ER-48MFI0jFR2S;
CRM8oCCMsCN0R(z4Ik8F0
;
RRRR-Q-RVsR5Ns88_osC2CRso0H#C)sRq)77RHk#MmoRB
piRRRRzs4nRRR:H5VRs8N8sC_soo2RCsMCN
0C-R-RRRRRRsRbF#OC#mR5B,piR7)q7R)2LHCoM-
-RRRRRRRRRRRRH5VRmiBpR'=R4N'RMm8RB'piCMPC002RE
CM-R-RRRRRRRRRRRRRRNRs8C_so=R<R7)q7N)58I8sHE80-84RF0IMF2Rj;-
-RRRRRRRRRRRRCRM8H
V;-R-RRRRRRMRC8sRbF#OC#-;
-MSC8CRoMNCs0zCR4;ns
R--RzRR4R(s:VRHRF5M0NRs8_8ss2CoRMoCC0sNCR
RRRRRRRRRRNRs8C_so=R<R7)q7
);S8CMRMoCC0sNC4Rzn
s;
-S-RRQV58IN8ss_CRo2sHCo#s0CR7Wq7k)R#oHMRmW_B
piRRRRzI4nRRR:H5VRI8N8sC_soo2RCsMCN
0CRRRRRRRRbOsFCR##5iBp,qRW727)RoLCHRM
RRRRRRRRRHRRVBR5p=iRR''4R8NMRiBp'CCPMR020MEC
RRRRRRRRRRRRRRRR8IN_osCRR<=W7q7)85N8HsI8-0E4FR8IFM0R;j2
RRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMRFbsO#C#;C
SMo8RCsMCNR0CzI4n;R
RR4Rz(:IRRRHV50MFR8IN8ss_CRo2oCCMsCN0
RRRRRRRRRRRR8IN_osCRR<=W7q7)S;
CRM8oCCMsCN0R(z4I
;
RRRR- -RGN0sRoDFHVORF7sRkRNDb0FsR#ONC-
S-0MFRCMC8RC8VRFsMsF_IE_OC
O	Sz--sRCo:sRbF#OC#p5BiL2RCMoH
S--RVRHRp5Bie'  RhaNRM8BRpi=4R''02RE
CM-R-SRQR7hl_0b=R<Rh7Q;-
-SRRR)7q7)l_0b=R<R7)q7
);-R-SRqRW7_7)0Rlb<W=Rq)77;-
-SRRRW0 _l<bR= RW;-
-SCRRMH8RV-;
-MSC8sRbF#OC#
;
SR--Q)VRCRN8qs88CR##=sRWHR0Cqs88C,##RbL$NR##7RQh0FFRkk0b0VRHRRW HC#RMDNLCS8
zGlkRb:RsCFO#W#5 l_0b),Rq)77_b0l,qRW7_7)0,lbRh7Q_b0l,FRsks0_C
o2SLRRCMoH
S--RRRRH5VRW7q7)l_0bRR=)7q7)l_0bMRN8 RW_b0lR'=R4R'20MEC
S--SsRRF_k0s4CoRR<=7_Qh0;lb
S--S#CDCS
SRFRsks0_CRo4<s=RF_k0s5CoI0H8ER-48MFI0jFR2-;
-CSSMH8RVS;
CRM8bOsFC;##
RSRRRR
R-RR-CRtMNCs00CRE)CRqOvRC#DDR8NMRD#CCRO0DHFoOFRVsqR)vnA4__141S4
zR4U:VRHRE5OFCHO_8IH0=ERRR42oCCMsCN0
RSRSRRRz	OE:VRHR85N8HsI8R0E>cR42CRoMNCs0RC
RRRRRkRRORD	:sRbF#OC#p5BiR2
RRRRRRRRLHCoMR
RRRRRRRRRH5VRB'piCMPC0MRN8pRBiRR='24'RC0EMR
RRRRRRRRRR_RsNs88_osC58N8s8IH04E-RI8FMR0F4Rc2<)=Rq)7758N8s8IH04E-RI8FMR0F4;c2
RRRRRRRRCRRMH8RVR;
RRRRRCRRMb8RsCFO#k#RO;D	
RSRCRM8oCCMsCN0REzO	R;
RSRRzR4g:FRVsRRHH5MR80CbEk_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0SC
-Q-RVNR58I8sHE80R4>RcM2RCRC80OFRs0CNCsRIHR0CCLMNDNCRMF8Rkk0b0MRCNCLDRD#CCRO0DHFoOR
RRRRRRzRS.:jRRRHV58N8s8IH0>ERR24cRMoCC0sNC-
S-HRVGFRVsNROD4DRd(UU,CR#D0CORRFV0#sH0CN0R0MFRHLCMsoRC#oH0CCs8S
SSFSskC0_M25HRR<='R4'IMECR_5sNs88_osC58N8s8IH04E-RI8FMR0F4Rc2=2RHR#CDCjR''S;
SISSF_k0CHM52=R<R''4RCIEMIR5Ns8_CNo58I8sHE80-84RF0IMFcR42RR=HC2RDR#C';j'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RWRCIEMIR5Ns8_CNo58I8sHE80-84RF0IMFcR42RR=HC2RDR#C';j'
RRRRRRRRMSC8CRoMNCs0zCR.
j;SR--Q5VRNs88I0H8E=R<R24cRRMFI0sHCMRCNCLDRRFsFbk0kC0RMDNLCCR#D0CORoDFHMORCCC88S
RRRRRS4z.RH:RVNR58I8sHE80RR<=4Rc2oCCMsCN0
SSSSksF0M_C5RH2<'=R4
';SSSSI0Fk_5CMH<2R=4R''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=W
 ;RRRRRRRRS8CMRMoCC0sNC.Rz4S;
-t-RCsMCNR0C0REC)RqvODCD#MRN8sR0H0-#N#0C
RRRRRRRR.Sz.RR:VRFs[MRHRH5I8_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
RRRRRRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVAv)q_d4nU4cX7RR:DCNLD#RHR""W;R
RRRRRRRRRRRRRRCRLo
HMRRRRRRRRRRRRSqA)vn_4dXUc4:7RRv)qA_4n114_4R
SRRRRRRRRRbRRFRs0lRNb5q7Q5Rj2=H>RMC_so25[,7Rq7R)q=D>RFII_Ns885R4d8MFI0jFR27,RQ=AR>jR""q,R7A7)RR=>D_FIs8N8sd54RI8FMR0Fj
2,SSSS Rhq='>R4R',1q1)RR=>',j'RqW RR=>I_s0CHM52B,RpRiq=B>RpRi, RhA='>R4R',1A1)RR=>',j'RAW RR=>',j'RiBpA>R=RiBp,S
SSRRRRq7m5Rj2=I>RF_k0L4k#5[H,27,RmjA52>R=RksF0k_L#H45,2[2;R

RRRRRRRRRRRRRsRRF_k0s5Co[<2R=FRskL0_k5#4H2,[RCIEMsR5F_k0CHM52RR='24'R#CDCZR''S;
SISSF_k0s5Co[<2R=FRIkL0_k5#4H2,KRCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRSRRCRM8oCCMsCN0R.z.;R
RRSRRCRM8oCCMsCN0Rgz4;R
RRMRC8CRoMNCs0zCR4RU;R
RRRRRRRRR
R-RR-CRtMNCs00CRE)CRqOvRC#DDR8NMRD#CCRO0DHFoOFRVsqR)vnA4__1.1S.
zR.d:VRHRE5OFCHO_8IH0=ERRR.2oCCMsCN0
RSRz	OERH:RVNR58I8sHE80R4>Rdo2RCsMCN
0CRRRRRRRRk	ODRb:RsCFO#B#5p
i2RRRRRRRRRoLCHRM
RRRRRRRRRRHV5iBp'CCPMN0RMB8Rp=iRR''42ER0CRM
RRRRRRRRRsRR_8N8sC_so85N8HsI8-0E4FR8IFM0R24dRR<=)7q7)85N8HsI8-0E4FR8IFM0R24d;R
RRRRRRRRRCRM8H
V;RRRRRRRRCRM8bOsFCR##k	OD;R
SR8CMRMoCC0sNCORzE
	;RRRRScz.RV:RFHsRRRHM5b8C0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CSR--Q5VRNs88I0H8ERR>4Rd2M8CCRR0FONsC0ICRsCH0RNCMLRDCNRM8Fbk0kC0RMDNLCCR#D0CORoDFHRO
RRRRRSRRzR.6:VRHR85N8HsI8R0E>dR42CRoMNCs0SC
-V-RHVGRFOsRNRDD4UdU(#,RCODC0VRFRH0s#00NCFRM0CRLHRMosHCo#s0CCR8
RRRRRRRRRRRRRsRRF_k0CHM52=R<R''4RCIEMsR5_8N8sC_so85N8HsI8-0E4FR8IFM0R24dRH=R2DRC#'CRj
';SSSSI0Fk_5CMH<2R=4R''ERIC5MRI_N8s5CoNs88I0H8ER-48MFI04FRd=2RRRH2CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R ERIC5MRI_N8s5CoNs88I0H8ER-48MFI04FRd=2RRRH2CCD#R''j;R
RRRRRRCRSMo8RCsMCNR0Cz;.6
-S-RRQV58N8s8IH0<ER=dR42FRMRHIs0CCRMDNLCsRFR0FkbRk0CLMND#CRCODC0FRDoRHOM8CCCR8
SRRRR.SznRR:H5VRNs88I0H8E=R<R24dRMoCC0sNCR
SRRRRRRRRRsRRF_k0CHM52=R<R''4;S
SSFSIkC0_M25HRR<=';4'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RW;R
RRRRRRCRSMo8RCsMCNR0Cz;.n
-S-RMtCC0sNCER0CqR)vCRODRD#NRM80-sH#00NCR#
RRRRRSRRzR.(:FRVsRR[H5MRI0H8Ek_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0RC
RRRRRRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)RAqUv_4Xg..:7RRLDNCHDR#WR""R;
RRRRRRRRRRRRRLRRCMoH
RRRRRRRRRRRR)SAqUv_4Xg..:7RRv)qA_4n11._.R
SRRRRRRRRRbRRFRs0lRNb5q7QRR=>HsM_C.o5*4[+RI8FMR0F.2*[,7Rq7R)q=D>RFII_Ns885R4.8MFI0jFR27,RQ=AR>jR"jR",q)77A>R=RIDF_8sN84s5.FR8IFM0R,j2
SSSRRRR Rhq='>R4R',1q1)RR=>',j'RqW RR=>I_s0CHM52B,RpRiq=B>RpRi, RhA='>R4R',1A1)RR=>',j'RAW RR=>',j'RiBpA>R=RiBp,S
SSRRRRq7m5R42=I>RF_k0L.k#5.H,*4[+27,Rmjq52>R=RkIF0k_L#H.5,[.*27,Rm4A52>R=RksF0k_L#H.5,[.*+,42RA7m5Rj2=s>RF_k0L.k#5RH,.2*[2R;
RRRRRRRRRRRRRsRRF_k0s5Co.2*[RR<=s0Fk_#Lk.,5H.2*[RCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRsRRF_k0s5Co.+*[4<2R=FRskL0_k5#.H*,.[2+4RCIEMsR5F_k0CHM52RR='24'R#CDCZR''S;
SISSF_k0s5Co.2*[RR<=I0Fk_#Lk.,5H.2*[RCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRIRRF_k0s5Co.+*[4<2R=FRIkL0_k5#.H*,.[2+4RCIEMIR5F_k0CHM52RR='24'R#CDCZR''
;
RRRRRRRRS8CMRMoCC0sNC.Rz(R;
RRRRS8CMRMoCC0sNC.RzcR;
RCRRMo8RCsMCNR0Cz;.dR
R
SRRRRR--tCCMsCN0RC0ERv)qRDOCDN#RM#8RCODC0FRDoRHOVRFs)Aqv41n_cc_1
.SzURR:H5VROHEFOIC_HE80Rc=R2CRoMNCs0SC
z	OE:VRHR85N8HsI8R0E>.R42CRoMNCs0
CRRRRRRRRRk	ODRb:RsCFO#B#5p
i2RRRRRRRRRoLCHRM
RRRRRRRRRRHV5iBp'CCPMN0RMB8Rp=iRR''42ER0CRM
RRRRRRRRRsRR_8N8sC_so85N8HsI8-0E4FR8IFM0R24.RR<=)7q7)85N8HsI8-0E4FR8IFM0R24.;R
RRRRRRRRRCRM8H
V;RRRRRRRRCRM8bOsFCR##k	OD;R
SR8CMRMoCC0sNCORzE
	;RRRRSgz.RV:RFHsRRRHM5b8C0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CSR--Q5VRNs88I0H8ERR>4R.2M8CCRR0FONsC0ICRsCH0RNCMLRDCNRM8Fbk0kC0RMDNLCCR#D0CORoDFHRO
RRRRRSRRzRdj:VRHR85N8HsI8R0E>.R42CRoMNCs0SC
-V-RHVGRFOsRNRDD4UdU(#,RCODC0VRFRH0s#00NCFRM0CRLHRMosHCo#s0CCR8
RRRRRRRRRRRRRsRRF_k0CHM52=R<R''4RCIEMsR5_8N8sC_so85N8HsI8-0E4FR8IFM0R24.RH=R2DRC#'CRj
';SSSSI0Fk_5CMH<2R=4R''ERIC5MRI_N8s5CoNs88I0H8ER-48MFI04FR.-2RRRH2CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R ERIC5MRI_N8s5CoNs88I0H8ER-48MFI04FR.=2RRRH2CCD#R''j;R
RRRRRRCRSMo8RCsMCNR0Cz;dj
-S-RRQV58N8s8IH0<ER=.R42FRMRHIs0CCRMDNLCsRFR0FkbRk0CLMND#CRCODC0FRDoRHOM8CCCR8
SRRRRdSz4RR:H5VRNs88I0H8E=R<R24.RMoCC0sNCS
SSFSskC0_M25HRR<=';4'
SSSSkIF0M_C5RH2<'=R4
';RRRRRRRRRRRRRRRRI_s0CHM52=R<R;W 
RRRRRRRRMSC8CRoMNCs0zCRd
4;SR--tCCMsCN0RC0ERv)qRDOCDN#RM08Rs#H-0CN0#R
RRRRRRzRSd:.RRsVFRH[RMIR5HE80_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNCR
RRRRRRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqA)vj_cgcnX7RR:DCNLD#RHR""W;R
RRRRRRRRRRRRRRCRLo
HMRRRRRRRRRRRRSqA)vj_cgcnX7RR:)Aqv41n_cc_1
RSRRRRRRRRRRFRbsl0RN5bR7RQq=H>RMC_so*5c[R+d8MFI0cFR*,[2R7q7)=qR>FRDIN_I858s484RF0IMF2Rj,QR7A>R=Rj"jj,j"R7q7)=AR>FRDIN_s858s484RF0IMF2Rj,S
SShS q>R=R''4,1R1)=qR>jR''W,R =qR>sRI0M_C5,H2RiBpq>R=RiBp,hR A>R=R''4,1R1)=AR>jR''W,R =AR>jR''B,RpRiA=B>Rp
i,SSSS75mqd=2R>FRIkL0_k5#cHc,R*d[+2
,RSSSS75mq.=2R>FRIkL0_k5#cH*,c[2+.,SR
S7SSm4q52>R=RkIF0k_L#Hc5,[c*+,42RS
SSmS7q25jRR=>I0Fk_#Lkc,5HR[c*2S,
S7SSmdA52>R=RksF0k_L#Hc5,*Rc[2+d,SR
S7SSm.A52>R=RksF0k_L#Hc5,[c*+,.2RS
SSmS7A254RR=>s0Fk_#Lkc,5Hc+*[4R2,
SSSSA7m5Rj2=s>RF_k0Lck#5RH,c2*[2S;
SsSSF_k0s5Coc2*[RR<=s0Fk_#Lkc,5Hc2*[RCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRsRRF_k0s5Coc+*[4<2R=FRskL0_k5#cH*,c[2+4RCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRsRRF_k0s5Coc+*[.<2R=FRskL0_k5#cH*,c[2+.RCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRsRRF_k0s5Coc+*[d<2R=FRskL0_k5#cH*,c[2+dRCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRIRRF_k0s5Coc2*[RR<=I0Fk_#Lkc,5Hc2*[RCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRIRRF_k0s5Coc+*[4<2R=FRIkL0_k5#cH*,c[2+4RCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRIRRF_k0s5Coc+*[.<2R=FRIkL0_k5#cH*,c[2+.RCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRIRRF_k0s5Coc+*[d<2R=FRIkL0_k5#cH*,c[2+dRCIEMIR5F_k0CHM52RR='24'R#CDCZR''
;
RRRRRRRRS8CMRMoCC0sNCdRz.R;
RRRRS8CMRMoCC0sNC.RzgR;
RCRRMo8RCsMCNR0Cz;.U
R
SR-RR-CRtMNCs00CRE)CRqOvRC#DDR8NMRD#CCRO0DHFoOFRVsqR)vnA4__1g1Sg
zRdd:VRHRE5OFCHO_8IH0=ERRRg2oCCMsCN0
OSzE:	RRRHV58N8s8IH0>ERR244RMoCC0sNCR
RRRRRRORkD:	RRFbsO#C#5iBp2R
RRRRRRLRRCMoH
RRRRRRRRHRRVBR5pCi'P0CMR8NMRiBpR'=R4R'20MEC
RRRRRRRRRRRRNs_8_8ss5CoNs88I0H8ER-48MFI04FR4<2R=qR)757)Ns88I0H8ER-48MFI04FR4
2;RRRRRRRRRMRC8VRH;R
RRRRRRMRC8sRbF#OC#ORkD
	;SCRRMo8RCsMCNR0Cz	OE;R
RRzRSd:cRRsVFRHHRM8R5CEb0_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNC-
S-VRQR85N8HsI8R0E>4R42CRMC08RFsROCCN0RHIs0CCRMDNLCMRN8kRF00bkRNCMLRDC#CCDOD0RFOoH
RRRRRRRRdSz6RR:H5VRNs88I0H8ERR>4R42oCCMsCN0
-S-RGVHRsVFRDONDdR4U,U(RD#CCRO0F0VRs0H#NR0CMRF0LMCHoCRso0H#C8sC
RRRRRRRRRRRRRRRRksF0M_C5RH2<'=R4I'RERCM5Ns_8_8ss5CoNs88I0H8ER-48MFI04FR4=2RRRH2CCD#R''j;S
SSFSIkC0_M25HRR<='R4'IMECRN5I8C_so85N8HsI8-0E4FR8IFM0R244RH=R2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0CHM52=R<RRW IMECRN5I8C_so85N8HsI8-0E4FR8IFM0R244RH=R2DRC#'CRj
';RRRRRRRRS8CMRMoCC0sNCdRz6S;
-Q-RVNR58I8sHE80RR<=4R42MIFRsCH0RNCMLRDCFFsRkk0b0MRCNCLDRD#CCRO0DHFoOCRMC88C
RRSRSRRzRdn:VRHR85N8HsI8R0E<4=R4o2RCsMCN
0CSRRRRRRRRRRRRksF0M_C5RH2<'=R4
';SSSSI0Fk_5CMH<2R=4R''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=W
 ;RRRRRRRRS8CMRMoCC0sNCdRznS;
-t-RCsMCNR0C0REC)RqvODCD#MRN8sR0H0-#N#0C
RRRRRRRRdSz(RR:VRFs[MRHRH5I8_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
RRRRRRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVAv)q_c.jU7XURD:RNDLCRRH#";W"
RRRRRRRRRRRRRRRRoLCHRM
RRRRRRRRRSRRAv)q_c.jU7XUR):Rq4vAng_1_
1gRRRRRRRRRRRRRRRRRFRbsl0RN5bR7RQq=H>RMC_so*5g[R+(8MFI0gFR*,[2R7q7)=qR>FRDIN_I858s48jRF0IMF2Rj,QR7A>R=Rj"jjjjjj,j"R7q7)=AR>FRDIN_s858s48jRF0IMF2Rj,S
SShS q>R=R''4,1R1)=qR>jR''W,R =qR>sRI0M_C5,H2RiBpq>R=RiBp,hR A>R=R''4,1R1)=AR>jR''W,R =AR>jR''B,RpRiA=B>RpRi,
SSSSq7m5R(2=I>RF_k0LUk#5UH,*([+2
,RSSSS75mqn=2R>FRIkL0_k5#UH*,U[2+n,SR
S7SSm6q52>R=RkIF0k_L#HU5,[U*+,62RS
SSmS7q25cRR=>I0Fk_#LkU,5HU+*[cR2,
SSSSq7m5Rd2=I>RF_k0LUk#5UH,*d[+2
,RSSSS75mq.=2R>FRIkL0_k5#UH*,U[2+.,SR
S7SSm4q52>R=RkIF0k_L#HU5,[U*+,42RS
SSmS7q25jRR=>I0Fk_#LkU,5HU2*[,SR
S7SSm(A52>R=RksF0k_L#HU5,[U*+,(2RS
SSmS7A25nRR=>s0Fk_#LkU,5HU+*[nR2,
SSSSA7m5R62=s>RF_k0LUk#5UH,*6[+2
,RSSSS75mAc=2R>FRskL0_k5#UH*,U[2+c,SR
S7SSmdA52>R=RksF0k_L#HU5,[U*+,d2RS
SSmS7A25.RR=>s0Fk_#LkU,5HU+*[.R2,
SSSSA7m5R42=s>RF_k0LUk#5UH,*4[+2
,RSSSS75mAj=2R>FRskL0_k5#UH*,U[R2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRu7Qq25jRR=>HsM_Cgo5*U[+27,RQRuA=">Rj
",RRRRRRRRRRRRRRRRRRRRRRRRRRRR7qmu5Rj2=I>RbHNs0L$_k5#UH2,[,mR7ujA52>R=RNsbs$H0_#LkU,5H[;22
RRRRRRRRRRRRRRRRksF0C_so*5g[<2R=FRskL0_k5#UH*,U[I2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRksF0C_so*5g[2+4RR<=s0Fk_#LkU,5HU+*[4I2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRksF0C_so*5g[2+.RR<=s0Fk_#LkU,5HU+*[.I2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRksF0C_so*5g[2+dRR<=s0Fk_#LkU,5HU+*[dI2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRksF0C_so*5g[2+cRR<=s0Fk_#LkU,5HU+*[cI2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRksF0C_so*5g[2+6RR<=s0Fk_#LkU,5HU+*[6I2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRksF0C_so*5g[2+nRR<=s0Fk_#LkU,5HU+*[nI2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRksF0C_so*5g[2+(RR<=s0Fk_#LkU,5HU+*[(I2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRksF0C_so*5g[2+URR<=ssbNH_0$LUk#5[H,2ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRI0Fk_osC5[g*2=R<RkIF0k_L#HU5,[U*2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRI0Fk_osC5[g*+R42<I=RF_k0LUk#5UH,*4[+2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRI0Fk_osC5[g*+R.2<I=RF_k0LUk#5UH,*.[+2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRI0Fk_osC5[g*+Rd2<I=RF_k0LUk#5UH,*d[+2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRI0Fk_osC5[g*+Rc2<I=RF_k0LUk#5UH,*c[+2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRI0Fk_osC5[g*+R62<I=RF_k0LUk#5UH,*6[+2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRI0Fk_osC5[g*+Rn2<I=RF_k0LUk#5UH,*n[+2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRI0Fk_osC5[g*+R(2<I=RF_k0LUk#5UH,*([+2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRI0Fk_osC5[g*+RU2<I=RbHNs0L$_k5#UH2,[RCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRSRRCRM8oCCMsCN0R(zd;R
RRSRRCRM8oCCMsCN0Rczd;R
RRMRC8CRoMNCs0zCRd
d;
RSRR-R-RMtCC0sNCER0CqR)vCRODRD#NRM8#CCDOD0RFOoHRsVFRv)qA_4n1_4U1
4USUzdRH:RVOR5EOFHCH_I8R0E=UR42CRoMNCs0SC
z	OERH:RVNR58I8sHE80R4>Rjo2RCsMCN
0CRRRRRRRRk	ODRb:RsCFO#B#5p
i2RRRRRRRRRoLCHRM
RRRRRRRRRRHV5iBp'CCPMN0RMB8Rp=iRR''42ER0CRM
RRRRRRRRRsRR_8N8sC_so85N8HsI8-0E4FR8IFM0R24jRR<=)7q7)85N8HsI8-0E4FR8IFM0R24j;R
RRRRRRRRRCRM8H
V;RRRRRRRRCRM8bOsFCR##k	OD;R
SRMRC8CRoMNCs0zCRO;E	
RRRRdSzgRR:VRFsHMRHRC58b_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
-S-RRQV58N8s8IH0>ERR24jRCMC8FR0RCOsNR0CI0sHCMRCNCLDR8NMR0FkbRk0CLMND#CRCODC0FRDo
HORRRRRRRRSjzcRH:RVNR58I8sHE80R4>Rjo2RCsMCN
0CSR--VRHGVRFsODNDRU4dUR(,#CCDOF0RVsR0HN#00MCRFL0RCoHMRosCHC#0s
C8RRRRRRRRRRRRRRRRs0Fk_5CMH<2R=4R''ERIC5MRs8_N8ss_CNo58I8sHE80-84RF0IMFjR42RR=HC2RDR#C';j'
SSSSkIF0M_C5RH2<'=R4I'RERCM58IN_osC58N8s8IH04E-RI8FMR0F4Rj2=RRH2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0CHM52=R<RRW IMECRN5I8C_so85N8HsI8-0E4FR8IFM0R24jRH=R2DRC#'CRj
';RRRRRRRRS8CMRMoCC0sNCcRzjS;
-Q-RVNR58I8sHE80RR<=4Rj2MIFRsCH0RNCMLRDCFFsRkk0b0MRCNCLDRD#CCRO0DHFoOCRMC88C
RRSRSRRzRc4:VRHR85N8HsI8R0E<4=Rjo2RCsMCN
0CSRRRRRRRRRRRRksF0M_C5RH2<'=R4
';SSSSI0Fk_5CMH<2R=4R''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=W
 ;RRRRRRRRS8CMRMoCC0sNCcRz4S;
-t-RCsMCNR0C0REC)RqvODCD#MRN8sR0H0-#N#0C
RRRRRRRRcSz.RR:VRFs[MRHRH5I8_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
RRRRRRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVAv)q_.4jcnX47RR:DCNLD#RHR""W;R
RRRRRRRRRRRRRRCRLo
HMRRRRRRRRRRRRSqA)vj_4.4cXn:7RRv)qA_4n1_4U1
4URRRRRRRRRRRRRRRRRFRbsl0RN5bR7RQq=H>RMC_soU54*4[+6FR8IFM0R*4U[R2,q)77q>R=RIDF_8IN8gs5RI8FMR0FjR2,7RQA=">Rjjjjjjjjjjjjjjjj"q,R7A7)RR=>D_FIs8N8sR5g8MFI0jFR2S,
S SSh=qR>4R''1,R1R)q='>RjR',WR q=I>RsC0_M25H,pRBi=qR>pRBi ,Rh=AR>4R''1,R1R)A='>RjR',WR A='>RjR',BApiRR=>B,piRS
SSmS7q6542>R=RkIF0k_L#54nHn,4*4[+6R2,
SSSSq7m524cRR=>I0Fk_#Lk4Hn5,*4n[c+42
,RSSSS75mq4Rd2=I>RF_k0L4k#n,5H4[n*+24d,SR
S7SSm4q5.=2R>FRIkL0_kn#454H,n+*[4,.2RS
SSmS7q4542>R=RkIF0k_L#54nHn,4*4[+4R2,
SSSSq7m524jRR=>I0Fk_#Lk4Hn5,*4n[j+42
,RSSSS75mqg=2R>FRIkL0_kn#454H,n+*[gR2,
SSSSq7m5RU2=I>RF_k0L4k#n,5H4[n*+,U2RS
SSmS7q25(RR=>I0Fk_#Lk4Hn5,*4n[2+(,SR
S7SSmnq52>R=RkIF0k_L#54nHn,4*n[+2
,RSSSS75mq6=2R>FRIkL0_kn#454H,n+*[6R2,
SSSSq7m5Rc2=I>RF_k0L4k#n,5H4[n*+,c2RS
SSmS7q25dRR=>I0Fk_#Lk4Hn5,*4n[2+d,SR
S7SSm.q52>R=RkIF0k_L#54nHn,4*.[+2
,RSSSS75mq4=2R>FRIkL0_kn#454H,n+*[4R2,
SSSSq7m5Rj2=I>RF_k0L4k#n,5H4[n*2
,RSSSS75mA4R62=s>RF_k0L4k#n,5H4[n*+246,SR
S7SSm4A5c=2R>FRskL0_kn#454H,n+*[4,c2RS
SSmS7Ad542>R=RksF0k_L#54nHn,4*4[+dR2,
SSSSA7m524.RR=>s0Fk_#Lk4Hn5,*4n[.+42
,RSSSS75mA4R42=s>RF_k0L4k#n,5H4[n*+244,SR
S7SSm4A5j=2R>FRskL0_kn#454H,n+*[4,j2RS
SSmS7A25gRR=>s0Fk_#Lk4Hn5,*4n[2+g,SR
S7SSmUA52>R=RksF0k_L#54nHn,4*U[+2
,RSSSS75mA(=2R>FRskL0_kn#454H,n+*[(R2,
SSSSA7m5Rn2=s>RF_k0L4k#n,5H4[n*+,n2RS
SSmS7A256RR=>s0Fk_#Lk4Hn5,*4n[2+6,SR
S7SSmcA52>R=RksF0k_L#54nHn,4*c[+2
,RSSSS75mAd=2R>FRskL0_kn#454H,n+*[dR2,
SSSSA7m5R.2=s>RF_k0L4k#n,5H4[n*+,.2RS
SSmS7A254RR=>s0Fk_#Lk4Hn5,*4n[2+4,SR
S7SSmjA52>R=RksF0k_L#54nHn,4*,[2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRQR7u=qR>MRH_osC5*4U[(+4RI8FMR0F4[U*+24n,QR7u=AR>jR"j
",RRRRRRRRRRRRRRRRRRRRRRRRRRRR7qmu5R42=I>RbHNs0L$_kn#45.H,*4[+27,Rm5uqj=2R>bRIN0sH$k_L#54nH*,.[
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRR7Amu5R42=s>RbHNs0L$_kn#45.H,*4[+27,Rm5uAj=2R>bRsN0sH$k_L#54nH*,.[;22
RRRRRRRRRRRRRRRRksF0C_soU54*R[2<s=RF_k0L4k#n,5H4[n*2ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRs0Fk_osC5*4U[2+4RR<=s0Fk_#Lk4Hn5,*4n[2+4RCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRsRRF_k0s5Co4[U*+R.2<s=RF_k0L4k#n,5H4[n*+R.2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRsks0_C4o5U+*[d<2R=FRskL0_kn#454H,n+*[dI2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRksF0C_soU54*c[+2=R<RksF0k_L#54nHn,4*c[+2ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRs0Fk_osC5*4U[2+6RR<=s0Fk_#Lk4Hn5,*4n[2+6RCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRsRRF_k0s5Co4[U*+Rn2<s=RF_k0L4k#n,5H4[n*+Rn2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRsks0_C4o5U+*[(<2R=FRskL0_kn#454H,n+*[(I2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRksF0C_soU54*U[+2=R<RksF0k_L#54nHn,4*U[+2ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRs0Fk_osC5*4U[2+gRR<=s0Fk_#Lk4Hn5,*4n[2+gRCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRsRRF_k0s5Co4[U*+24jRR<=s0Fk_#Lk4Hn5,*4n[j+42ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRs0Fk_osC5*4U[4+42=R<RksF0k_L#54nHn,4*4[+4I2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRksF0C_soU54*4[+.<2R=FRskL0_kn#454H,n+*[4R.2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRsks0_C4o5U+*[4Rd2<s=RF_k0L4k#n,5H4[n*+24dRCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRsRRF_k0s5Co4[U*+24cRR<=s0Fk_#Lk4Hn5,*4n[c+42ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRs0Fk_osC5*4U[6+42=R<RksF0k_L#54nHn,4*4[+6I2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRksF0C_soU54*4[+n<2R=bRsN0sH$k_L#54nH*,.[I2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRksF0C_soU54*4[+(<2R=bRsN0sH$k_L#54nH*,.[2+4RCIEMsR5F_k0CHM52RR='24'R#CDCZR''
;
RRRRRRRRRRRRRRRRI0Fk_osC5*4U[<2R=FRIkL0_kn#454H,n2*[RCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRIRRF_k0s5Co4[U*+R42<I=RF_k0L4k#n,5H4[n*+R42IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRIks0_C4o5U+*[.<2R=FRIkL0_kn#454H,n+*[.I2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRkIF0C_soU54*d[+2=R<RkIF0k_L#54nHn,4*d[+2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRI0Fk_osC5*4U[2+cRR<=I0Fk_#Lk4Hn5,*4n[2+cRCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRIRRF_k0s5Co4[U*+R62<I=RF_k0L4k#n,5H4[n*+R62IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRIks0_C4o5U+*[n<2R=FRIkL0_kn#454H,n+*[nI2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRkIF0C_soU54*([+2=R<RkIF0k_L#54nHn,4*([+2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRI0Fk_osC5*4U[2+URR<=I0Fk_#Lk4Hn5,*4n[2+URCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRIRRF_k0s5Co4[U*+Rg2<I=RF_k0L4k#n,5H4[n*+Rg2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRIks0_C4o5U+*[4Rj2<I=RF_k0L4k#n,5H4[n*+24jRCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRIRRF_k0s5Co4[U*+244RR<=I0Fk_#Lk4Hn5,*4n[4+42ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRI0Fk_osC5*4U[.+42=R<RkIF0k_L#54nHn,4*4[+.I2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRkIF0C_soU54*4[+d<2R=FRIkL0_kn#454H,n+*[4Rd2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRIks0_C4o5U+*[4Rc2<I=RF_k0L4k#n,5H4[n*+24cRCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRIRRF_k0s5Co4[U*+246RR<=I0Fk_#Lk4Hn5,*4n[6+42ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRI0Fk_osC5*4U[n+42=R<RNIbs$H0_#Lk4Hn5,[.*2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRI0Fk_osC5*4U[(+42=R<RNIbs$H0_#Lk4Hn5,[.*+R42IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R

RRRRRSRRCRM8oCCMsCN0R.zc;R
RRSRRCRM8oCCMsCN0Rgzd;R
RRMRC8CRoMNCs0zCRd
U;
RSRR-R-RMtCC0sNCER0CqR)vCRODRD#NRM8#CCDOD0RFOoHRsVFRv)qA_4n1_dn1
dnSUzdNRR:H5VROHEFOIC_HE80Rd=Rno2RCsMCN
0CSEzO	RR:H5VRNs88I0H8ERR>go2RCsMCN
0CSRRRRDkO	RR:bOsFC5##B2pi
RSSLHCoMS
SRVRHRp5BiP'CCRM0NRM8BRpi=4R''02RE
CMSRSRR_RsNs88_osC58N8s8IH04E-RI8FMR0Fg<2R=qR)757)Ns88I0H8ER-48MFI0gFR2S;
SCRRMH8RVS;
S8CMRFbsO#C#RDkO	S;
RCRRMo8RCsMCNR0Cz	OE;R
SRzRRdRgN:FRVsRRHH5MR80CbEk_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0SC
-Q-RVNR58I8sHE80Rg>R2CRMC08RFsROCCN0RHIs0CCRMDNLCMRN8kRF00bkRNCMLRDC#CCDOD0RFOoH
SSSzNcjRH:RVNR58I8sHE80Rg>R2CRoMNCs0SC
-V-RHVGRFOsRNRDD4UdU(#,RCODC0VRFRH0s#00NCFRM0CRLHRMosHCo#s0CCS8
SsSSF_k0CHM52=R<R''4RCIEMsR5_8N8sC_so85N8HsI8-0E4FR8IFM0RRg2=2RHR#CDCjR''S;
SISSF_k0CHM52=R<R''4RCIEMIR5Ns8_CNo58I8sHE80-84RF0IMF2RgRH=RRC2RDR#C';j'
SSSS0Is_5CMH<2R= RWRCIEMIR5Ns8_CNo58I8sHE80-84RF0IMF2RgRH=R2DRC#'CRj
';SCSSMo8RCsMCNR0CzNcj;-
S-VRQR85N8HsI8R0E<g=R2FRMRHIs0CCRMDNLCsRFR0FkbRk0CLMND#CRCODC0FRDoRHOM8CCCS8
ScSz4:NRRRHV58N8s8IH0<ER=2RgRMoCC0sNCS
SSFSskC0_M25HRR<=';4'
SSSSkIF0M_C5RH2<'=R4
';SSSSI_s0CHM52=R<R;W 
SSSCRM8oCCMsCN0R4zcNS;
-t-RCsMCNR0C0REC)RqvODCD#MRN8sR0H0-#N#0C
SSSzNc.RV:RF[sRRRHM58IH0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CRRRRRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FAVR)_qv6X4.dR.7:NRDLRCDH"#RW
";RRRRRRRRRRRRRRRRLHCoMS
SS)SAq6v_4d.X.:7RRv)qA_4n1_dn1
dnRRRRRRRRRRRRRRRRRRRRb0FsRblNRQ57q>R=R_HMs5Cod[n*+Rd48MFI0dFRn2*[,7Rq7R)q=D>RFII_Ns8858URF0IMF2Rj,QR7A>R=Rj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjj,j"R7q7)=AR>FRDIN_s858sUFR8IFM0R,j2
SSSSq hRR=>',4'R)11q>R=R''j, RWq>R=R0Is_5CMHR2,BqpiRR=>B,piRA hRR=>',4'R)11A>R=R''j, RWA>R=R''j,pRBi=AR>pRBiS,
S7SSmdq54=2R>FRIkL0_k.#d5dH,.+*[d,42RS
SSmS7qj5d2>R=RkIF0k_L#5d.H.,d*d[+j
2,SSSS75mq.Rg2=I>RF_k0Ldk#.,5Hd[.*+2.g,SR
S7SSm.q5U=2R>FRIkL0_k.#d5dH,.+*[.,U2RS
SSmS7q(5.2>R=RkIF0k_L#5d.H.,d*.[+(
2,SSSS75mq.Rn2=I>RF_k0Ldk#.,5Hd[.*+2.n,SR
S7SSm.q56=2R>FRIkL0_k.#d5dH,.+*[.,62RS
SSmS7qc5.2>R=RkIF0k_L#5d.H.,d*.[+c
2,SSSS75mq.Rd2=I>RF_k0Ldk#.,5Hd[.*+2.d,SR
S7SSm.q5.=2R>FRIkL0_k.#d5dH,.+*[.,.2RS
SSmS7q45.2>R=RkIF0k_L#5d.H.,d*.[+4
2,SSSS75mq.Rj2=I>RF_k0Ldk#.,5Hd[.*+2.j,SR
S7SSm4q5g=2R>FRIkL0_k.#d5dH,.+*[4,g2RS
SSmS7qU542>R=RkIF0k_L#5d.H.,d*4[+U
2,SSSS75mq4R(2=I>RF_k0Ldk#.,5Hd[.*+24(,SR
S7SSm4q5n=2R>FRIkL0_k.#d5dH,.+*[4,n2RS
SSmS7q6542>R=RkIF0k_L#5d.H.,d*4[+6
2,SSSS75mq4Rc2=I>RF_k0Ldk#.,5Hd[.*+24c,SR
S7SSm4q5d=2R>FRIkL0_k.#d5dH,.+*[4,d2RS
SSmS7q.542>R=RkIF0k_L#5d.H.,d*4[+.
2,SSSS75mq4R42=I>RF_k0Ldk#.,5Hd[.*+244,SR
S7SSm4q5j=2R>FRIkL0_k.#d5dH,.+*[4,j2RS
SSmS7q25gRR=>I0Fk_#LkdH.5,*d.[2+g,S
SSmS7q25URR=>I0Fk_#LkdH.5,*d.[2+U,SR
S7SSm(q52>R=RkIF0k_L#5d.H.,d*([+2
,RSSSS75mqn=2R>FRIkL0_k.#d5dH,.+*[n
2,SSSS75mq6=2R>FRIkL0_k.#d5dH,.+*[6R2,
SSSSq7m5Rc2=I>RF_k0Ldk#.,5Hd[.*+,c2RS
SSmS7q25dRR=>I0Fk_#LkdH.5,*d.[2+d,S
SSmS7q25.RR=>I0Fk_#LkdH.5,*d.[2+.,SR
S7SSm4q52>R=RkIF0k_L#5d.H.,d*4[+2
,RSSSS75mqj=2R>FRIkL0_k.#d5dH,.2*[,S
SSmS7A45d2>R=RksF0k_L#5d.H.,d*d[+4R2,
SSSSA7m52djRR=>s0Fk_#LkdH.5,*d.[j+d2S,
S7SSm.A5g=2R>FRskL0_k.#d5dH,.+*[.,g2RS
SSmS7AU5.2>R=RksF0k_L#5d.H.,d*.[+UR2,
SSSSA7m52.(RR=>s0Fk_#LkdH.5,*d.[(+.2S,
S7SSm.A5n=2R>FRskL0_k.#d5dH,.+*[.,n2RS
SSmS7A65.2>R=RksF0k_L#5d.H.,d*.[+6R2,
SSSSA7m52.cRR=>s0Fk_#LkdH.5,*d.[c+.2S,
S7SSm.A5d=2R>FRskL0_k.#d5dH,.+*[.,d2RS
SSmS7A.5.2>R=RksF0k_L#5d.H.,d*.[+.R2,
SSSSA7m52.4RR=>s0Fk_#LkdH.5,*d.[4+.2S,
S7SSm.A5j=2R>FRskL0_k.#d5dH,.+*[.,j2RS
SSmS7Ag542>R=RksF0k_L#5d.H.,d*4[+gR2,
SSSSA7m524URR=>s0Fk_#LkdH.5,*d.[U+42S,
S7SSm4A5(=2R>FRskL0_k.#d5dH,.+*[4,(2RS
SSmS7An542>R=RksF0k_L#5d.H.,d*4[+nR2,
SSSSA7m5246RR=>s0Fk_#LkdH.5,*d.[6+42S,
S7SSm4A5c=2R>FRskL0_k.#d5dH,.+*[4,c2RS
SSmS7Ad542>R=RksF0k_L#5d.H.,d*4[+dR2,
SSSSA7m524.RR=>s0Fk_#LkdH.5,*d.[.+42S,
S7SSm4A54=2R>FRskL0_k.#d5dH,.+*[4,42RS
SSmS7Aj542>R=RksF0k_L#5d.H.,d*4[+jR2,
SSSSA7m5Rg2=s>RF_k0Ldk#.,5Hd[.*+,g2
SSSSA7m5RU2=s>RF_k0Ldk#.,5Hd[.*+,U2RS
SSmS7A25(RR=>s0Fk_#LkdH.5,*d.[2+(,SR
S7SSmnA52>R=RksF0k_L#5d.H.,d*n[+2S,
S7SSm6A52>R=RksF0k_L#5d.H.,d*6[+2
,RSSSS75mAc=2R>FRskL0_k.#d5dH,.+*[cR2,
SSSSA7m5Rd2=s>RF_k0Ldk#.,5Hd[.*+,d2
SSSSA7m5R.2=s>RF_k0Ldk#.,5Hd[.*+,.2RS
SSmS7A254RR=>s0Fk_#LkdH.5,*d.[2+4,SR
S7SSmjA52>R=RksF0k_L#5d.H.,d*,[2
RRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRQRuq=H>RMC_son5d*d[+6FR8IFM0R*dn[.+d27,RQRuA=">Rjjjj"R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRu7mq25dRR=>IsbNH_0$Ldk#.,5Hc+*[dR2,7qmu5R.2=I>RbHNs0L$_k.#d5cH,*.[+2R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRu7mq254RR=>IsbNH_0$Ldk#.,5Hc+*[4R2,7qmu5Rj2=I>RbHNs0L$_k.#d5cH,*,[2
RRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRm5uAd=2R>bRsN0sH$k_L#5d.H*,c[2+d,mR7u.A52>R=RNsbs$H0_#LkdH.5,[c*+,.2
RRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRm5uA4=2R>bRsN0sH$k_L#5d.H*,c[2+4,mR7ujA52>R=RNsbs$H0_#LkdH.5,[c*2
2;RRRRRRRRRRRRRRRRRFRsks0_Cdo5n2*[RR<=s0Fk_#LkdH.5,*d.[I2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRsRRF_k0s5Cod[n*+R42<s=RF_k0Ldk#.,5Hd[.*+R42IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRs0Fk_osC5*dn[2+.RR<=s0Fk_#LkdH.5,*d.[2+.RCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRksF0C_son5d*d[+2=R<RksF0k_L#5d.H.,d*d[+2ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRsks0_Cdo5n+*[c<2R=FRskL0_k.#d5dH,.+*[cI2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRsRRF_k0s5Cod[n*+R62<s=RF_k0Ldk#.,5Hd[.*+R62IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRs0Fk_osC5*dn[2+nRR<=s0Fk_#LkdH.5,*d.[2+nRCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRksF0C_son5d*([+2=R<RksF0k_L#5d.H.,d*([+2ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRsks0_Cdo5n+*[U<2R=FRskL0_k.#d5dH,.+*[UI2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRsRRF_k0s5Cod[n*+Rg2<s=RF_k0Ldk#.,5Hd[.*+Rg2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRs0Fk_osC5*dn[j+42=R<RksF0k_L#5d.H.,d*4[+jI2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRsRRF_k0s5Cod[n*+244RR<=s0Fk_#LkdH.5,*d.[4+42ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRsks0_Cdo5n+*[4R.2<s=RF_k0Ldk#.,5Hd[.*+24.RCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRksF0C_son5d*4[+d<2R=FRskL0_k.#d5dH,.+*[4Rd2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRs0Fk_osC5*dn[c+42=R<RksF0k_L#5d.H.,d*4[+cI2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRsRRF_k0s5Cod[n*+246RR<=s0Fk_#LkdH.5,*d.[6+42ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRsks0_Cdo5n+*[4Rn2<s=RF_k0Ldk#.,5Hd[.*+24nRCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRksF0C_son5d*4[+(<2R=FRskL0_k.#d5dH,.+*[4R(2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRs0Fk_osC5*dn[U+42=R<RksF0k_L#5d.H.,d*4[+UI2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRsRRF_k0s5Cod[n*+24gRR<=s0Fk_#LkdH.5,*d.[g+42ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRsks0_Cdo5n+*[.Rj2<s=RF_k0Ldk#.,5Hd[.*+2.jRCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRksF0C_son5d*.[+4<2R=FRskL0_k.#d5dH,.+*[.R42IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRs0Fk_osC5*dn[.+.2=R<RksF0k_L#5d.H.,d*.[+.I2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRsRRF_k0s5Cod[n*+2.dRR<=s0Fk_#LkdH.5,*d.[d+.2ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRsks0_Cdo5n+*[.Rc2<s=RF_k0Ldk#.,5Hd[.*+2.cRCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRksF0C_son5d*.[+6<2R=FRskL0_k.#d5dH,.+*[.R62IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRs0Fk_osC5*dn[n+.2=R<RksF0k_L#5d.H.,d*.[+nI2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRsRRF_k0s5Cod[n*+2.(RR<=s0Fk_#LkdH.5,*d.[(+.2ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRsks0_Cdo5n+*[.RU2<s=RF_k0Ldk#.,5Hd[.*+2.URCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRksF0C_son5d*.[+g<2R=FRskL0_k.#d5dH,.+*[.Rg2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRs0Fk_osC5*dn[j+d2=R<RksF0k_L#5d.H.,d*d[+jI2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRsRRF_k0s5Cod[n*+2d4RR<=s0Fk_#LkdH.5,*d.[4+d2ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRsks0_Cdo5n+*[dR.2<s=RbHNs0L$_k.#d5cH,*R[2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRs0Fk_osC5*dn[d+d2=R<RNsbs$H0_#LkdH.5,[c*+R42IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRs0Fk_osC5*dn[c+d2=R<RNsbs$H0_#LkdH.5,[c*+R.2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRs0Fk_osC5*dn[6+d2=R<RNsbs$H0_#LkdH.5,[c*+Rd2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRR
RRRRRRRRRRRRRRRRIRRF_k0s5Cod[n*2=R<RkIF0k_L#5d.H.,d*R[2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRI0Fk_osC5*dn[2+4RR<=I0Fk_#LkdH.5,*d.[2+4RCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRkIF0C_son5d*.[+2=R<RkIF0k_L#5d.H.,d*.[+2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRIks0_Cdo5n+*[d<2R=FRIkL0_k.#d5dH,.+*[dI2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRIRRF_k0s5Cod[n*+Rc2<I=RF_k0Ldk#.,5Hd[.*+Rc2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRI0Fk_osC5*dn[2+6RR<=I0Fk_#LkdH.5,*d.[2+6RCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRkIF0C_son5d*n[+2=R<RkIF0k_L#5d.H.,d*n[+2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRIks0_Cdo5n+*[(<2R=FRIkL0_k.#d5dH,.+*[(I2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRIRRF_k0s5Cod[n*+RU2<I=RF_k0Ldk#.,5Hd[.*+RU2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRI0Fk_osC5*dn[2+gRR<=I0Fk_#LkdH.5,*d.[2+gRCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRkIF0C_son5d*4[+j<2R=FRIkL0_k.#d5dH,.+*[4Rj2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRI0Fk_osC5*dn[4+42=R<RkIF0k_L#5d.H.,d*4[+4I2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRIRRF_k0s5Cod[n*+24.RR<=I0Fk_#LkdH.5,*d.[.+42ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRIks0_Cdo5n+*[4Rd2<I=RF_k0Ldk#.,5Hd[.*+24dRCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRkIF0C_son5d*4[+c<2R=FRIkL0_k.#d5dH,.+*[4Rc2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRI0Fk_osC5*dn[6+42=R<RkIF0k_L#5d.H.,d*4[+6I2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRIRRF_k0s5Cod[n*+24nRR<=I0Fk_#LkdH.5,*d.[n+42ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRIks0_Cdo5n+*[4R(2<I=RF_k0Ldk#.,5Hd[.*+24(RCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRkIF0C_son5d*4[+U<2R=FRIkL0_k.#d5dH,.+*[4RU2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRI0Fk_osC5*dn[g+42=R<RkIF0k_L#5d.H.,d*4[+gI2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRIRRF_k0s5Cod[n*+2.jRR<=I0Fk_#LkdH.5,*d.[j+.2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRIks0_Cdo5n+*[.R42<I=RF_k0Ldk#.,5Hd[.*+2.4RCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRkIF0C_son5d*.[+.<2R=FRIkL0_k.#d5dH,.+*[.R.2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRI0Fk_osC5*dn[d+.2=R<RkIF0k_L#5d.H.,d*.[+dI2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRIRRF_k0s5Cod[n*+2.cRR<=I0Fk_#LkdH.5,*d.[c+.2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRIks0_Cdo5n+*[.R62<I=RF_k0Ldk#.,5Hd[.*+2.6RCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRkIF0C_son5d*.[+n<2R=FRIkL0_k.#d5dH,.+*[.Rn2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRI0Fk_osC5*dn[(+.2=R<RkIF0k_L#5d.H.,d*.[+(I2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRIRRF_k0s5Cod[n*+2.URR<=I0Fk_#LkdH.5,*d.[U+.2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRIks0_Cdo5n+*[.Rg2<I=RF_k0Ldk#.,5Hd[.*+2.gRCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRkIF0C_son5d*d[+j<2R=FRIkL0_k.#d5dH,.+*[dRj2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRI0Fk_osC5*dn[4+d2=R<RkIF0k_L#5d.H.,d*d[+4I2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRIRRF_k0s5Cod[n*+2d.RR<=IsbNH_0$Ldk#.,5Hc2*[RCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRkIF0C_son5d*d[+d<2R=bRIN0sH$k_L#5d.H*,c[2+4RCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRkIF0C_son5d*d[+c<2R=bRIN0sH$k_L#5d.H*,c[2+.RCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRkIF0C_son5d*d[+6<2R=bRIN0sH$k_L#5d.H*,c[2+dRCIEMIR5F_k0CHM52RR='24'R#CDCZR''
;
SCSSMo8RCsMCNR0CzNc.;S
SCRM8oCCMsCN0RgzdNS;
CRM8oCCMsCN0RUzdNR;
R8CMRMoCC0sNCcRzd
;
RcRzcRR:H5VRMRF0s8N8sC_soo2RCsMCNR0C-o-RCsMCNR0C#CCDOs0RNRl
R-RR-VRQR8N8s8IH0<ERRN6R#o#HMjR''FR0RkkM#RC8L#H0
RRRRRzjRH:RVNR58I8sHE80R4=R2CRoMNCs0RC
RRRRRDRRFsI_Ns88_<#R=jR"jjjj"RR&s_N8s_Co#25j;R
RRRRRRFRDIN_I8_8s#=R<Rj"jj"jjRI&RNs8_C#o_5;j2
RRRR8CMRMoCC0sNCjRz;R
RR4RzRRR:H5VRNs88I0H8ERR=.o2RCsMCN
0CRRRRRRRRD_FIs8N8sR_#<"=Rjjjj"RR&s_N8s_Co#R548MFI0jFR2R;
RRRRRDRRFII_Ns88_<#R=jR"j"jjRI&RNs8_C#o_584RF0IMF2Rj;R
RRMRC8CRoMNCs0zCR4R;
RzRR.:RRRRHV58N8s8IH0=ERRRd2oCCMsCN0
RRRRRRRRIDF_8sN8#s_RR<="jjj"RR&s_N8s_Co#R5.8MFI0jFR2R;
RRRRRDRRFII_Ns88_<#R=jR"jRj"&NRI8C_so5_#.FR8IFM0R;j2
RRRR8CMRMoCC0sNC.Rz;R
RRdRzRRR:H5VRNs88I0H8ERR=co2RCsMCN
0CRRRRRRRRD_FIs8N8sR_#<"=RjRj"&NRs8C_so5_#dFR8IFM0R;j2
RRRRRRRRIDF_8IN8#s_RR<=""jjRI&RNs8_C#o_58dRF0IMF2Rj;R
RRMRC8CRoMNCs0zCRdS;
z:cSRRHV58N8s8IH0=ERRR62oCCMsCN0
DSSFsI_Ns88_<#R=jR''RR&s_N8s_Co#R5c8MFI0jFR2S;
SIDF_8IN8#s_RR<='Rj'&NRI8C_so5_#cFR8IFM0R;j2
MSC8CRoMNCs0zCRcR;
RzRR6:RRRRHV58N8s8IH0>ERRR62oCCMsCN0
RRRRRRRRIDF_8sN8#s_RR<=s_N8s_Co#R568MFI0jFR2R;
RRRRRDRRFII_Ns88_<#R=NRI8C_so5_#6FR8IFM0R;j2
RRRR8CMRMoCC0sNC6Rz;R

R-RR-VRQRH58MC_sos2RC#oH0RCs7RQhkM#HopRBiR
RRnRzRRR:H5VR8_HMs2CoRMoCC0sNCR
RRRRRRsRbF#OC#BR5pRi,72QhRoLCHRM
RRRRRRRRRHRRVBR5p=iRR''4R8NMRiBp'CCPMR020MEC
RRRRRRRRRRRRRRRR_HMs_Co#=R<Rh7Q;R
RRRRRRRRRRMRC8VRH;R
RRRRRRMRC8sRbF#OC#R;
RCRRMo8RCsMCNR0Cz
n;RRRRzR(R:VRHRF5M0HR8MC_soo2RCsMCN
0CRRRRRRRRRRRRHsM_C#o_RR<=7;Qh
RRRR8CMRMoCC0sNC(Rz;R

R-RR-VRQR85sF_k0s2CoRosCHC#0smR7zkaR#oHMRpmBiR
RRURzs:RRRRHV5Fs8ks0_CRo2oCCMsCN0
RRRRRRRRFbsO#C#R_5)miBp,FRsks0_C#o_2CRLo
HMRRRRRRRRRRRRH5VR)B_mp=iRR''4R8NMRm)_B'piCMPC002RE
CMRRRRRRRRRRRRRRRR)m_7z<aR=FRsks0_C#o_;R
RRRRRRRRRRMRC8VRH;R
RRRRRRMRC8sRbF#OC#R;
RCRRMo8RCsMCNR0Cz;Us
RRRRszgRRR:H5VRMRF0sk8F0C_soo2RCsMCN
0CRRRRRRRRRRRR)m_7z<aR=FRsks0_C#o_;R
RRMRC8CRoMNCs0zCRg
s;
USzI:RRRRHV5FI8ks0_CRo2oCCMsCN0
RRRRRRRRFbsO#C#R_5WmiBp,FRIks0_C#o_2CRLo
HMRRRRRRRRRRRRH5VRWB_mp=iRR''4R8NMRmW_B'piCMPC002RE
CMRRRRRRRRRRRRRRRRWm_7z<aR=FRIks0_C#o_;R
RRRRRRRRRRMRC8VRH;R
RRRRRRMRC8sRbF#OC#R;
RCRRMo8RCsMCNR0Cz;UI
RRRRIzgRRR:H5VRMRF0Ik8F0C_soo2RCsMCN
0CRRRRRRRRRRRRWm_7z<aR=FRIks0_C#o_;R
RRMRC8CRoMNCs0zCRg
I;
RRRRR--Q5VRs8N8sC_sos2RC#oH0RCsq)77RHk#MBoRpRi
RzRR4RjR:VRHRN5s8_8ss2CoRMoCC0sNCR
RRRRRRsRbF#OC#)R5_pmBi),Rq)772CRLo
HMRRRRRRRRRRRRH5VR)B_mp=iRR''4R8NMRm)_B'piCMPC002RE
CMRRRRRRRRRRRRRRRRs_N8s_Co#=R<R7)q7N)58I8sHE80-84RF0IMF2Rj;R
RRRRRRRRRRMRC8VRH;R
RRRRRRMRC8sRbF#OC#R;
RCRRMo8RCsMCNR0Cz;4j
RRRR4z4RH:RVMR5Fs0RNs88_osC2CRoMNCs0RC
RRRRRRRRRsRRNs8_C#o_RR<=)7q7)R;
RCRRMo8RCsMCNR0Cz;44
R
RR-R-RRQV58IN8ss_CRo2sHCo#s0CR7q7)#RkHRMoB
piRRRRzR4.RH:RVIR5Ns88_osC2CRoMNCs0RC
RRRRRbRRsCFO#5#RB,piR7Wq7R)2LHCoMR
RRRRRRRRRRVRHRp5BiRR='R4'NRM8B'piCMPC002RE
CMRRRRRRRRRRRRRRRRI_N8s_Co#=R<R7Wq7N)58I8sHE80-84RF0IMF2Rj;R
RRRRRRRRRRMRC8VRH;R
RRRRRRMRC8sRbF#OC#R;
RCRRMo8RCsMCNR0Cz;4.
RRRRdz4RH:RVMR5FI0RNs88_osC2CRoMNCs0RC
RRRRRRRRRIRRNs8_C#o_RR<=W7q7)R;
RCRRMo8RCsMCNR0Cz;4d
RRRRRRRRR
RR-R-RMtCC0sNCER0CqR)vCRODRD#NRM8#CCDOD0RFOoH
RRRRcz4RV:RFHsRRRHM5lMk_DOCDc_nR4-R2FR8IFM0RojRCsMCN
0CRRRR-Q-RVNR58I8sHE80R6>R2CRMC08RFsROCCN0RHIs0CCRMDNLCMRN8kRF00bkRNCMLRDC#CCDOD0RFOoH
RRRRRRRR6z4RH:RVNR58I8sHE80Rn>R2CRoMNCs0RC
RRRRRRRRRRRRRsRRF_k0C#M_5RH2<'=R4I'RERCM58sN_osC_N#58I8sHE80-84RF0IMF2RnRH=R2DRC#'CRj
';SSSSI0Fk__CM#25HRR<='R4'IMECRN5I8C_so5_#Ns88I0H8ER-48MFI0nFR2RR=HC2RDR#C';j'
RRRRRRRRRRRRRRRR0Is__CM#25HRR<=WI RERCM58IN_osC_N#58I8sHE80-84RF0IMF2RnRH=R2DRC#'CRj
';RRRRRRRRCRM8oCCMsCN0R6z4;R
RR-R-RRQV58N8s8IH0<ER=2R6RRMFI0sHCMRCNCLDRRFsFbk0kC0RMDNLCCR#D0CORoDFHMORCCC88R
RRRRRR4RznRR:H5VRNs88I0H8E=R<RRn2oCCMsCN0
RRRRRRRRRRRRRRRRksF0M_C_H#52=R<R''4;S
SSFSIkC0_M5_#H<2R=4R''R;
RRRRRRRRRRRRRIRRsC0_M5_#H<2R= RW;R
RRRRRRMRC8CRoMNCs0zCR4
n;RRRR-t-RCsMCNR0C0REC)RqvODCD#MRN8sR0H0-#N#0C
RRRRRRRR(z4RV:RF[sRRRHM58IH0-ERRR428MFI0jFRRMoCC0sNCR
RRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqz)vRnc:NRDLRCDH"#R1"7aRH&RMo0CCHs'lCNo58IH0RE2&7R""RR&HCM0o'CsHolNC*5HnRc2&WR""RR&HCM0o'CsHolNC25[R"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05+5H4n2*c8,RCEb02&2RR""XRH&RMo0CCHs'lCNo54[+2R;
RRRRRRRRRLRRCMoH
RRRRRRRRRRRRqz)vRnc:)RXqcvnXR47
RRRRRRRRRRRRRRRRsbF0NRlb7R5RR=>HsM_C#o_5,[2RRqj=D>RFII_Ns88_j#52q,R4>R=RIDF_8IN8#s_5,42RRq.=D>RFII_Ns88_.#52R,
RRRRRRRRRRRRRRRRRRRRRRRRRRqd=D>RFII_Ns88_d#52q,Rc>R=RIDF_8IN8#s_5,c2RRq6=D>RFII_Ns88_6#52
,RSSSSSRSR7qu)j>R=RIDF_8sN8#s_5,j2R)7uq=4R>FRDIN_s8_8s#254,uR7)Rq.=D>RFsI_Ns88_.#52S,
SSSSS7RRud)qRR=>D_FIs8N8s5_#dR2,7qu)c>R=RIDF_8sN8#s_5,c2R)7uq=6R>FRDIN_s8_8s#256,SR
SSSSSWRR >R=R0Is__CM#25H,BRWp=iR>pRBi7,Ru=mR>FRskL0_kn#_cH#5,,[2Rm1uRR=>I0Fk_#Lk_#nc5[H,2
2;RRRRRRRRRRRRRRRRs0Fk_osC_[#52=R<RksF0k_L#c_n#,5H[I2RERCM5ksF0M_C_H#52RR='24'R#CDCZR''S;
SISSF_k0s_Co#25[RR<=I0Fk_#Lk_#nc5[H,2ERIC5MRI0Fk__CM#25HR'=R4R'2CCD#R''Z;R
RRRRRRMRC8CRoMNCs0zCR4
(;RRRRR8CMRMoCC0sNC4RzcR;RRRRRRRRRRRR
RRRRRR
RR-R-RMtCC0sNCRRNdI.RFRs88bCCRv)qRDOCDVRHRbNbssFbHCN0RRRRRRRRRRRRR
RRRRRRzR4U:VRHRk5MlC_ODdD_.RR=4o2RCsMCN
0CRRRR-Q-RVNR58I8sHE80R(>R2CRMC08RFsROCCN0RHIs0CCRMDNLCMRN8kRF00bkRNCMLRDC#CCDOD0RFOoH
RRRRRRRRgz4NRR:H5VRNs88I0H8ERR>no2RCsMCN
0CRRRRRRRRRRRRRRRRs0Fk__CMd<.R=4R''ERIC5MR58sN_osC_N#58I8sHE80-84RF0IMF2RnRM=RkOl_C_DDnRc2NRM858sN_osC_6#52RR='2j'2DRC#'CRj
';SSSSI0Fk__CMd<.R=4R''ERIC5MR58IN_osC_N#58I8sHE80-84RF0IMF2RnRM=RkOl_C_DDnRc2NRM858IN_osC_6#52RR='2j'2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0CdM_.=R<RRW IMECRI55Ns8_C#o_58N8s8IH04E-RI8FMR0Fn=2RRlMk_DOCDc_n2MRN8IR5Ns8_C#o_5R62=jR''R22CCD#R''j;R
RRRRRRMRC8CRoMNCs0zCR4;gN
RRRRRRRRgz4LRR:H5VRNs88I0H8ERR=nMRN8kRMlC_ODnD_cRR=jo2RCsMCN
0CRRRRRRRRRRRRRRRRs0Fk__CMd<.R=4R''ERIC5MR58sN_osC_6#52RR='2j'2DRC#'CRj
';SSSSI0Fk__CMd<.R=4R''ERIC5MR58IN_osC_6#52RR='2j'2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0CdM_.=R<RRW IMECRI55Ns8_C#o_5R62=jR''R22CCD#R''j;R
RRRRRRMRC8CRoMNCs0zCR4;gLRRRR-Q-RVNR58I8sHE80RR<=6M2RFsRIHR0CCLMNDFCRskRF00bkRNCMLRDC#CCDOD0RFOoHRCMC8
C8RRRRRRRRzR.j:VRHR85N8HsI8R0E<6=R2CRoMNCs0RC
RRRRRRRRRRRRRsRRF_k0CdM_.=R<R''4;S
SSFSIkC0_M._dRR<=';4'
RRRRRRRRRRRRRRRR0Is__CMd<.R= RW;R
RRRRRRMRC8CRoMNCs0zCR.
j;RRRR-t-RCsMCNR0C0REC)RqvODCDR8NMRH0s-N#00RC
RRRRRzRR.:4RRsVFRH[RMIR5HE80R4-R2FR8IFM0RojRCsMCN
0CRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FzVR)dqv.RR:DCNLD#RHR7"1a&"RR0HMCsoC'NHloIC5HE802RR&"R7"&MRH0CCosl'HN5oCM_klODCD_*ncnRc2&WR""RR&HCM0o'CsHolNC25[R"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05lMk_DOCDc_n*Rnc+.Rd,CR8b20E2RR&"RX"&MRH0CCosl'HN5oC[2+4;R
RRRRRRRRRRCRLo
HMRRRRRRRRRRRRzv)qd:.RRqX)vXd.4
7RRRRRRRRRRRRRRRRRb0FsRblNRR57=H>RMC_so5_#[R2,q=jR>FRDIN_I8_8s#25j,4RqRR=>D_FII8N8s5_#4R2,q=.R>FRDIN_I8_8s#25.,R
RRRRRRRRRRRRRRRRRRRRRRRRRq=dR>FRDIN_I8_8s#25d,cRqRR=>D_FII8N8s5_#cR2,
SSSSRSSR)7uq=jR>FRDIN_s8_8s#25j,uR7)Rq4=D>RFsI_Ns88_4#527,Ru.)qRR=>D_FIs8N8s5_#.
2,SSSSSRSR7qu)d>R=RIDF_8sN8#s_5,d2R)7uq=cR>FRDIN_s8_8s#25c,SR
SSSSSWRR >R=R0Is__CMdR.,WiBpRR=>B,piRm7uRR=>s0Fk_#Lk_#d.5lMk_DOCD._d,,[2Rm1uRR=>I0Fk_#Lk_#d.5lMk_DOCD._d,2[2;R
RRRRRRRRRRRRRRFRsks0_C#o_5R[2<s=RF_k0L_k#d5.#M_klODCD_,d.[I2RERCM5ksF0M_C_Rd.=4R''C2RDR#C';Z'
SSSSkIF0C_so5_#[<2R=FRIkL0_kd#_.M#5kOl_C_DDd[.,2ERIC5MRI0Fk__CMd=.RR''42DRC#'CRZ
';RRRRRRRRR8CMRMoCC0sNC.Rz4R;
RRRRCRM8oCCMsCN0RUz4;RRRRRRRR
RR
RRRRR--tCCMsCN0R4NRnFRIs88RCRCb)RqvODCDRRHVNsbbFHbsNR0CRRRRRRRRRRRRRRR
RzRR.:.RRRHV5lMk_DOCDn_4R4=R2CRoMNCs0RC
R-RR-VRQR85N8HsI8R0E>2R6RCMC8FR0RCOsNR0CI0sHCMRCNCLDR8NMR0FkbRk0CLMND#CRCODC0FRDo
HORRRRRRRRzN.dRH:RVNR58I8sHE80Rn>RR8NMRlMk_DOCD._dR4=R2CRoMNCs0RC
RRRRRRRRRRRRRsRRF_k0C4M_n=R<R''4RCIEM5R5s_N8s_Co#85N8HsI8-0E4FR8IFM0RRn2=kRMlC_ODnD_cN2RM58Rs_N8s_Co#256R'=R4R'2NRM858sN_osC_c#52RR='2j'2DRC#'CRj
';SSSSI0Fk__CM4<nR=4R''ERIC5MR58IN_osC_N#58I8sHE80-84RF0IMF2RnRM=RkOl_C_DDnRc2NRM858IN_osC_6#52RR='24'R8NMRN5I8C_so5_#c=2RR''j2C2RDR#C';j'
RRRRRRRRRRRRRRRR0Is__CM4<nR= RWRCIEM5R5I_N8s_Co#85N8HsI8-0E4FR8IFM0RRn2=kRMlC_ODnD_cN2RM58RI_N8s_Co#256R'=R4R'2NRM858IN_osC_c#52RR='2j'2DRC#'CRj
';RRRRRRRRCRM8oCCMsCN0Rdz.NR;
RRRRRzRR.RdL:VRHR85N8HsI8R0E>RRnNRM8M_klODCD_Rd./4=R2CRoMNCs0RC
RRRRRRRRRRRRRsRRF_k0C4M_n=R<R''4RCIEM5R5s_N8s_Co#85N8HsI8-0E4FR8IFM0RRn2=kRMlC_ODnD_cN2RM58Rs_N8s_Co#256R'=RjR'2NRM858sN_osC_c#52RR='2j'2DRC#'CRj
';SSSSI0Fk__CM4<nR=4R''ERIC5MR58IN_osC_N#58I8sHE80-84RF0IMF2RnRM=RkOl_C_DDnRc2NRM858IN_osC_6#52RR='2j'R8NMRN5I8C_so5_#c=2RR''j2C2RDR#C';j'
RRRRRRRRRRRRRRRR0Is__CM4<nR= RWRCIEM5R5I_N8s_Co#85N8HsI8-0E4FR8IFM0RRn2=kRMlC_ODnD_cN2RM58RI_N8s_Co#256R'=RjR'2NRM858IN_osC_c#52RR='2j'2DRC#'CRj
';RRRRRRRRCRM8oCCMsCN0Rdz.LR;
RRRRRzRR.RdO:VRHR85N8HsI8R0E=RRnNRM8M_klODCD_Rd.=2R4RMoCC0sNCR
RRRRRRRRRRRRRRFRskC0_Mn_4RR<='R4'IMECRs55Ns8_C#o_5R62=4R''N2RM58Rs_N8s_Co#25cR'=Rj2'2R#CDCjR''S;
SISSF_k0C4M_n=R<R''4RCIEM5R5I_N8s_Co#256R'=R4R'2NRM858IN_osC_c#52RR='2j'2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0C4M_n=R<RRW IMECRI55Ns8_C#o_5R62=4R''N2RM58RI_N8s_Co#25cR'=Rj2'2R#CDCjR''R;
RRRRRCRRMo8RCsMCNR0CzO.d;R
RRRRRR.Rzd:8RRRHV58N8s8IH0=ERRN6RMM8RkOl_C_DDd/.R=2R4RMoCC0sNCR
RRRRRRRRRRRRRRFRskC0_Mn_4RR<='R4'IMECRs55Ns8_C#o_58N8s8IH04E-RI8FMR0Fc=2RRlMk_DOCD._d2C2RDR#C';j'
SSSSkIF0M_C_R4n<'=R4I'RERCM5N5I8C_so5_#Ns88I0H8ER-48MFI0cFR2RR=M_klODCD_2d.2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0C4M_n=R<RRW IMECRI55Ns8_C#o_58N8s8IH04E-RI8FMR0Fc=2RRlMk_DOCD._d2C2RDR#C';j'
RRRRRRRR8CMRMoCC0sNC.RzdR8;R-RR-VRQR85N8HsI8R0E<6=R2FRMRHIs0CCRMDNLCsRFR0FkbRk0CLMND#CRCODC0FRDoRHOM8CCCR8
RRRRRzRR.:cRRRHV58N8s8IH0<ER=2RcRMoCC0sNCR
RRRRRRRRRRRRRRFRskC0_Mn_4RR<=';4'
SSSSkIF0M_C_R4n<'=R4
';RRRRRRRRRRRRRRRRI_s0C4M_n=R<R;W 
RRRRRRRR8CMRMoCC0sNC.RzcR;
R-RR-CRtMNCs00CRE)CRqOvRCRDDNRM80-sH#00NCR
RRRRRR.Rz6RR:VRFs[MRHRH5I8R0E-2R4RI8FMR0FjCRoMNCs0RC
RRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)Rzqnv4RD:RNDLCRRH#"a17"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloMC5kOl_C_DDnnc*cRR+M_klODCD_*d.dR.2&WR""RR&HCM0o'CsHolNC25[R"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05lMk_DOCDc_n*Rnc+kRMlC_ODdD_..*dR4+Rn8,RCEb02&2RR""XRH&RMo0CCHs'lCNo54[+2R;
RRRRRRRRRLRRCMoH
RRRRRRRRRRRRqz)vR4n:qR)vX4n4
7RRRRRRRRRRRRRRRRRb0FsRblNRR57=H>RMC_so5_#[R2,q=jR>FRDIN_I8_8s#25j,4RqRR=>D_FII8N8s5_#4R2,q=.R>FRDIN_I8_8s#25.,R
RRRRRRRRRRRRRRRRRRRRRRRRRq=dR>FRDIN_I8_8s#25d,uR7)Rqj=D>RFsI_Ns88_j#527,Ru4)qRR=>D_FIs8N8s5_#4R2,7qu).>R=RIDF_8sN8#s_5,.2
SSSSRSSR)7uq=dR>FRDIN_s8_8s#25d, RWRR=>I_s0C4M_nW,RBRpi=B>RpRi,7Rum=s>RF_k0L_k#45n#M_klODCD_,4n[R2,1Rum=I>RF_k0L_k#45n#M_klODCD_,4n[;22
RRRRRRRRRRRRRRRRksF0C_so5_#[<2R=FRskL0_k4#_nM#5kOl_C_DD4[n,2ERIC5MRs0Fk__CM4=nRR''42DRC#'CRZ
';SSSSI0Fk_osC_[#52=R<RkIF0k_L#n_4#k5MlC_OD4D_n2,[RCIEMIR5F_k0C4M_nRR='24'R#CDCZR''R;
RRRRRCRRMo8RCsMCNR0Cz;.6
RRRR8CMRMoCC0sNC.Rz.R;RRRR
R8CMRMoCC0sNCcRzcC;
MN8RsHOE00COkRsCMsF_IE_OC;O	
-
-
-----
--p-RNR#0HDlbCMlC0HN0FHMR#CR8VDNk0-
--#-RCODC0N_sls
NO0EHCkO0s#CRCODC0N_slVRFRv)q_u)W_H)R#k
VMHO0FoMRCC0_M88_CEb05x#HCRR:HCM0oRCs;CR8bR0E:MRH0CCoss2RCs0kMMRH0CCos#RH
sPNHDNLCHRlMH_#x:CRR0HMCsoCRR:=jL;
CMoH
lRRH#M_HRxC:8=RCEb0;R
RH5VR#CHxR8<RCEb02ER0CRM
RlRRH#M_HRxC:#=RH;xC
CRRMH8RVR;
R0sCkRsMl_HM#CHx;M
C8CRo0M_C8C_8b;0E
MOF#M0N0kRMlC_ODRD#:MRH0CCos=R:R855CEb0R4-R2n/42R;RRRRRRRRRR-R-RFyRVqR)vX4n4O7RC#DDRCMC8
C80C$bR0Fk_#Lk_b0$C#RHRsNsN5$RM_klODCD#FR8IFM0RRj,I0H8ER-48MFI0jFR2VRFR8#0_oDFH
O;#MHoNsDRF_k0LRk#:kRF0k_L#$_0bRC;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFVsF_8k50RHkMb0FR0RH0s-N#002C#
o#HMRNDs0Fk_RCM:0R#8F_Do_HOP0COFMs5kOl_C#DDRI8FMR0FjR2;RRRRR-R-RNCML#DCRsVFRH0s-N#00
C##MHoNIDRF_k0C:MRR8#0_oDFHPO_CFO0sk5MlC_ODRD#8MFI0jFR2#;
HNoMDFRIkL0_k:#RR0Fk_#Lk_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$FIVR_k8F0HR5M0bkRR0F0-sH#00NC
#2#MHoNIDRsC0_MRR:#_08DHFoOC_POs0F5lMk_DOCD8#RF0IMF2Rj;RRRRRRRRR--I0sHCMRCNCLD#FRVsNRCOsERFFIRVqR)vCROD
D##MHoNHDRMC_soRR:#_08DHFoOC_POs0F58IH04E-RI8FMR0FjR2;RRRRRRRRRR--k8#CRR0FsHCo#s0CRh7QRH
#oDMNRksF0C_soRR:#_08DHFoOC_POs0F58IH04E-RI8FMR0FjR2;RRRRR-RR-#RkC08RFCRso0H#C)sR_z7maH
#oDMNRkIF0C_soRR:#_08DHFoOC_POs0F58IH04E-RI8FMR0FjR2;RRRRR-RR-#RkC08RFCRso0H#CWsR_z7maH
#oDMNR8sN_osCR#:R0D8_FOoH_OPC05FsNs88I0H8ER-48MFI0jFR2R;RR-RR-#RkC08RFCRso0H#C)sRq)77
o#HMRNDI_N8sRCo:0R#8F_Do_HOP0COFNs58I8sHE80-84RF0IMF2Rj;RRRR-R-RCk#8FR0RosCHC#0sqRW7
7)#MHoNDDRFsI_Ns88R#:R0D8_FOoH_OPC05FsdFR8IFM0R;j2RRRRRRRRRRRRRR--s8N8sHRL0H#RM0bkRR0F)RqvODCD#cR5R0LH#CRsJskHC
82#MHoNDDRFII_Ns88R#:R0D8_FOoH_OPC05FsdFR8IFM0R;j2RRRRRRRRRRRRRR--I8N8sHRL0H#RM0bkRR0F)RqvODCD#cR5R0LH#CRsJskHC
82Ns00H0LkC3R\s_NlF#VVCR0\:0R#soHM;L

CMoH
R
RR-R-RRQVNs88I0H8ERR<c#RN#MHoR''jRR0Fk#MkCL8RH
0#RRRRzR4R:VRHR85N8HsI8R0E=2R4RMoCC0sNCR
RRRRRRFRDIN_s8R8s<"=Rj"jjRs&RNs8_Cjo52R;
RRRRRDRRFII_Ns88RR<="jjj"RR&I_N8s5Coj
2;RRRRCRM8oCCMsCN0R;z4
RRRRRz.RH:RVNR58I8sHE80R.=R2CRoMNCs0RC
RRRRRDRRFsI_Ns88RR<=""jjRs&RNs8_C4o5RI8FMR0Fj
2;RRRRRRRRD_FII8N8s=R<Rj"j"RR&I_N8s5Co4FR8IFM0R;j2
RRRR8CMRMoCC0sNC.Rz;R
RRdRzRRR:H5VRNs88I0H8ERR=do2RCsMCN
0CRRRRRRRRD_FIs8N8s=R<R''jRs&RNs8_C.o5RI8FMR0Fj
2;RRRRRRRRD_FII8N8s=R<R''jRI&RNs8_C.o5RI8FMR0Fj
2;RRRRCRM8oCCMsCN0R;zd
RRRRRzcRH:RVNR58I8sHE80Rd>R2CRoMNCs0RC
RRRRRDRRFsI_Ns88RR<=s_N8s5CodFR8IFM0R;j2
RRRRRRRRIDF_8IN8<sR=NRI8C_soR5d8MFI0jFR2R;
RCRRMo8RCsMCNR0Cz
c;
RRRRR--Q5VR8_HMs2CoRosCHC#0sQR7h#RkHRMoB
piRRRRzR6R:VRHRH58MC_soo2RCsMCN
0CRRRRRRRRbOsFCR##5iBp,QR7hL2RCMoH
RRRRRRRRRRRRRHV5iBpR'=R4N'RMB8RpCi'P0CM2ER0CRM
RRRRRRRRRRRRRHRRMC_so=R<Rh7Q;R
RRRRRRRRRRMRC8VRH;R
RRRRRRMRC8sRbF#OC#R;
RCRRMo8RCsMCNR0Cz
6;RRRRzRnR:VRHRF5M0HR8MC_soo2RCsMCN
0CRRRRRRRRRRRRHsM_C<oR=QR7hR;
RCRRMo8RCsMCNR0Cz
n;
RRRRR--Q5VRs0Fk_osC2CRso0H#C7sRmRzakM#HoBRmpRi
RzRR(RsR:VRHR85sF_k0s2CoRMoCC0sNCR
RRRRRRsRbF#OC#)R5_pmBis,RF_k0s2CoRoLCHRM
RRRRRRRRRHRRV)R5_pmBiRR='R4'NRM8)B_mpCi'P0CM2ER0CRM
RRRRRRRRRRRRR)RR_z7ma=R<RksF0C_soR;
RRRRRRRRRCRRMH8RVR;
RRRRRCRRMb8RsCFO#
#;RRRRCRM8oCCMsCN0Rsz(;R
RRURzs:RRRRHV50MFRFs8ks0_CRo2oCCMsCN0
RRRRRRRRRRRR7)_mRza<s=RF_k0s;Co
RRRR8CMRMoCC0sNCURzs
;
RRRR-Q-RVsR5F_k0s2CoRosCHC#0smR7zkaR#oHMRpmBiR
RR(RzI:RRRRHV5FI8ks0_CRo2oCCMsCN0
RRRRRRRRFbsO#C#R_5WmiBp,FRIks0_CRo2LHCoMR
RRRRRRRRRRVRHR_5WmiBpR'=R4N'RMW8R_pmBiP'CC2M0RC0EMR
RRRRRRRRRRRRRR_RW7amzRR<=I0Fk_osC;R
RRRRRRRRRRMRC8VRH;R
RRRRRRMRC8sRbF#OC#R;
RCRRMo8RCsMCNR0Cz;(I
RRRRIzURRR:H5VRMRF0Ik8F0C_soo2RCsMCN
0CRRRRRRRRRRRRWm_7z<aR=FRIks0_C
o;RRRRCRM8oCCMsCN0RIzU;R

R-RR-VRQRN5s8_8ss2CoRosCHC#0sqR)7R7)kM#HoBRmpRi
RzRRg:RRRRHV58sN8ss_CRo2oCCMsCN0
RRRRRRRRFbsO#C#R_5)miBp,qR)727)RoLCHRM
RRRRRRRRRHRRV)R5_pmBiRR='R4'NRM8)B_mpCi'P0CM2ER0CRM
RRRRRRRRRRRRRsRRNs8_C<oR=qR)757)Ns88I0H8ER-48MFI0jFR2R;
RRRRRRRRRCRRMH8RVR;
RRRRRCRRMb8RsCFO#
#;RRRRCRM8oCCMsCN0R;zg
RRRRjz4RH:RVMR5Fs0RNs88_osC2CRoMNCs0RC
RRRRRRRRRsRRNs8_C<oR=qR)7;7)
RRRR8CMRMoCC0sNC4RzjR;
RRRRR
RRRRRR-Q-RVIR5Ns88_osC2CRso0H#CWsRq)77RHk#MBoRpRi
RzRR4R6R:VRHRN5I8_8ss2CoRMoCC0sNCR
RRRRRRsRbF#OC#BR5pRi,W7q7)L2RCMoH
RRRRRRRRRRRRRHV5iBpR'=R4N'RMB8RpCi'P0CM2ER0CRM
RRRRRRRRRRRRRIRRNs8_C<oR=qRW757)Ns88I0H8ER-48MFI0jFR2R;
RRRRRRRRRCRRMH8RVR;
RRRRRCRRMb8RsCFO#
#;RRRRCRM8oCCMsCN0R6z4;R
RR4RznRR:H5VRMRF0I8N8sC_soo2RCsMCN
0CRRRRRRRRRRRRI_N8sRCo<W=Rq)77;R
RRMRC8CRoMNCs0zCR4
n;
RRRRR--tCCMsCN0RC0ERv)qRDOCDN#RM#8RCODC0FRDo
HORRRRzR44:FRVsRRHHMMRkOl_C#DDRI8FMR0FjCRoMNCs0RC
RRRRR-RR-VRQR85N8HsI8R0E>2RcRCMC8FR0RCOsNR0CI0sHCMRCNCLDR8NMR0FkbRk0CLMND#CRCODC0FRDo
HORRRRRRRRzR4.:VRHR85N8HsI8R0E>2RcRMoCC0sNCR
RRRRRRRRRRRRRRFRskC0_M25HRR<='R4'IMECRN5s8C_so85N8HsI8-0E4FR8IFM0RRc2=2RHR#CDCjR''R;
RRRRRRRRRRRRRIRRF_k0CHM52=R<R''4RCIEMIR5Ns8_CNo58I8sHE80-84RF0IMF2RcRH=R2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0CHM52=R<RRW IMECRN5I8C_so85N8HsI8-0E4FR8IFM0RRc2=2RHR#CDCjR''R;
RRRRRCRRMo8RCsMCNR0Cz;4.
RRRRRRRRR--Q5VRNs88I0H8E=R<RRc2MIFRsCH0RNCMLRDCFFsRkk0b0MRCNCLDRD#CCRO0DHFoOCRMC88C
RRRRRRRRdz4RH:RVNR58I8sHE80RR<=co2RCsMCN
0CRRRRRRRRRRRRRRRRs0Fk_5CMH<2R=4R''R;
RRRRRRRRRRRRRIRRF_k0CHM52=R<R''4;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R R;
RRRRRRRRRCRRMo8RCsMCNR0Cz;4d
RRRRR--tsMCNR0C0REC)RqvODCD#MRN8sR0H0-#N#0C
RRRRRRRRcz4RV:RF[sRRRHM58IH0-ERRR428MFI0jFRRMoCC0sNCR
RRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqz)vRR:DCNLD#RHR7"1a&"RR0HMCsoC'NHloIC5HE802RR&"R7"&MRH0CCosl'HN5oCHn*42RR&"RW"&MRH0CCosl'HN5oC[&2RR"" RH&RMo0CCHs'lCNo50oC_8CM_b8C05E5H2+4*,4nRb8C02E2R"&RX&"RR0HMCsoC'NHlo[C5+;42
RRRRRRRRRRRRoLCHRM
RRRRRRRRRzRR):qvRv)q44nX7RR
RRRRRRRRRRRRRbRRFRs0lRNb5=7R>MRH_osC5,[2RRqj=D>RFII_Ns885,j2RRq4=D>RFII_Ns885,42RRq.=D>RFII_Ns885,.2
RRRRRRRRRRRRRRRRRRRRRRRRqRRd>R=RIDF_8IN8ds527,Ruj)qRR=>D_FIs8N8s25j,uR7)Rq4=D>RFsI_Ns885,42RR
RRRRRRRRRRRRRRRRRRRRRRRRR7qu).>R=RIDF_8sN8.s527,Rud)qRR=>D_FIs8N8s25d, RWRR=>I_s0CHM52
,RRRRRRRRRRRRRRRRRRRRRRRRRRBRWp=iR>pRBi7,Ru=mR>FRskL0_kH#5,,[2Rm1uRR=>I0Fk_#Lk5[H,2
2;RRRRRRRRRRRRs0Fk_osC5R[2<s=RF_k0L5k#H2,[RCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRIRRF_k0s5Co[<2R=FRIkL0_kH#5,R[2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRMRC8CRoMNCs0zCR4
c;RRRRRRRRCRM8oCCMsCN0R4z4;R
RRRRRRRRRRRRRRRRRRRRRRRRRR
RRCRM8NEsOHO0C0CksRD#CC_O0s;Nl




