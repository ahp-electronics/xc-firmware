--
@ER--B$FbsEHo0OR52gR4g-cRRj.jd$R1MHbDO$H0ROQM
R--fN]C8:CsR#//$DMbH0OH$N/lb0DN.Uj4J4.b/blNb#Cs/DGHH/MGD/HLoCCMs/HOo_CMoCCMs.HO/lsNM__sIE3P8Ry4f-
-
-
-

---1-RHDlbCqR)vHRI0#ERHDMoC7Rq71) 1FRVsFRL0sERCRN8NRM8I0sHC-
-RsaNoRC0:HRXDGHM

---4-Rj4/jR01CRQW)av _m_7 qIR5sCH0RsbF002RF R)qw7_Qa)1RRHM8NCVkRD0V
Fs-R-RRMOFVODH0CRs#kFD0MHFRsbkbCF#3CR)VRCs0eFRHCs0GQ-QRtwuqNR]MF8LF-	
-RRRBbEN0.CsR#"zHRMoAODF	CR1D0CO)RqvvFClsR$"#0COH3FM
H
DLssN$CRHC
C;kR#CHCCC38#0_oDFH4O_43ncN;DD
Ck#RCHCC03#8F_Do_HO#MHoCN83D
D;DsHLNRs$k#MHH
l;kR#Ck#MHHPl3ObFlFMMC0N#3D
D;CHM00)$Rq_vh)R_WHS#
oCCMsRHO5R
SRVRRNDlH$RR:#H0sM:oR=MR"F"MC;S
SI0H8ERR:HCM0oRCs:4=R;SR
S8N8s8IH0:ERR0HMCsoCRR:=nR;RRRRRR-R-RoLHRFCMkRoEVRFs80CbES
S80CbERR:HCM0oRCs:c=RUS;
Sk8F0C_soRR:LDFFCRNM:V=RNCD#;RRRR-RR-NRE#kRF00bkRosC
8SSHsM_C:oRRFLFDMCNRR:=V#NDCR;RRRRRR-R-R#ENR08NNMRHbRk0s
CoRRRRRRRRs_#08NN0R#:R0MsHoS;
S_IslCF8:0R#soHMRR:="QW)aw _Qa)1"S;
S8sN8ss_C:oRRFLFDMCNRR:=V#NDCR;RRRRR-E-RNs#RCRN8Ns88CR##s
CoSNSI8_8ssRCo:FRLFNDCM:RR=NRVDR#CRRRRRR--ERN#I0sHC8RN8#sC#CRsoS
S2S;
b0FsRS5
Sz7maF:Rk#0R0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2S;
S7)q7:)RRRHM#_08DHFoOC_POs0F58N8s8IH04E-RI8FMR0Fj
2;SQS7h:RRRRHM#_08DHFoOC_POs0F58IH04E-RI8FMR0Fj
2;SqSW7R7):MRHR8#0_oDFHPO_CFO0s85N8HsI8-0E4FR8IFM0R;j2
WSS :RRRRHM#_08DHFoOR;RRRRRRR--I0sHCMRCNCLDRsVFRlsN
BSSp:iRRRHM#_08DHFoOR;RRRRRRR--OODF	FRVsNRslN,R8,8sRM8H
mSSBRpi:MRHR8#0_oDFHRO;RRRRRR--FRb0OODF	FRVs_RI80Fk
RRRRRRRRR h:MRHR8#0_oDFHRO;RRRRR-RR-MRCNCLD
RRRRRRRR W_hRR:H#MR0D8_FOoH;RRRRRRRRR--CLMNDRC
RRRRR)RR1:aRRRHM#_08DHFoORRRRRRRRR--#
#sRRRRRRRR2C;
MC8RM00H$qR)v)h__
W;

---w-RH0s#RbHlDCClM00NHRFMl0k#RRLCODNDCN8RsjOE

--NEsOHO0C0CksRFLDOs	_NFlRVqR)v)h__HWR#k
VMHO0FVMRk_MOH0MH5:LRRFLFDMCN2CRs0MksRs#0HRMoHL#
CMoH
HRRVLR52ER0CRM
RsRRCs0kMh5"FCRsNI8/sCH0RMOFVODH0EROC3O	Rl1Hk0DNHRFMllH#NE0OR#bF#DHLC!R!"
2;RDRC#RC
RsRRCs0kMB5"F8kDR0MFRbHlDCClMA0RD	FORv)q3#RQRC0ERNsC88RN8#sC#CRso0H#C8sCRHk#M0oRE#CRNRlCOODF	#RNRC0ERv)q?;"2
CRRMH8RVC;
MV8Rk_MOH0MH;k
VMHO0FoMRCC0_M88_CEb05x#HCRR:HCM0oRCs;CR8bR0E:MRH0CCoss2RCs0kMMRH0CCos#RH
sPNHDNLCHRlMH_#x:CRR0HMCsoCRR:=jL;
CMoH
lRRH#M_HRxC:8=RCEb0;R
RH5VR#CHxR8<RCEb02ER0CRM
RlRRH#M_HRxC:#=RH;xC
CRRMH8RVR;
R0sCkRsMl_HM#CHx;R
RCRM8o_C0C_M880CbEN;
0H0sLCk0RMoCC0sNFss_CsbF0RR:#H0sM
o;-0-N0LsHkR0CoCCMsFN0sC_sb0FsRRFVLODF	N_slRR:NEsOHO0C0CksRRH#VOkM_HHM0N5s8_8ss2Co;-
-RoLCHLMRD	FORlsNRbHlDCClM00NHRFM#MHoN
D#VOkM0MHFRs#0H.Mo#5DPNRR:#H0sMRo2skC0s#MR0D8_FOoH_OPC0RFsHP#
NNsHLRDC#RDP:0R#8F_Do_HOP0COFNs5'oEHE'-NDRFI8MFI0jFR2P;
NNsHLRDCHRR:HCM0o;Cs
oLCHRM
RsVFRHHRMRRj0#FRDEP'HRoEDbFF
RRRRRHV5NN5'oEHE2-HR'=R4R'20MEC
RSR#5DPH:2R=4R''S;
CCD#
RSR#5DPH:2R=jR''S;
CRM8H
V;RMRC8FRDF
b;RCRs0MksRP#D;M
C80R#soHM.P#D;k
VMHO0F#MRD#P.0MsHoR5N:0R#8F_Do_HOP0COFRs2skC0s#MR0MsHo#RH
sPNHDNLCRR#:0R#soHM5EN'H-oENF'DIR+48MFI04FR2P;
NNsHLRDCHRR:HCM0o;Cs
oLCHRM
RsVFRHHRM'RNDRFI0NFR'oEHEFRDFRb
RHRRVNR55RH2=4R''02RE
CMS#RR5NH-'IDF+R42:'=R4
';S#CDCR
SRH#5-DN'F4I+2=R:R''j;C
SMH8RVR;
R8CMRFDFbR;
R0sCkRsM#C;
M#8RD#P.0MsHoN;
0H0sLCk0R_GObbsF#RR:#H0sM
o;-F-OMN#0M#0RsDPNR#:R0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2=R:Rs#0H.Mo#5DPs_#08NN02-;
-CRLoRHMLODF	NRsllRHblDCCNM00MHFRo#HM#ND
MVkOF0HMCRo0E_OFCHO_8IH0IE5HE80RH:RMo0CCRs2skC0sHMRMo0CCHsR#N
PsLHNDPCRN:DRR0HMCsoCRR:=jP;
NNsHLRDC8dHP.8,RHnP4,HR8PRU,8cHP,HR8PR.,84HPRH:RMo0CC
s;LHCoMR
R8dHP.=R:RH5I8-0E4d2/nR;
RP8H4:nR=IR5HE80-/424
U;RHR8P:UR=IR5HE80-/42gR;
RP8Hc=R:RH5I8-0E4c2/;R
R8.HPRR:=58IH04E-2;/.
8RRHRP4:5=RI0H8E2-4;R
RH5VR84HPRj>R2ER0CRM
RPRRN:DR=NRPDRR+4R;
R8CMR;HV
HRRV8R5HRP.>2RjRC0EMR
RRNRPD=R:RDPNR4+R;R
RCRM8H
V;RVRHRH58P>cRRRj20MEC
RRRRDPNRR:=PRND+;R4
CRRMH8RVR;
RRHV5P8HURR>j02RE
CMRRRRPRND:P=RN+DRR
4;RMRC8VRH;R
RH5VR84HPnRR>j02RE
CMRRRRPRND:P=RN+DRR
4;RMRC8VRH;-
-RVRHRH58PRd.>2RjRC0EM-
-RRRRPRND:P=RN+DRR
4;-R-RCRM8H
V;RVRHRN5PDRR>.02RE
CMRRRRskC0s5MR.*R*RDPNR.+RRR**5DPNRd-R2
2;RDRC#RC
RsRRCs0kM.R5RR**P2ND;R
RCRM8H
V;CRM8o_C0OHEFOIC_HE80;k
VMHO0FoMRCO0_EOFHCC_8b50E80CbERR:HCM0o2CsR0sCkRsMHCM0oRCsHP#
NNsHLRDC8E_OFCHO_b8C0:ERR0HMCsoCRR:=jL;
CMoH
HRRV8R5CEb0RU>R42g.RC0EMR
RR_R8OHEFO8C_CEb0RR:=4UndcR;
R#CDH5VR80CbE=R<RgU4.MRN8CR8bR0E>jRcg2nRRC0EMR
RR_R8OHEFO8C_CEb0RR:=U.4g;R
RCHD#V8R5CEb0RR<=cnjgR8NMRb8C0>ERRc.jU02RE
CMRRRR8E_OFCHO_b8C0:ER=jRcg
n;RDRC#RHV5b8C0<ER=jR.cNURM88RCEb0R4>RjR.c2ER0CRM
R8RR_FOEH_OC80CbE=R:Rc.jUR;
R#CDH5VR80CbE=R<R.4jcMRN8CR8bR0E>4R6.02RE
CMRRRR8E_OFCHO_b8C0:ER=jR4.
c;RDRC#RHV5b8C0<ER=4R6.02RE
CMRRRR8E_OFCHO_b8C0:ER=4R6.R;
R8CMR;HV
sRRCs0kM_R8OHEFO8C_CEb0;M
C8CRo0E_OFCHO_b8C0
E;VOkM0MHFR0oC_8IH0lE_FU8_5FOEH_OCI:8RR0HMCsoC2CRs0MksR0HMCsoCR
H#PHNsNCLDR8IH0lE_FU8_RH:RMo0CC
s;LHCoMR
RH5VROHEFOIC_8RR>U02RE
CMRRRRI0H8EF_l8R_U:O=REOFHC8_IR5-ROHEFOIC_8FRl82RU;R
RCCD#
RRRR8IH0lE_FU8_RR:=OHEFOIC_8R;
R8CMR;HV
sRRCs0kMHRI8_0El_F8UC;
Mo8RCI0_HE80_8lF_
U;
MOF#M0N0_RIOHEFOIC_HE80RH:RMo0CC:sR=CRo0E_OFCHO_8IH0IE5HE802O;
F0M#NRM0IE_OFCHO_b8C0:ERR0HMCsoCRR:=4UndcC/o0H_I8_0El_F8U_5IOHEFOIC_HE802O;
F0M#NRM08E_OFCHO_b8C0:ERR0HMCsoCRR:=o_C0OHEFO8C_CEb05b8C0;E2
MOF#M0N0_R8OHEFOIC_HE80RH:RMo0CC:sR=4R5ncdU/O8_EOFHCC_8b20ER5+R5d4nU8c/_FOEH_OC80CbE/2RR;U2
k
VMHO0FoMRCM0_kOl_C#DD5RI8:MRH0CCosE;OFCHO_RI8:MRH0CCoss2RCs0kMMRH0CCos#RH
sPNHDNLCkRMlC_ODRD#:MRH0CCosL;
CMoH
MRRkOl_C#DDRR:=5-I84O2/EOFHC8_IR4+R;R
RskC0sMMRkOl_C#DD;M
C8CRo0k_MlC_OD;D#
k
VMHO0FoMRC#0_H5xCIRMO:MRH0CCos8;RM:ORR0HMCsoC2CRs0MksR0HMCsoCR
H#LHCoMR
RR0sCkRsMIRMO*MR8OC;
Mo8RC#0_H;xC
k
VMHO0FoMRCL0_F8FD5#8_HRxC:MRH0CCosI;R_x#HCRR:HCM0o;CsRO8_IRR:HCM0o;CsROI_IRR:HCM0o2CsR0sCkRsMHCM0oRCsHL#
CMoH
RHV5#8_HRxC<I=R_x#HC02RE
CMRCRs0MksRO8_IC;
D
#CRCRs0MksROI_IC;
MH8RVC;
Mo8RCL0_F8FD;O

F0M#NRM0OHEFOIC_HE80RH:RMo0CC:sR=CRo0F_LF5D8o_C0#CHx50oC_lMk_DOCDI#5HE80,_R8OHEFOIC_HE802C,o0k_MlC_OD5D#80CbE8,R_FOEH_OC80CbE,22
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRCRo0H_#xoC5CM0_kOl_C#DD58IH0RE,IE_OFCHO_8IH0,E2o_C0M_klODCD#C58b,0EROI_EOFHCC_8b20E2S,
SSSSSSSSS8SR_FOEH_OCI0H8EI,R_FOEH_OCI0H8E
2;O#FM00NMR8IH0ME_kOl_C#DDRH:RMo0CC:sR=CRo0F_LF5D8o_C0#CHx50oC_lMk_DOCDI#5HE80,_R8OHEFOIC_HE802C,o0k_MlC_OD5D#80CbE8,R_FOEH_OC80CbE,22
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR0oC_x#HCC5o0k_MlC_OD5D#I0H8EI,R_FOEH_OCI0H8Eo2,CM0_kOl_C#DD5b8C0RE,IE_OFCHO_b8C02E2,S
SSSSSSSSSSRRRRH5I8-0E482/_FOEH_OCI0H8E5,RI0H8E2-4/OI_EOFHCH_I820ER4+R;F
OMN#0M80RCEb0_lMk_DOCD:#RR0HMCsoCRR:=o_C0LDFF8C5o0H_#xoC5CM0_kOl_C#DD58IH0RE,8E_OFCHO_8IH0,E2o_C0M_klODCD#C58b,0ERO8_EOFHCC_8b20E2R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRCRo0H_#xoC5CM0_kOl_C#DD58IH0RE,IE_OFCHO_8IH0,E2o_C0M_klODCD#C58b,0EROI_EOFHCC_8b20E2S,
SSSSSSSSSRRR5b8C04E-2_/8OHEFO8C_CEb0,8R5CEb0-/42IE_OFCHO_b8C0RE2+;R4SOR
F0M#NRM0xFCsR#:R0D8_FOoH_OPC05FsOHEFOIC_HE80*8IH0ME_kOl_C#DD-8IH04E-RI8FMR0Fj:2R=FR50sEC#>R=R''j2O;
F0M#NRM0#NsPDD_#PRR:#_08DHFoOC_POs0F5FOEH_OCI0H8EH*I8_0EM_klODCD#R-48MFI0jFR2=R:RsxCFRR&#H0sM#o.DsP5#80_N20N;F
OMN#0M#0RsDPNR#:R0MsHoE5OFCHO_8IH0IE*HE80_lMk_DOCD8#RF0IMF2R4RR:=#.DP#H0sM#o5sDPN_P#D2-;
-CRLoRHMLODF	NRsllRHblDCCNM00MHFRo#HM#ND
b0$CkRF0k_L#04_$RbCHN#Rs$sNRC58b_0EM_klODCD#R-48MFI0jFR,HRI8_0EM_klODCD#R-48MFI0jFR2VRFR8#0_oDFH
O;#MHoNFDRkL0_kR#4:kRF0k_L#04_$;bCRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$FsVR_k8F0HR5M0bkRR0F0-sH#00NC
#20C$bR0Fk_#Lk.$_0bHCR#sRNsRN$5b8C0ME_kOl_C#DD-84RF0IMF,RjRI.*HE80_lMk_DOCD4#+RI8FMR0FjF2RV0R#8F_Do;HO
o#HMRNDF_k0L.k#RF:RkL0_k_#.0C$b;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFVsF_8k50RHkMb0FR0RH0s-N#002C#
b0$CkRF0k_L#0c_$RbCHN#Rs$sNRC58b_0EM_klODCD#R-48MFI0jFR,*RcI0H8Ek_MlC_OD+D#dFR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNR0Fk_#LkcRR:F_k0Lck#_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFR8s_FRk05bHMk00RFsR0H0-#N#0C2$
0bFCRkL0_k_#U0C$bRRH#NNss$8R5CEb0_lMk_DOCD4#-RI8FMR0FjU,R*8IH0ME_kOl_C#DD+8(RF0IMF2RjRRFV#_08DHFoO#;
HNoMDkRF0k_L#:URR0Fk_#LkU$_0bRC;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RV_Rs80FkRM5HbRk000FRs#H-0CN0#02
$RbCbHNs0L$_k_#U0C$bRRH#NNss$8R5CEb0_lMk_DOCD4#-RI8FMR0FjI,RHE80_lMk_DOCD4#-RI8FMR0FjF2RV0R#8F_Do;HO
o#HMRNDbHNs0L$_kR#U:NRbs$H0_#LkU$_0bRC;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFVsF_8k50RHkMb0FR0RH0s-N#002C#
b0$CkRF0k_L#_4n0C$bRRH#NNss$8R5CEb0_lMk_DOCD4#-RI8FMR0Fj4,RnH*I8_0EM_klODCD#6+4RI8FMR0FjF2RV0R#8F_Do;HO
o#HMRNDF_k0L4k#nRR:F_k0L4k#n$_0bRC;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFVsF_8k50RHkMb0FR0RH0s-N#002C#
b0$CNRbs$H0_#Lk40n_$RbCHN#Rs$sNRC58b_0EM_klODCD#R-48MFI0jFR,*R.I0H8Ek_MlC_OD+D#4FR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNRsbNH_0$L4k#nRR:bHNs0L$_kn#4_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFR8s_FRk05bHMk00RFsR0H0-#N#0C2$
0bFCRkL0_k.#d_b0$C#RHRsNsN5$R80CbEk_MlC_OD-D#4FR8IFM0RRj,dI.*HE80_lMk_DOCDd#+4FR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNR0Fk_#Lkd:.RR0Fk_#Lkd0._$;bCRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFR8s_FRk05bHMk00RFsR0H0-#N#0C2$
0bbCRN0sH$k_L#_d.0C$bRRH#NNss$8R5CEb0_lMk_DOCD4#-RI8FMR0Fjc,R*8IH0ME_kOl_C#DD+8dRF0IMF2RjRRFV#_08DHFoO#;
HNoMDNRbs$H0_#Lkd:.RRsbNH_0$Ldk#.$_0bRC;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RV_Rs80FkRM5HbRk000FRs#H-0CN0##2
HNoMDkRF0M_CR#:R0D8_FOoH_OPC05Fs80CbEk_MlC_OD-D#4FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--CLMNDRC#VRFs0-sH#00NC##
HNoMDsRI0M_CR#:R0D8_FOoH_OPC05Fs80CbEk_MlC_OD-D#4FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--I0sHCMRCNCLD#FRVsNRCOsERFFIRVqR)vCROD
D##MHoNHDRMC_soRR:#_08DHFoOC_POs0F58IH0dE+6FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-#RkC08RFCRso0H#C7sRQ
hR#MHoNFDRks0_C:oRR8#0_oDFHPO_CFO0sH5I8+0Ed86RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-#RkC08RFCRso0H#C7sRm
za#MHoNFDRks0_CRo4:0R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RCk#8FR0RFOEFR#CLIC0CRCM7RQhNRM8Fbk0kF0RVDRAFRO	)
qv#MHoNsDRNs8_C:oRR8#0_oDFHPO_CFO0s85N8HsI8-0E4FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-#RkC08RFCRso0H#C)sRq)77
o#HMRNDI_N8sRCo:0R#8F_Do_HOP0COFNs58I8sHE80-84RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-k-R#RC80sFRC#oH0RCsW7q7)H
#oDMNRIDF_8sN8:sRR8#0_oDFHPO_CFO0sd54RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-R8sN8LsRHR0#HkMb0FR0Rv)qRDOCD5#RcHRL0s#RCHJks2C8
o#HMRNDD_FII8N8sRR:#_08DHFoOC_POs0F5R4d8MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--I8N8sHRL0H#RM0bkRR0F)RqvODCD#cR5R0LH#CRsJskHC
82#MHoN)DRq)77_b0lR#:R0D8_FOoH_OPC05FsNs88I0H8ER-48MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--k8#CRR0FbCHbDCHMR7)q7#)
HNoMDqRW7_7)0Rlb:0R#8F_Do_HOP0COFNs58I8sHE80-84RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-k-R#RC80bFRHDbCHRMCW7q7)H
#oDMNRh7Q_b0lR#:R0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-#RkC08RFHRbbHCDM7CRQ#h
HNoMD RW_b0lR#:R0D8_FOoH;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-k-R#RC80bFRHDbCHRMCW- 
-MRC8DRLFRO	sRNlHDlbCMlC0HN0F#MRHNoMD-#
-CRLoRHM#CCDOs0RNHlRlCbDl0CMNF0HMHR#oDMN#k
VMHO0FoMRCM0_knl_cC58b:0ER0HMCsoC2CRs0MksR0HMCsoCR
H#PHNsNCLDRDPNRH:RMo0CC:sR=;Rj
oLCHRM
RDPNRR:=80CbEc/n;R
RH5VR5b8C0lERFn8Rc>2RR2cURC0EMR
RRNRPD=R:RDPNR4+R;R
RCRM8H
V;RCRs0MksRDPN;M
C8CRo0k_Mlc_n;k
VMHO0FoMRCD0_CFV0P_Csd8.5CEb0RH:RMo0CCRs2skC0sHMRMo0CCHsR#C
Lo
HMRCRs0Mks5b8C0lERFn8Rc
2;CRM8o_C0D0CVFsPC_;d.
MVkOF0HMCRo0C_DVP0FC8s5CEb0RH:RMo0CCRs;lRNG:MRH0CCoss2RCs0kMMRH0CCos#RH
sPNHDNLCNRPDRR:HCM0oRCs:j=R;C
Lo
HMRVRHRC58bR0E-NRlG=R>RRj20MEC
RRRRDPNRR:=80CbERR-l;NG
CRRD
#CRRRRPRND:8=RCEb0;R
RCRM8H
V;RCRs0Mks5DPN2C;
Mo8RCD0_CFV0P;Cs
MVkOF0HMCRo0k_Ml._d5b8C0:ERR0HMCsoC2CRs0MksR0HMCsoCR
H#PHNsNCLDRDPNRH:RMo0CC:sR=;Rj
oLCHRM
RRHV5b8C0<ER=URcR8NMRb8C0>ERR24nRC0EMR
RRPRRN:DR=;R4
CRRMH8RVR;
R0sCkRsMP;ND
8CMR0oC_lMk_;d.
MVkOF0HMCRo0k_Mln_45b8C0:ERR0HMCsoC2CRs0MksR0HMCsoCR
H#PHNsNCLDRDPNRH:RMo0CC:sR=;Rj
oLCHRM
RRHV5b8C0<ER=nR4R8NMRb8C0>ERRRj20MEC
RRRRNRPD=R:R
4;RMRC8VRH;R
RskC0sPMRN
D;CRM8o_C0M_kl4
n;O#FM00NMRlMk_DOCDc_nRH:RMo0CC:sR=CRo0k_Mlc_n5b8C0;E2
MOF#M0N0CRDVP0FCds_.RR:HCM0oRCs:o=RCD0_CFV0P_Csd8.5CEb02O;
F0M#NRM0M_klODCD_Rd.:MRH0CCos=R:R0oC_lMk_5d.D0CVFsPC_2d.;F
OMN#0MD0RCFV0P_Cs4:nRR0HMCsoCRR:=o_C0D0CVFsPC5VDC0CFPs._d,.Rd2O;
F0M#NRM0M_klODCD_R4n:MRH0CCos=R:R0oC_lMk_54nD0CVFsPC_24n;0

$RbCF_k0L_k#0C$b_#ncRRH#NNss$MR5kOl_C_DDn8cRF0IMF,RjR8IH04E-RI8FMR0FjF2RV0R#8F_Do;HO
b0$CkRF0k_L#$_0bdC_.H#R#sRNsRN$5lMk_DOCD._dRI8FMR0FjI,RHE80-84RF0IMF2RjRRFV#_08DHFoO0;
$RbCF_k0L_k#0C$b_#4nRRH#NNss$MR5kOl_C_DD48nRF0IMF,RjR8IH04E-RI8FMR0FjF2RV0R#8F_Do;HO
o#HMRNDF_k0L_k#nRc#:kRF0k_L#$_0bnC_cR#;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RVFR8k50RHkMb0FR0RH0s-N#002C#
o#HMRNDF_k0L_k#dR.#:kRF0k_L#$_0bdC_.R#;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RVFR8k50RHkMb0FR0RH0s-N#002C#
o#HMRNDF_k0L_k#4Rn#:kRF0k_L#$_0b4C_nR#;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RVFR8k50RHkMb0FR0RH0s-N#002C#
o#HMRNDF_k0C#M_R#:R0D8_FOoH_OPC05FsM_klODCD_Rnc8MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-MRCNCLD#FRVssR0H0-#N#0C
o#HMRNDF_k0CdM_.RR:#_08DHFoO#;
HNoMDkRF0M_C_R4n:0R#8F_Do;HO
o#HMRNDI_s0C#M_R#:R0D8_FOoH_OPC05FsM_klODCD_Rnc8MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-sRIHR0CCLMNDRC#VRFsCENORIsFRRFV)RqvODCD#H
#oDMNR0Is__CMd:.RR8#0_oDFH
O;#MHoNIDRsC0_Mn_4R#:R0D8_FOoH;H
#oDMNR_HMs_Co#RR:#_08DHFoOC_POs0F58IH04E-RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RCk#8FR0RosCHC#0sQR7h#R
HNoMDkRF0C_soR_#:0R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-#RkC08RFCRso0H#C7sRm
za#MHoNsDRNs8_C#o_R#:R0D8_FOoH_OPC05FsNs88I0H8ER-48MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--k8#CRR0FsHCo#s0CR7q7)H
#oDMNR8IN_osC_:#RR8#0_oDFHPO_CFO0s85N8HsI8-0E4FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-#RkC08RFCRso0H#CqsR7
7)#MHoNDDRFsI_Ns88_:#RR8#0_oDFHPO_CFO0sR568MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--Ns88R0LH#MRHbRk00)FRqOvRC#DDRR5cL#H0RJsCkCHs8#2
HNoMDFRDIN_I8_8s#RR:#_08DHFoOC_POs0F586RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-N-R8R8sL#H0RbHMk00RFqR)vCRODRD#5LcRHR0#skCJH8sC2-
-R8CMRD#CCRO0sRNlHDlbCMlC0HN0F#MRHNoMDN#
0H0sLCk0Rs\3NFl_VCV#0:\RRs#0H;Mo
C
Lo
HMRRRR-Q-RV8RN8HsI8R0E<EROFCHO_8IH0NER#o#HMjR''FR0RkkM#RC8L#H0
RRRRRzjRH:RVNR58I8sHE80R4=R2CRoMNCs0SC
RRRRD_FIs8N8s=R<Rj"jjjjjjjjjj"jjRs&RNs8_Cjo52S;
RRRRD_FII8N8s=R<Rj"jjjjjjjjjj"jjRI&RNs8_Cjo52S;
CRM8oCCMsCN0R;zj
RRRRRz4RH:RVNR58I8sHE80R.=R2CRoMNCs0SC
SIDF_8sN8<sR=jR"jjjjjjjjj"jjRs&RNs8_C4o5RI8FMR0Fj
2;SRRRRIDF_8IN8<sR=jR"jjjjjjjjj"jjRI&RNs8_C4o5RI8FMR0Fj
2;S8CMRMoCC0sNC4Rz;R
RR.RzRRR:H5VRNs88I0H8ERR=do2RCsMCN
0CSFSDIN_s8R8s<"=Rjjjjjjjjj"jjRs&RNs8_C.o5RI8FMR0Fj
2;SRRRRIDF_8IN8<sR=jR"jjjjjjjjjRj"&NRI8C_soR5.8MFI0jFR2S;
CRM8oCCMsCN0R;z.
RRRRRzdRH:RVNR58I8sHE80Rc=R2CRoMNCs0SC
SIDF_8sN8<sR=jR"jjjjjjjjj&"RR8sN_osC58dRF0IMF2Rj;R
SRDRRFII_Ns88RR<="jjjjjjjj"jjRI&RNs8_Cdo5RI8FMR0Fj
2;S8CMRMoCC0sNCdRz;R
RRcRzRRR:H5VRNs88I0H8ERR=6o2RCsMCN
0CSRRRRIDF_8sN8<sR=jR"jjjjjjjj"RR&s_N8s5CocFR8IFM0R;j2
RSRRFRDIN_I8R8s<"=Rjjjjjjjjj&"RR8IN_osC58cRF0IMF2Rj;C
SMo8RCsMCNR0Cz
c;RRRRzR6R:VRHR85N8HsI8R0E=2RnRMoCC0sNCR
SRDRRFsI_Ns88RR<="jjjjjjjj&"RR8sN_osC586RF0IMF2Rj;S
SD_FII8N8s=R<Rj"jjjjjjRj"&NRI8C_soR568MFI0jFR2S;
CRM8oCCMsCN0R;z6
RRRRRznRH:RVNR58I8sHE80R(=R2CRoMNCs0SC
RRRRD_FIs8N8s=R<Rj"jjjjjj&"RR8sN_osC58nRF0IMF2Rj;S
SD_FII8N8s=R<Rj"jjjjjj&"RR8IN_osC58nRF0IMF2Rj;C
SMo8RCsMCNR0Cz
n;RRRRzR(R:VRHR85N8HsI8R0E=2RURMoCC0sNCR
SRDRRFsI_Ns88RR<="jjjj"jjRs&RNs8_C(o5RI8FMR0Fj
2;SFSDIN_I8R8s<"=RjjjjjRj"&NRI8C_soR5(8MFI0jFR2S;
CRM8oCCMsCN0R;z(
RRRRRzURH:RVNR58I8sHE80Rg=R2CRoMNCs0SC
RRRRD_FIs8N8s=R<Rj"jj"jjRs&RNs8_CUo5RI8FMR0Fj
2;SFSDIN_I8R8s<"=Rjjjjj&"RR8IN_osC58URF0IMF2Rj;C
SMo8RCsMCNR0Cz
U;RRRRzRgR:VRHR85N8HsI8R0E=jR42CRoMNCs0SC
RRRRD_FIs8N8s=R<Rj"jjRj"&NRs8C_soR5g8MFI0jFR2S;
SIDF_8IN8<sR=jR"j"jjRI&RNs8_Cgo5RI8FMR0Fj
2;S8CMRMoCC0sNCgRz;R
RR4Rzj:RRRRHV58N8s8IH0=ERR244RMoCC0sNCR
SRDRRFsI_Ns88RR<="jjj"RR&s_N8s5Co48jRF0IMF2Rj;S
SD_FII8N8s=R<Rj"jj&"RR8IN_osC5R4j8MFI0jFR2S;
CRM8oCCMsCN0Rjz4;R
RR4Rz4:RRRRHV58N8s8IH0=ERR24.RMoCC0sNCR
SRDRRFsI_Ns88RR<=""jjRs&RNs8_C4o54FR8IFM0R;j2
DSSFII_Ns88RR<=""jjRI&RNs8_C4o54FR8IFM0R;j2
MSC8CRoMNCs0zCR4
4;RRRRzR4.RH:RVNR58I8sHE80R4=Rdo2RCsMCN
0CSRRRRIDF_8sN8<sR=jR''RR&s_N8s5Co48.RF0IMF2Rj;S
SD_FII8N8s=R<R''jRI&RNs8_C4o5.FR8IFM0R;j2
MSC8CRoMNCs0zCR4
.;RRRRzR4dRH:RVNR58I8sHE80R4>Rdo2RCsMCN
0CSRRRRIDF_8sN8<sR=NRs8C_sod54RI8FMR0Fj
2;SRRRRIDF_8IN8<sR=NRI8C_sod54RI8FMR0Fj
2;S8CMRMoCC0sNC4Rzd
;
RRRR-Q-RV8R5HsM_CRo2sHCo#s0CRh7QRHk#MBoRpRi
RzRR4RcR:VRHRH58MC_soo2RCsMCN
0CRRRRRRRRbOsFCR##5iBp,QR7hL2RCMoH
RRRRRRRRRRRRRHV5iBpR'=R4N'RMB8RpCi'P0CM2ER0CRM
RRRRRRRRRRRRRHRRMC_so=R<Rj5"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jjR7&RQ;h2
RRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMRFbsO#C#;C
SMo8RCsMCNR0Cz;4c
RRRR6z4RRR:H5VRMRF08_HMs2CoRMoCC0sNCR
RRRRRRRRRRMRH_osCRR<=5j"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjRj"&QR7h
2;S8CMRMoCC0sNC4Rz6
;
RRRR7amzRR<=F_k0s5CoI0H8ER-48MFI0jFR2
;
RRRR-Q-RVsR5Ns88_osC2CRso0H#C)sRq)77RHk#MmoRB
piRRRRzs4nRRR:H5VRs8N8sC_soo2RCsMCN
0C-R-RRRRRRsRbF#OC#mR5B,piR7)q7R)2LHCoM-
-RRRRRRRRRRRRH5VRmiBpR'=R4N'RMm8RB'piCMPC002RE
CM-R-RRRRRRRRRRRRRRNRs8C_so=R<R7)q7N)58I8sHE80-84RF0IMF2Rj;-
-RRRRRRRRRRRRCRM8H
V;-R-RRRRRRMRC8sRbF#OC#-;
-MSC8CRoMNCs0zCR4;ns
R--RzRR4R(s:VRHRF5M0NRs8_8ss2CoRMoCC0sNCR
RRRRRRRRRRNRs8C_so=R<R7)q7
);S8CMRMoCC0sNC4Rzn
s;
-S-RRQV58IN8ss_CRo2sHCo#s0CR7Wq7k)R#oHMRmW_B
piRRRRzI4nRRR:H5VRI8N8sC_soo2RCsMCN
0CRRRRRRRRbOsFCR##5iBp,qRW727)RoLCHRM
RRRRRRRRRHRRVBR5p=iRR''4R8NMRiBp'CCPMR020MEC
RRRRRRRRRRRRRRRR8IN_osCRR<=W7q7)85N8HsI8-0E4FR8IFM0R;j2
RRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMRFbsO#C#;C
SMo8RCsMCNR0CzI4n;R
RR4Rz(:IRRRHV50MFR8IN8ss_CRo2oCCMsCN0
RRRRRRRRRRRR8IN_osCRR<=W7q7)S;
CRM8oCCMsCN0R(z4I
;
RRRR-t-RCsMCNR0C0REC)RqvODCD#MRN8CR#D0CORoDFHVORF)sRq4vAn4_1_
14SUz4RH:RVOR5EOFHCH_I8R0E=2R4RMoCC0sNCR
RRzRS4:gRRsVFRHHRM8R5CEb0_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNC-
S-VRQR85N8HsI8R0E>cR42CRMC08RFsROCCN0RHIs0CCRMDNLCMRN8kRF00bkRNCMLRDC#CCDOD0RFOoH
RRRRRRRR.SzjRR:H5VRNs88I0H8ERR>4Rc2oCCMsCN0
-S-RGVHRsVFRDONDdR4U,U(RD#CCRO0F0VRs0H#NR0CMRF0LMCHoCRso0H#C8sC
SSSS0Fk_5CMH<2R=4R''ERIC5MRs_N8s5CoNs88I0H8ER-48MFI04FRc=2RRRH2CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R ERIC5MRI_N8s5CoNs88I0H8ER-48MFI04FRc=2RRRH2CCD#R''j;R
RRRRRRCRSMo8RCsMCNR0Cz;.j
-S-RRQV58N8s8IH0<ER=cR42FRMRHIs0CCRMDNLCsRFR0FkbRk0CLMND#CRCODC0FRDoRHOM8CCCR8
SRRRR.Sz4RR:H5VRNs88I0H8E=R<R24cRMoCC0sNCS
SSkSF0M_C5RH2<'=R4
';RRRRRRRRRRRRRRRRI_s0CHM52=R<R;W 
RRRRRRRRMSC8CRoMNCs0zCR.
4;SR--tCCMsCN0RC0ERv)qRDOCDN#RM08Rs#H-0CN0#R
RRRRRRzRS.:.RRsVFRH[RMIR5HE80_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNCS
SS0N0skHL0GCROs_bFRb#FAVR)_qv4Undc7X4RD:RNDLCRRH#"QW)av _m_7 q =)qw7_Qa)1,)R1e_qpAR="&sR#P5ND[2+4R"&R,)RWQ_a v m7_"A=RI&RsF_l8
C;RRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FAVR)_qv4Undc7X4RD:RNDLCRRH#"aA7"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloHC5*d4nURc2&WR""RR&HCM0o'CsHolNC25[R"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05R5H+2R4*d4nURc,80CbER22&XR""RR&HCM0o'CsHolNC+5[4
2;SLSSCMoH
RRRRRRRRRRRR)SAq4v_ncdUXR47:qR)vnA4__141S4
RRRRRRRRRRRRb0FsRblNRQ57q25jRR=>HsM_C[o52q,R7q7)RR=>D_FII8N8sd54RI8FMR0FjR2,7RQA=">RjR",q)77A>R=RIDF_8sN84s5dFR8IFM0R,j2
SSSSq hRR=>Wh_ ,1R1)=qR>jR''W,R =qR>sRI0M_C5,H2RiBpq>R=RiBp,hR A>R=R, hR)11A>R=Ra)1, RWA>R=R''j,pRBi=AR>BRmp
i,SRSSR7RRm=qR>bRFCRM,75mAj=2R>kRF0k_L#H45,2[2;R

RRRRRRRRRRRRRFRRks0_C[o52=R<R0Fk_#Lk4,5H[I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRS8CMRMoCC0sNC.Rz.R;
RRRRS8CMRMoCC0sNC4RzgR;
RCRRMo8RCsMCNR0Cz;4URRRR
RRRR
RRRRRR-t-RCsMCNR0C0REC)RqvODCD#MRN8CR#D0CORoDFHVORF)sRq4vAn._1_
1.Sdz.RH:RVOR5EOFHCH_I8R0E=2R.RMoCC0sNCR
RRzRS.:cRRsVFRHHRM8R5CEb0_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNC-
S-VRQR85N8HsI8R0E>dR42CRMC08RFsROCCN0RHIs0CCRMDNLCMRN8kRF00bkRNCMLRDC#CCDOD0RFOoH
RRRRRRRR.Sz6RR:H5VRNs88I0H8ERR>4Rd2oCCMsCN0
-S-RGVHRsVFRDONDdR4U,U(RD#CCRO0F0VRs0H#NR0CMRF0LMCHoCRso0H#C8sC
RRRRRRRRRRRRRRRR0Fk_5CMH<2R=4R''ERIC5MRs_N8s5CoNs88I0H8ER-48MFI04FRd=2RRRH2CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R ERIC5MRI_N8s5CoNs88I0H8ER-48MFI04FRd=2RRRH2CCD#R''j;R
RRRRRRCRSMo8RCsMCNR0Cz;.6
-S-RRQV58N8s8IH0<ER=dR42FRMRHIs0CCRMDNLCsRFR0FkbRk0CLMND#CRCODC0FRDoRHOM8CCCR8
SRRRR.SznRR:H5VRNs88I0H8E=R<R24dRMoCC0sNCR
SRRRRRRRRRFRRkC0_M25HRR<=';4'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RW;R
RRRRRRCRSMo8RCsMCNR0Cz;.n
-S-RMtCC0sNCER0CqR)vCRODRD#NRM80-sH#00NCR#
RRRRRSRRzR.(:FRVsRR[H5MRI0H8Ek_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0SC
S0SN0LsHkR0CGbO_s#FbRRFVAv)q_gU4.7X.RD:RNDLCRRH#"QW)av _m_7 q =)qw7_Qa)1,)R1e_qpAR="&sR#P5ND.+*[.FR8IFM0R[.*+R42&,R"RQW)av _m_7 AR="&sRI_8lFCR;
RRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)RAqUv_4Xg..:7RRLDNCHDR#AR"7Ra"&MRH0CCosl'HN5oCI0H8E&2RR""7RH&RMo0CCHs'lCNo5UH*42g.R"&RW&"RR0HMCsoC'NHlo[C5*R.2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50E5+HRR*42U.4g,CR8b20E2RR&"RX"&MRH0CCosl'HN5oC54[+22*.;S
SSoLCHRM
RRRRRRRRRSRRAv)q_gU4.7X.R):Rq4vAn._1_
1.SRRRRRRRRRRRRsbF0NRlb7R5Q=qR>MRH_osC5[.*+84RF0IMF*R.[R2,q)77q>R=RIDF_8IN84s5.FR8IFM0R,j2RA7QRR=>""jj,7Rq7R)A=D>RFsI_Ns885R4.8MFI0jFR2S,
SRSRRhR q>R=R W_h1,R1R)q='>RjR',WR q=I>RsC0_M25H,pRBi=qR>pRBi ,Rh=AR>hR ,1R1)=AR>1R)aW,R =AR>jR''B,RpRiA=m>RB,pi
SSSRRRR7Rmq=F>Rb,CMRA7m5R42=F>RkL0_k5#.H*,.[2+4,mR7A25jRR=>F_k0L.k#5RH,.2*[2R;
RRRRRRRRRRRRRFRRks0_C.o5*R[2<F=RkL0_k5#.H*,.[I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co.+*[4<2R=kRF0k_L#H.5,[.*+R42IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRMSC8CRoMNCs0zCR.
(;RRRRRMSC8CRoMNCs0zCR.
c;RRRRCRM8oCCMsCN0Rdz.;
RR
RSRR-R-RMtCC0sNCER0CqR)vCRODRD#NRM8#CCDOD0RFOoHRsVFRv)qA_4n11c_cz
S.:URRRHV5FOEH_OCI0H8ERR=co2RCsMCN
0CRRRRSgz.RV:RFHsRRRHM5b8C0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CSR--Q5VRNs88I0H8ERR>4R.2M8CCRR0FONsC0ICRsCH0RNCMLRDCNRM8Fbk0kC0RMDNLCCR#D0CORoDFHRO
RRRRRSRRzRdj:VRHR85N8HsI8R0E>.R42CRoMNCs0SC
-V-RHVGRFOsRNRDD4UdU(#,RCODC0VRFRH0s#00NCFRM0CRLHRMosHCo#s0CCR8
RRRRRRRRRRRRRFRRkC0_M25HRR<='R4'IMECRN5s8C_so85N8HsI8-0E4FR8IFM0R24.RH=R2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0CHM52=R<RRW IMECRN5I8C_so85N8HsI8-0E4FR8IFM0R24.RH=R2DRC#'CRj
';RRRRRRRRS8CMRMoCC0sNCdRzjS;
-Q-RVNR58I8sHE80RR<=4R.2MIFRsCH0RNCMLRDCFFsRkk0b0MRCNCLDRD#CCRO0DHFoOCRMC88C
RRSRSRRzRd4:VRHR85N8HsI8R0E<4=R.o2RCsMCN
0CSSSSF_k0CHM52=R<R''4;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R R;
RRRRRSRRCRM8oCCMsCN0R4zd;-
S-CRtMNCs00CRE)CRqOvRC#DDR8NMRH0s-N#00
C#RRRRRRRRS.zdRV:RF[sRRRHM58IH0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CSNSS0H0sLCk0R_GObbsF#VRFRqA)vj_cgcnX7RR:DCNLD#RHR)"WQ_a v m7_)q= _q7w1Q)a1,R)peq_"A=R#&RsDPN5[c*+8cRF0IMF*Rc[2+4R"&R,)RWQ_a v m7_"A=RI&RsF_l8
C;RRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FAVR)_qvcnjgXRc7:NRDLRCDH"#RA"7aRH&RMo0CCHs'lCNo58IH0RE2&7R""RR&HCM0o'CsHolNC*5Hcnjg2RR&"RW"&MRH0CCosl'HN5oC[2*cR"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05R5H+2R4*gcjn8,RCEb02&2RR""XRH&RMo0CCHs'lCNo5+5[4c2*2S;
SCSLo
HMRRRRRRRRRRRRSqA)vj_cgcnX7RR:)Aqv41n_cc_1
RSRRRRRRRRRRFRbsl0RN5bR7RQq=H>RMC_so*5c[R+d8MFI0cFR*,[2R7q7)=qR>FRDIN_I858s484RF0IMF2Rj,QR7A>R=Rj"jj,j"R7q7)=AR>FRDIN_s858s484RF0IMF2Rj,S
SShS q>R=R W_h1,R1R)q='>RjR',WR q=I>RsC0_M25H,pRBi=qR>pRBi ,Rh=AR>hR ,1R1)=AR>1R)aW,R =AR>jR''B,RpRiA=m>RB,pi
SSSSq7mRR=>FMbC,mR7A25dRR=>F_k0Lck#5RH,c+*[dR2,75mA.=2R>kRF0k_L#Hc5,[c*+,.2RS
SSmS7A254RR=>F_k0Lck#5cH,*4[+27,RmjA52>R=R0Fk_#Lkc,5HR[c*2
2;RRRRRRRRRRRRRRRRF_k0s5Coc2*[RR<=F_k0Lck#5cH,*R[2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5[c*+R42<F=RkL0_k5#cH*,c[2+4RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so*5c[2+.RR<=F_k0Lck#5cH,*.[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cco5*d[+2=R<R0Fk_#Lkc,5Hc+*[dI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';
RRRRRRRRMSC8CRoMNCs0zCRd
.;RRRRRMSC8CRoMNCs0zCR.
g;RRRRCRM8oCCMsCN0RUz.;S

RRRR-t-RCsMCNR0C0REC)RqvODCD#MRN8CR#D0CORoDFHVORF)sRq4vAng_1_
1gSdzdRH:RVOR5EOFHCH_I8R0E=2RgRMoCC0sNCR
RRzRSd:cRRsVFRHHRM8R5CEb0_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNC-
S-VRQR85N8HsI8R0E>4R42CRMC08RFsROCCN0RHIs0CCRMDNLCMRN8kRF00bkRNCMLRDC#CCDOD0RFOoH
RRRRRRRRdSz6RR:H5VRNs88I0H8ERR>4R42oCCMsCN0
-S-RGVHRsVFRDONDdR4U,U(RD#CCRO0F0VRs0H#NR0CMRF0LMCHoCRso0H#C8sC
RRRRRRRRRRRRRRRR0Fk_5CMH<2R=4R''ERIC5MRs_N8s5CoNs88I0H8ER-48MFI04FR4=2RRRH2CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R ERIC5MRI_N8s5CoNs88I0H8ER-48MFI04FR4=2RRRH2CCD#R''j;R
RRRRRRCRSMo8RCsMCNR0Cz;d6
-S-RRQV58N8s8IH0<ER=4R42FRMRHIs0CCRMDNLCsRFR0FkbRk0CLMND#CRCODC0FRDoRHOM8CCCR8
SRRRRdSznRR:H5VRNs88I0H8E=R<R244RMoCC0sNCR
SRRRRRRRRRFRRkC0_M25HRR<=';4'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RW;R
RRRRRRCRSMo8RCsMCNR0Cz;dn
-S-RMtCC0sNCER0CqR)vCRODRD#NRM80-sH#00NCR#
RRRRRSRRzRd(:FRVsRR[H5MRI0H8Ek_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0SC
S0SN0LsHkR0CGbO_s#FbRRFVAv)q_c.jU7XURD:RNDLCRRH#"QW)av _m_7 q =)qw7_Qa)1,)R1e_qpAR="&sR#P5NDg+*[gFR8IFM0R[g*+R42&,R"RQW)av _m_7 AR="&sRI_8lFCR;
RRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)RAq.v_jXcUU:7RRLDNCHDR#AR"7Ra"&MRH0CCosl'HN5oCI0H8E&2RR""7RH&RMo0CCHs'lCNo5.H*j2cUR"&RW&"RR0HMCsoC'NHlo[C5*Rg2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50E5+HRR*42.Ujc,CR8b20E2RR&"RX"&MRH0CCosl'HN5oC54[+22*g;S
SSoLCHRM
RRRRRRRRRSRRAv)q_c.jU7XUR):Rq4vAng_1_
1gRRRRRRRRRRRRRRRRRFRbsl0RN5bR7RQq=H>RMC_so*5g[R+(8MFI0gFR*,[2R7q7)=qR>FRDIN_I858s48jRF0IMF2Rj,QR7A>R=Rj"jjjjjj,j"R7q7)=AR>FRDIN_s858s48jRF0IMF2Rj,R
RRRRRRRRRRRRRRRRRRRRRRRRRRhR q>R=R W_h1,R1R)q='>RjR',WR q=I>RsC0_M25H,pRBi=qR>pRBi ,Rh=AR>hR ,1R1)=AR>1R)aW,R =AR>jR''B,RpRiA=m>RB,piRR
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7q>R=RCFbM7,Rm(A52>R=R0Fk_#LkU,5HU+*[(R2,75mAn=2R>kRF0k_L#HU5,[U*+,n2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7A256RR=>F_k0LUk#5UH,*6[+27,RmcA52>R=R0Fk_#LkU,5HU+*[cR2,75mAd=2R>kRF0k_L#HU5,[U*+,d2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7A25.RR=>F_k0LUk#5UH,*.[+27,Rm4A52>R=R0Fk_#LkU,5HU+*[4R2,75mAj=2R>kRF0k_L#HU5,[U*2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRR7qQu5Rj2=H>RMC_so*5g[2+U,QR7u=AR>jR""R,
RRRRRRRRRRRRRRRRRRRRRRRRR7RRmRuq=F>Rb,CMRu7mA25jRR=>bHNs0L$_k5#UH2,[2R;
RRRRRRRRRRRRRFRRks0_Cgo5*R[2<F=RkL0_k5#UH*,U[I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cog+*[4<2R=kRF0k_L#HU5,[U*+R42IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5[g*+R.2<F=RkL0_k5#UH*,U[2+.RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so*5g[2+dRR<=F_k0LUk#5UH,*d[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cgo5*c[+2=R<R0Fk_#LkU,5HU+*[cI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cog+*[6<2R=kRF0k_L#HU5,[U*+R62IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5[g*+Rn2<F=RkL0_k5#UH*,U[2+nRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so*5g[2+(RR<=F_k0LUk#5UH,*([+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cgo5*U[+2=R<RsbNH_0$LUk#5[H,2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRSRRCRM8oCCMsCN0R(zd;R
RRSRRCRM8oCCMsCN0Rczd;R
RRMRC8CRoMNCs0zCRd
d;
RSRR-R-RMtCC0sNCER0CqR)vCRODRD#NRM8#CCDOD0RFOoHRsVFRv)qA_4n1_4U1
4USUzdRH:RVOR5EOFHCH_I8R0E=UR42CRoMNCs0RC
RSRRzRdg:FRVsRRHH5MR80CbEk_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0SC
-Q-RVNR58I8sHE80R4>RjM2RCRC80OFRs0CNCsRIHR0CCLMNDNCRMF8Rkk0b0MRCNCLDRD#CCRO0DHFoOR
RRRRRRzRSc:jRRRHV58N8s8IH0>ERR24jRMoCC0sNC-
S-HRVGFRVsNROD4DRd(UU,CR#D0CORRFV0#sH0CN0R0MFRHLCMsoRC#oH0CCs8R
RRRRRRRRRRRRRRkRF0M_C5RH2<'=R4I'RERCM58sN_osC58N8s8IH04E-RI8FMR0F4Rj2=2RHR#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=WI RERCM58IN_osC58N8s8IH04E-RI8FMR0F4Rj2=2RHR#CDCjR''R;
RRRRRSRRCRM8oCCMsCN0Rjzc;-
S-VRQR85N8HsI8R0E<4=RjM2RFsRIHR0CCLMNDFCRskRF00bkRNCMLRDC#CCDOD0RFOoHRCMC8
C8RRSRRzRSc:4RRRHV58N8s8IH0<ER=jR42CRoMNCs0SC
RRRRRRRRRRRRF_k0CHM52=R<R''4;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R R;
RRRRRSRRCRM8oCCMsCN0R4zc;-
S-CRtMNCs00CRE)CRqOvRC#DDR8NMRH0s-N#00
C#RRRRRRRRS.zcRV:RF[sRRRHM58IH0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CSNSS0H0sLCk0R_GObbsF#VRFRqA)vj_4.4cXn:7RRLDNCHDR#WR") Qa_7vm =_q)7 q_)wQ1Ra,1q)ep=_A"RR&#NsPDU54*4[+UFR8IFM0R*4U[2+4R"&R,)RWQ_a v m7_"A=RI&RsF_l8
C;RRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FAVR)_qv4cj.X74nRD:RNDLCRRH#"aA7"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloHC5*.4jc&2RR""WRH&RMo0CCHs'lCNo54[*U&2RR"" RH&RMo0CCHs'lCNo50oC_8CM_b8C05E5HRR+442*j,.cRb8C02E2R"&RX&"RR0HMCsoC'NHlo5C5[2+4*24U;S
SSoLCHRM
RRRRRRRRRSRRAv)q_.4jcnX47RR:)Aqv41n_41U_4RU
RRRRRRRRRRRRRRRRRsbF0NRlb7R5Q=qR>MRH_osC5*4U[6+4RI8FMR0F4[U*2q,R7q7)RR=>D_FII8N8sR5g8MFI0jFR27,RQ=AR>jR"jjjjjjjjjjjjj"jj,7Rq7R)A=D>RFsI_Ns8858gRF0IMF2Rj,R
RRRRRRRRRRRRRRRRRRRRRRRRRRhR q>R=R W_h1,R1R)q='>RjR',WR q=I>RsC0_M25H,pRBi=qR>pRBi ,Rh=AR>hR ,1R1)=AR>1R)aW,R =AR>jR''B,RpRiA=m>RB,piRR
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7q>R=RCFbM7,Rm4A56=2R>kRF0k_L#54nHn,4*4[+6R2,75mA4Rc2=F>RkL0_kn#454H,n+*[4,c2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7Ad542>R=R0Fk_#Lk4Hn5,*4n[d+427,Rm4A5.=2R>kRF0k_L#54nHn,4*4[+.R2,75mA4R42=F>RkL0_kn#454H,n+*[4,42RR
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7Aj542>R=R0Fk_#Lk4Hn5,*4n[j+427,RmgA52>R=R0Fk_#Lk4Hn5,*4n[2+g,mR7A25URR=>F_k0L4k#n,5H4[n*+,U2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7A25(RR=>F_k0L4k#n,5H4[n*+,(2RA7m5Rn2=F>RkL0_kn#454H,n+*[nR2,75mA6=2R>kRF0k_L#54nHn,4*6[+2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mAc=2R>kRF0k_L#54nHn,4*c[+27,RmdA52>R=R0Fk_#Lk4Hn5,*4n[2+d,mR7A25.RR=>F_k0L4k#n,5H4[n*+,.2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7A254RR=>F_k0L4k#n,5H4[n*+,42RA7m5Rj2=F>RkL0_kn#454H,n2*[,RR
RRRRRRRRRRRRRRRRRRRRRRRRR7RRQRuq=H>RMC_soU54*4[+(FR8IFM0R*4U[n+427,RQRuA=">Rj,j"Ru7mq>R=RCFbMR,
RRRRRRRRRRRRRRRRRRRRRRRRR7RRm5uA4=2R>NRbs$H0_#Lk4Hn5,[.*+,42Ru7mA25jRR=>bHNs0L$_kn#45.H,*2[2;R
RRRRRRRRRRRRRRkRF0C_soU54*R[2<F=RkL0_kn#454H,n2*[RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*4[+2=R<R0Fk_#Lk4Hn5,*4n[2+4RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*.[+2=R<R0Fk_#Lk4Hn5,*4n[2+.RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*d[+2=R<R0Fk_#Lk4Hn5,*4n[2+dRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*c[+2=R<R0Fk_#Lk4Hn5,*4n[2+cRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*6[+2=R<R0Fk_#Lk4Hn5,*4n[2+6RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*n[+2=R<R0Fk_#Lk4Hn5,*4n[2+nRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*([+2=R<R0Fk_#Lk4Hn5,*4n[2+(RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*U[+2=R<R0Fk_#Lk4Hn5,*4n[2+URCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*g[+2=R<R0Fk_#Lk4Hn5,*4n[2+gRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*4[+j<2R=kRF0k_L#54nHn,4*4[+jI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+244RR<=F_k0L4k#n,5H4[n*+244RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*4[+.<2R=kRF0k_L#54nHn,4*4[+.I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+24dRR<=F_k0L4k#n,5H4[n*+24dRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*4[+c<2R=kRF0k_L#54nHn,4*4[+cI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+246RR<=F_k0L4k#n,5H4[n*+246RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*4[+n<2R=NRbs$H0_#Lk4Hn5,[.*2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[4R(2<b=RN0sH$k_L#54nH*,.[2+4RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R

RRRRRSRRCRM8oCCMsCN0R.zc;R
RRSRRCRM8oCCMsCN0Rgzd;R
RRMRC8CRoMNCs0zCRd
U;
RSRR-R-RMtCC0sNCER0CqR)vCRODRD#NRM8#CCDOD0RFOoHRsVFRv)qA_4n1_dn1
dnSUzdNRR:H5VROHEFOIC_HE80Rd=Rno2RCsMCN
0CSRRRRgzdNRR:VRFsHMRHRC58b_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
-S-RRQV58N8s8IH0>ERRRg2M8CCRR0FONsC0ICRsCH0RNCMLRDCNRM8Fbk0kC0RMDNLCCR#D0CORoDFHSO
ScSzj:NRRRHV58N8s8IH0>ERRRg2oCCMsCN0
-S-RGVHRsVFRDONDdR4U,U(RD#CCRO0F0VRs0H#NR0CMRF0LMCHoCRso0H#C8sC
SSSS0Fk_5CMH<2R=4R''ERIC5MRs_N8s5CoNs88I0H8ER-48MFI0gFR2RR=HC2RDR#C';j'
SSSS0Is_5CMH<2R= RWRCIEMIR5Ns8_CNo58I8sHE80-84RF0IMF2RgRH=R2DRC#'CRj
';SCSSMo8RCsMCNR0CzNcj;-
S-VRQR85N8HsI8R0E<g=R2FRMRHIs0CCRMDNLCsRFR0FkbRk0CLMND#CRCODC0FRDoRHOM8CCCS8
ScSz4:NRRRHV58N8s8IH0<ER=2RgRMoCC0sNCS
SSkSF0M_C5RH2<'=R4
';SSSSI_s0CHM52=R<R;W 
SSSCRM8oCCMsCN0R4zcNS;
-t-RCsMCNR0C0REC)RqvODCD#MRN8sR0H0-#N#0C
SSSzNc.RV:RF[sRRRHM58IH0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CSNSS0H0sLCk0R_GObbsF#VRFRqA)v4_6..Xd7RR:DCNLD#RHR)"WQ_a v m7_)q= _q7w1Q)a1,R)peq_"A=R#&RsDPN5*dn[n+dRI8FMR0Fd[n*+R42&,R"RQW)av _m_7 AR="&sRI_8lFCR;
RRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)RAq6v_4d.X.:7RRLDNCHDR#AR"7Ra"&MRH0CCosl'HN5oCI0H8E&2RR""7RH&RMo0CCHs'lCNo56H*4R.2&WR""RR&HCM0o'CsHolNC*5[dRn2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50E5+HRR*426,4.Rb8C02E2R"&RX&"RR0HMCsoC'NHlo5C5[2+4*2dn;S
SSoLCHRM
RRRRRRRRRRRRRRRRRRRRRRRRRqA)v4_6..Xd7RR:)Aqv41n_d1n_dRn
RRRRRRRRRRRRRRRRRRRRRRRRRbRRFRs0lRNb5q7QRR=>HsM_Cdo5n+*[d84RF0IMFnRd*,[2R7q7)=qR>FRDIN_I858sUFR8IFM0R,j2RA7QRR=>"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjR",q)77A>R=RIDF_8sN8Us5RI8FMR0Fj
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRhR q>R=R W_h1,R1R)q='>RjR',WR q=I>RsC0_M25H,pRBi=qR>pRBi ,Rh=AR>hR ,1R1)=AR>1R)aW,R =AR>jR''B,RpRiA=m>RB,pi
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRm=qR>bRFCRM,75mAdR42=F>RkL0_k.#d5dH,.+*[d,42RA7m52djRR=>F_k0Ldk#.,5Hd[.*+2dj,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mA.Rg2=F>RkL0_k.#d5dH,.+*[.,g2RA7m52.URR=>F_k0Ldk#.,5Hd[.*+2.U,mR7A(5.2>R=R0Fk_#LkdH.5,*d.[(+.2R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRA7m52.nRR=>F_k0Ldk#.,5Hd[.*+2.n,mR7A65.2>R=R0Fk_#LkdH.5,*d.[6+.27,Rm.A5c=2R>kRF0k_L#5d.H.,d*.[+c
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7Ad5.2>R=R0Fk_#LkdH.5,*d.[d+.27,Rm.A5.=2R>kRF0k_L#5d.H.,d*.[+.R2,75mA.R42=F>RkL0_k.#d5dH,.+*[.,42
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRm.A5j=2R>kRF0k_L#5d.H.,d*.[+jR2,75mA4Rg2=F>RkL0_k.#d5dH,.+*[4,g2RA7m524URR=>F_k0Ldk#.,5Hd[.*+24U,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mA4R(2=F>RkL0_k.#d5dH,.+*[4,(2RA7m524nRR=>F_k0Ldk#.,5Hd[.*+24n,mR7A6542>R=R0Fk_#LkdH.5,*d.[6+42R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRA7m524cRR=>F_k0Ldk#.,5Hd[.*+24c,mR7Ad542>R=R0Fk_#LkdH.5,*d.[d+427,Rm4A5.=2R>kRF0k_L#5d.H.,d*4[+.
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7A4542>R=R0Fk_#LkdH.5,*d.[4+427,Rm4A5j=2R>kRF0k_L#5d.H.,d*4[+jR2,75mAg=2R>kRF0k_L#5d.H.,d*g[+2R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRA7m5RU2=F>RkL0_k.#d5dH,.+*[UR2,75mA(=2R>kRF0k_L#5d.H.,d*([+27,RmnA52>R=R0Fk_#LkdH.5,*d.[2+n,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mA6=2R>kRF0k_L#5d.H.,d*6[+27,RmcA52>R=R0Fk_#LkdH.5,*d.[2+c,mR7A25dRR=>F_k0Ldk#.,5Hd[.*+,d2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRm.A52>R=R0Fk_#LkdH.5,*d.[2+.,mR7A254RR=>F_k0Ldk#.,5Hd[.*+,42RA7m5Rj2=F>RkL0_k.#d5dH,.2*[,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR7qQuRR=>HsM_Cdo5n+*[d86RF0IMFnRd*d[+.R2,7AQuRR=>"jjjjR",7qmuRR=>FMbC,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR7Amu5Rd2=b>RN0sH$k_L#5d.H*,c[2+d,mR7u.A52>R=RsbNH_0$Ldk#.,5Hc+*[.
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7u4A52>R=RsbNH_0$Ldk#.,5Hc+*[4R2,7Amu5Rj2=b>RN0sH$k_L#5d.H*,c[;22
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n2*[RR<=F_k0Ldk#.,5Hd[.*2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[2+4RR<=F_k0Ldk#.,5Hd[.*+R42IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[.<2R=kRF0k_L#5d.H.,d*.[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[2+dRR<=F_k0Ldk#.,5Hd[.*+Rd2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[c<2R=kRF0k_L#5d.H.,d*c[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[2+6RR<=F_k0Ldk#.,5Hd[.*+R62IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[n<2R=kRF0k_L#5d.H.,d*n[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[2+(RR<=F_k0Ldk#.,5Hd[.*+R(2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[U<2R=kRF0k_L#5d.H.,d*U[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[2+gRR<=F_k0Ldk#.,5Hd[.*+Rg2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[4Rj2<F=RkL0_k.#d5dH,.+*[4Rj2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[4R42<F=RkL0_k.#d5dH,.+*[4R42IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[4R.2<F=RkL0_k.#d5dH,.+*[4R.2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[4Rd2<F=RkL0_k.#d5dH,.+*[4Rd2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[4Rc2<F=RkL0_k.#d5dH,.+*[4Rc2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[4R62<F=RkL0_k.#d5dH,.+*[4R62IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[4Rn2<F=RkL0_k.#d5dH,.+*[4Rn2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[4R(2<F=RkL0_k.#d5dH,.+*[4R(2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[4RU2<F=RkL0_k.#d5dH,.+*[4RU2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[4Rg2<F=RkL0_k.#d5dH,.+*[4Rg2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[.Rj2<F=RkL0_k.#d5dH,.+*[.Rj2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[.R42<F=RkL0_k.#d5dH,.+*[.R42IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[.R.2<F=RkL0_k.#d5dH,.+*[.R.2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[.Rd2<F=RkL0_k.#d5dH,.+*[.Rd2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[.Rc2<F=RkL0_k.#d5dH,.+*[.Rc2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[.R62<F=RkL0_k.#d5dH,.+*[.R62IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[.Rn2<F=RkL0_k.#d5dH,.+*[.Rn2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[.R(2<F=RkL0_k.#d5dH,.+*[.R(2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[.RU2<F=RkL0_k.#d5dH,.+*[.RU2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[.Rg2<F=RkL0_k.#d5dH,.+*[.Rg2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[dRj2<F=RkL0_k.#d5dH,.+*[dRj2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[dR42<F=RkL0_k.#d5dH,.+*[dR42IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[dR.2<b=RN0sH$k_L#5d.H*,c[I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*d[+d<2R=NRbs$H0_#LkdH.5,[c*+R42IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[dRc2<b=RN0sH$k_L#5d.H*,c[2+.RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*+2d6RR<=bHNs0L$_k.#d5cH,*d[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''
;
SCSSMo8RCsMCNR0CzNc.;S
SCRM8oCCMsCN0RgzdNS;
CRM8oCCMsCN0RUzdN
;
CRM8NEsOHO0C0CksRFLDOs	_N
l;
ONsECH0Os0kCFRM__sIOOEC	VRFRv)qh__)W#RH
MVkOF0HMkRVMHO_M5H0LRR:LDFFC2NMR0sCkRsM#H0sMHoR#C
Lo
HMRVRHR25LRC0EMR
RRCRs0Mks5F"hRNsC8s/IHR0COVFMD0HORCOEOR	31kHlDHN0FlMRHN#l0ROEb#F#HCLDR"!!2R;
R#CDCR
RRCRs0Mks5F"BkRD8MRF0HDlbCMlC0DRAFRO	)3qvRRQ#0RECs8CNR8N8s#C#RosCHC#0sRC8kM#HoER0CNR#lOCRD	FORRN#0REC)?qv"
2;RMRC8VRH;M
C8kRVMHO_M;H0
MVkOF0HMCRo0M_C8C_8b50E#CHxRH:RMo0CC;sRRb8C0:ERR0HMCsoC2CRs0MksR0HMCsoCR
H#PHNsNCLDRMlH_x#HCRR:HCM0oRCs:j=R;C
Lo
HMRHRlMH_#x:CR=CR8b;0E
HRRV#R5HRxC<CR8b20ERC0EMR
RRHRlMH_#x:CR=HR#x
C;RMRC8VRH;R
RskC0slMRH#M_H;xC
CRRMo8RCC0_M88_CEb0;0
N0LsHkR0CoCCMsFN0sC_sb0FsR#:R0MsHo-;
-0N0skHL0oCRCsMCNs0F_bsCFRs0FMVRFI_s_COEO:	RRONsECH0Os0kC#RHRMVkOM_HHs05Ns88_osC2-;
-CRLoRHMLODF	NRsllRHblDCCNM00MHFRo#HM#ND
MVkOF0HM0R#soHM.P#D5:NRRs#0H2MoR0sCkRsM#_08DHFoOC_POs0FR
H#PHNsNCLDRP#DR#:R0D8_FOoH_OPC05FsNH'EoNE-'IDFRI8FMR0Fj
2;PHNsNCLDR:HRR0HMCsoC;C
Lo
HMRFRVsRRHHjMRRR0F#'DPEEHoRFDFbR
RRVRHR55NNH'EoHE-2RR='24'RC0EMR
SRP#D5RH2:'=R4
';S#CDCR
SRP#D5RH2:'=Rj
';S8CMR;HV
CRRMD8RF;Fb
sRRCs0kMDR#PC;
M#8R0MsHoD.#PV;
k0MOHRFM#.DP#H0sMNo5R#:R0D8_FOoH_OPC02FsR0sCkRsM#H0sMHoR#N
PsLHND#CRR#:R0MsHo'5NEEHo-DN'F4I+RI8FMR0F4
2;PHNsNCLDR:HRR0HMCsoC;C
Lo
HMRFRVsRRHHNMR'IDFRR0FNH'EoDERF
FbRRRRH5VRN25HR'=R4R'20MEC
RSR#-5HNF'DI2+4RR:=';4'
DSC#SC
R5R#H'-ND+FI4:2R=jR''S;
CRM8H
V;RMRC8FRDF
b;RCRs0MksR
#;CRM8#.DP#H0sM
o;Ns00H0LkCORG_Fbsb:#RRs#0H;Mo
O--F0M#NRM0#NsPDRR:#_08DHFoOC_POs0F58IH04E-RI8FMR0Fj:2R=0R#soHM.P#D50s#_08NN
2;-L-RCMoHRFLDOs	RNHlRlCbDl0CMNF0HMHR#oDMN#k
VMHO0FoMRCO0_EOFHCH_I850EI0H8ERR:HCM0o2CsR0sCkRsMHCM0oRCsHP#
NNsHLRDCPRND:MRH0CCos=R:R
j;PHNsNCLDRP8HdR.,84HPn8,RH,PURP8Hc8,RH,P.RP8H4RR:HCM0o;Cs
oLCHRM
RP8Hd:.R=IR5HE80-/42d
n;RHR8PR4n:5=RI0H8E2-4/;4U
8RRHRPU:5=RI0H8E2-4/
g;RHR8P:cR=IR5HE80-/42cR;
RP8H.=R:RH5I8-0E4.2/;R
R84HPRR:=58IH04E-2R;
RRHV5P8H4RR>j02RE
CMRRRRPRND:P=RN+DRR
4;RMRC8VRH;R
RH5VR8.HPRj>R2ER0CRM
RPRRN:DR=NRPDRR+4R;
R8CMR;HV
HRRV8R5HRPc>2RjRC0EMR
RRNRPD=R:RDPNR4+R;R
RCRM8H
V;RVRHRH58P>URRRj20MEC
RRRRDPNRR:=PRND+;R4
CRRMH8RVR;
RRHV5P8H4>nRRRj20MEC
RRRRDPNRR:=PRND+;R4
CRRMH8RV-;
-HRRV8R5H.PdRj>R2ER0C-M
-RRRRDPNRR:=PRND+;R4
R--R8CMR;HV
HRRVPR5N>DRRR.20MEC
RRRR0sCkRsM5*.R*NRPDRR+.*R*RN5PDRR-d;22
CRRD
#CRRRRskC0s5MR.*R*RDPN2R;
R8CMR;HV
8CMR0oC_FOEH_OCI0H8EV;
k0MOHRFMo_C0OHEFO8C_CEb05b8C0:ERR0HMCsoC2CRs0MksR0HMCsoCR
H#PHNsNCLDRO8_EOFHCC_8bR0E:MRH0CCos=R:R
j;LHCoMR
RH5VR80CbERR>U.4g2ER0CRM
R8RR_FOEH_OC80CbE=R:Rd4nU
c;RDRC#RHV5b8C0<ER=4RUgN.RM88RCEb0Rc>RjRgn2ER0CRM
R8RR_FOEH_OC80CbE=R:RgU4.R;
R#CDH5VR80CbE=R<RgcjnMRN8CR8bR0E>jR.cRU20MEC
RRRRO8_EOFHCC_8bR0E:c=Rj;gn
CRRDV#HRC58bR0E<.=RjRcUNRM880CbERR>4cj.R02RE
CMRRRR8E_OFCHO_b8C0:ER=jR.c
U;RDRC#RHV5b8C0<ER=jR4.NcRM88RCEb0R6>R4R.20MEC
RRRRO8_EOFHCC_8bR0E:4=Rj;.c
CRRDV#HRC58bR0E<6=R4R.20MEC
RRRRO8_EOFHCC_8bR0E:6=R4
.;RMRC8VRH;R
RskC0s8MR_FOEH_OC80CbEC;
Mo8RCO0_EOFHCC_8b;0E
MVkOF0HMCRo0H_I8_0El_F8UE5OFCHO_RI8:MRH0CCoss2RCs0kMMRH0CCos#RH
sPNHDNLCHRI8_0El_F8URR:HCM0o;Cs
oLCHRM
RRHV5FOEH_OCI>8RRRU20MEC
RRRR8IH0lE_FU8_RR:=OHEFOIC_8RR-5FOEH_OCIl8RFU8R2R;
R#CDCR
RRHRI8_0El_F8U=R:RFOEH_OCI
8;RMRC8VRH;R
RskC0sIMRHE80_8lF_
U;CRM8o_C0I0H8EF_l8;_U
F
OMN#0MI0R_FOEH_OCI0H8ERR:HCM0oRCs:o=RCO0_EOFHCH_I850EI0H8E
2;O#FM00NMROI_EOFHCC_8bR0E:MRH0CCos=R:Rd4nUoc/CI0_HE80_8lF_IU5_FOEH_OCI0H8E
2;O#FM00NMRO8_EOFHCC_8bR0E:MRH0CCos=R:R0oC_FOEH_OC80CbEC58b20E;F
OMN#0M80R_FOEH_OCI0H8ERR:HCM0oRCs:5=R4Undc_/8OHEFO8C_CEb02RR+5n54d/Uc8E_OFCHO_b8C0RE2/2RU;V

k0MOHRFMo_C0M_klODCD#85IRH:RMo0CCOs;EOFHC8_IRH:RMo0CCRs2skC0sHMRMo0CCHsR#N
PsLHNDMCRkOl_C#DDRH:RMo0CC
s;LHCoMR
RM_klODCD#=R:R85I-/42OHEFOIC_8RR+4R;
R0sCkRsMM_klODCD#C;
Mo8RCM0_kOl_C#DD;V

k0MOHRFMo_C0#CHx5OIMRH:RMo0CCRs;8RMO:MRH0CCoss2RCs0kMMRH0CCos#RH
oLCHRM
RCRs0MksROIMR8*RM
O;CRM8o_C0#CHx;V

k0MOHRFMo_C0LDFF8_58#CHxRH:RMo0CCRs;IH_#x:CRR0HMCsoC;_R8O:IRR0HMCsoC;_RIO:IRR0HMCsoC2CRs0MksR0HMCsoCR
H#LHCoMV
HR_58#CHxRR<=IH_#xRC20MEC
sRRCs0kM_R8O
I;CCD#
sRRCs0kM_RIO
I;CRM8H
V;CRM8o_C0LDFF8
;
O#FM00NMRFOEH_OCI0H8ERR:HCM0oRCs:o=RCL0_F8FD50oC_x#HCC5o0k_MlC_OD5D#I0H8E8,R_FOEH_OCI0H8Eo2,CM0_kOl_C#DD5b8C0RE,8E_OFCHO_b8C02E2,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRoRRC#0_H5xCo_C0M_klODCD#H5I8,0EROI_EOFHCH_I820E,0oC_lMk_DOCD8#5CEb0,_RIOHEFO8C_CEb02
2,SSSSSSSSSRSS8E_OFCHO_8IH0RE,IE_OFCHO_8IH0;E2
MOF#M0N0HRI8_0EM_klODCD#RR:HCM0oRCs:o=RCL0_F8FD50oC_x#HCC5o0k_MlC_OD5D#I0H8E8,R_FOEH_OCI0H8Eo2,CM0_kOl_C#DD5b8C0RE,8E_OFCHO_b8C02E2,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRCRo0H_#xoC5CM0_kOl_C#DD58IH0RE,IE_OFCHO_8IH0,E2o_C0M_klODCD#C58b,0EROI_EOFHCC_8b20E2S,
SSSSSSSSSRSRRIR5HE80-/428E_OFCHO_8IH0RE,58IH04E-2_/IOHEFOIC_HE802RR+4O;
F0M#NRM080CbEk_MlC_ODRD#:MRH0CCos=R:R0oC_FLFDo85C#0_H5xCo_C0M_klODCD#H5I8,0ERO8_EOFHCH_I820E,0oC_lMk_DOCD8#5CEb0,_R8OHEFO8C_CEb02
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRoRRC#0_H5xCo_C0M_klODCD#H5I8,0EROI_EOFHCH_I820E,0oC_lMk_DOCD8#5CEb0,_RIOHEFO8C_CEb02
2,SSSSSSSSSRSRRC58b-0E482/_FOEH_OC80CbE5,R80CbE2-4/OI_EOFHCC_8b20ER4+R;
SRO#FM00NMRsxCFRR:#_08DHFoOC_POs0F5FOEH_OCI0H8EH*I8_0EM_klODCD#H-I8-0E4FR8IFM0RRj2:5=RFC0Es=#R>jR''
2;O#FM00NMRP#sN#D_D:PRR8#0_oDFHPO_CFO0sE5OFCHO_8IH0IE*HE80_lMk_DOCD4#-RI8FMR0Fj:2R=CRxs&FRRs#0H.Mo#5DPs_#08NN02O;
F0M#NRM0#NsPDRR:#H0sMOo5EOFHCH_I8*0EI0H8Ek_MlC_ODRD#8MFI04FR2=R:RP#D.s#0H5Mo#NsPDD_#P
2;-L-RCMoHRFLDOs	RNHlRlCbDl0CMNF0HMHR#oDMN#$
0bFCRkL0_k_#40C$bRRH#NNss$8R5CEb0_lMk_DOCD4#-RI8FMR0FjI,RHE80_lMk_DOCD4#-RI8FMR0FjF2RV0R#8F_Do;HO
o#HMRNDF_k0L4k#RF:RkL0_k_#40C$b;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFVsF_8k50RHkMb0FR0RH0s-N#002C#
b0$CkRF0k_L#0._$RbCHN#Rs$sNRC58b_0EM_klODCD#R-48MFI0jFR,*R.I0H8Ek_MlC_OD+D#4FR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNR0Fk_#Lk.RR:F_k0L.k#_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFR8s_FRk05bHMk00RFsR0H0-#N#0C2$
0bFCRkL0_k_#c0C$bRRH#NNss$8R5CEb0_lMk_DOCD4#-RI8FMR0Fjc,R*8IH0ME_kOl_C#DD+8dRF0IMF2RjRRFV#_08DHFoO#;
HNoMDkRF0k_L#:cRR0Fk_#Lkc$_0bRC;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RV_Rs80FkRM5HbRk000FRs#H-0CN0#02
$RbCF_k0LUk#_b0$C#RHRsNsN5$R80CbEk_MlC_OD-D#4FR8IFM0RRj,UH*I8_0EM_klODCD#R+(8MFI0jFR2VRFR8#0_oDFH
O;#MHoNFDRkL0_kR#U:kRF0k_L#0U_$;bCRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$FsVR_k8F0HR5M0bkRR0F0-sH#00NC
#20C$bRsbNH_0$LUk#_b0$C#RHRsNsN5$R80CbEk_MlC_OD-D#4FR8IFM0RRj,I0H8Ek_MlC_OD-D#4FR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNRsbNH_0$LUk#Rb:RN0sH$k_L#0U_$;bCRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFR8s_FRk05bHMk00RFsR0H0-#N#0C2$
0bFCRkL0_kn#4_b0$C#RHRsNsN5$R80CbEk_MlC_OD-D#4FR8IFM0RRj,4In*HE80_lMk_DOCD4#+6FR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNR0Fk_#Lk4:nRR0Fk_#Lk40n_$;bCRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$FsVR_k8F0HR5M0bkRR0F0-sH#00NC
#20C$bRsbNH_0$L4k#n$_0bHCR#sRNsRN$5b8C0ME_kOl_C#DD-84RF0IMF,RjRI.*HE80_lMk_DOCD4#+RI8FMR0FjF2RV0R#8F_Do;HO
o#HMRNDbHNs0L$_kn#4Rb:RN0sH$k_L#_4n0C$b;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFVsF_8k50RHkMb0FR0RH0s-N#002C#
b0$CkRF0k_L#_d.0C$bRRH#NNss$8R5CEb0_lMk_DOCD4#-RI8FMR0Fjd,R.H*I8_0EM_klODCD#4+dRI8FMR0FjF2RV0R#8F_Do;HO
o#HMRNDF_k0Ldk#.RR:F_k0Ldk#.$_0bRC;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RV_Rs80FkRM5HbRk000FRs#H-0CN0#02
$RbCbHNs0L$_k.#d_b0$C#RHRsNsN5$R80CbEk_MlC_OD-D#4FR8IFM0RRj,cH*I8_0EM_klODCD#R+d8MFI0jFR2VRFR8#0_oDFH
O;#MHoNbDRN0sH$k_L#Rd.:NRbs$H0_#Lkd0._$;bCRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$FsVR_k8F0HR5M0bkRR0F0-sH#00NC
#2#MHoNFDRkC0_MRR:#_08DHFoOC_POs0F5b8C0ME_kOl_C#DD-84RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RNCML#DCRsVFRH0s-N#00
C##MHoNIDRsC0_MRR:#_08DHFoOC_POs0F5b8C0ME_kOl_C#DD-84RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RHIs0CCRMDNLCV#RFCsRNROEsRFIF)VRqOvRC#DD
o#HMRNDHsM_C:oRR8#0_oDFHPO_CFO0sH5I8+0Ed86RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-k-R#RC80sFRC#oH0RCs7RQh
o#HMRNDF_k0sRCo:0R#8F_Do_HOP0COFIs5HE80+Rd68MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-k-R#RC80sFRC#oH0RCs7amz
o#HMRNDF_k0s4CoR#:R0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-#RkC08RFEROFCF#R0LCIMCCRh7QR8NMR0FkbRk0FAVRD	FORv)q
o#HMRNDs_N8sRCo:0R#8F_Do_HOP0COFNs58I8sHE80-84RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-k-R#RC80sFRC#oH0RCs)7q7)H
#oDMNR8IN_osCR#:R0D8_FOoH_OPC05FsNs88I0H8ER-48MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--k8#CRR0FsHCo#s0CR7Wq7#)
HNoMDFRDIN_s8R8s:0R#8F_Do_HOP0COF4s5dFR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-NRs8R8sL#H0RbHMk00RFqR)vCRODRD#5LcRHR0#skCJH8sC2H
#oDMNRIDF_8IN8:sRR8#0_oDFHPO_CFO0sd54RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-R8IN8LsRHR0#HkMb0FR0Rv)qRDOCD5#RcHRL0s#RCHJks2C8
o#HMRND)7q7)l_0bRR:#_08DHFoOC_POs0F58N8s8IH04E-RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RCk#8FR0RbbHCMDHCqR)7
7)#MHoNWDRq)77_b0lR#:R0D8_FOoH_OPC05FsNs88I0H8ER-48MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--k8#CRR0FbCHbDCHMR7Wq7#)
HNoMDQR7hl_0bRR:#_08DHFoOC_POs0F58IH04E-RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-k-R#RC80bFRHDbCHRMC7
Qh#MHoNWDR l_0bRR:#_08DHFoOR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--k8#CRR0FbCHbDCHMR
W -C-RML8RD	FORlsNRbHlDCClM00NHRFM#MHoN
D#-L-RCMoHRD#CCRO0sRNlHDlbCMlC0HN0F#MRHNoMDV#
k0MOHRFMo_C0M_kln8c5CEb0:MRH0CCoss2RCs0kMMRH0CCos#RH
sPNHDNLCNRPDRR:HCM0oRCs:j=R;C
Lo
HMRNRPD=R:Rb8C0nE/cR;
RRHV5C58bR0ElRF8nRc2>URc2ER0CRM
RPRRN:DR=NRPDRR+4R;
R8CMR;HV
sRRCs0kMNRPDC;
Mo8RCM0_knl_cV;
k0MOHRFMo_C0D0CVFsPC_5d.80CbERR:HCM0o2CsR0sCkRsMHCM0oRCsHL#
CMoH
sRRCs0kMC58bR0ElRF8n;c2
8CMR0oC_VDC0CFPs._d;k
VMHO0FoMRCD0_CFV0P5Cs80CbERR:HCM0o;CsRGlNRH:RMo0CCRs2skC0sHMRMo0CCHsR#N
PsLHNDPCRN:DRR0HMCsoCRR:=jL;
CMoH
HRRV8R5CEb0Rl-RN>GR=2RjRC0EMR
RRNRPD=R:Rb8C0-ERRGlN;R
RCCD#
RRRRDPNRR:=80CbER;
R8CMR;HV
sRRCs0kMN5PD
2;CRM8o_C0D0CVFsPC;k
VMHO0FoMRCM0_kdl_.C58bR0E:MRH0CCoss2RCs0kMMRH0CCos#RH
sPNHDNLCNRPDRR:HCM0oRCs:j=R;C
Lo
HMRVRHRC58bR0E<c=RUMRN8CR8bR0E>nR42ER0CRM
RRRRPRND:4=R;R
RCRM8H
V;RCRs0MksRDPN;M
C8CRo0k_Ml._d;k
VMHO0FoMRCM0_k4l_nC58bR0E:MRH0CCoss2RCs0kMMRH0CCos#RH
sPNHDNLCNRPDRR:HCM0oRCs:j=R;C
Lo
HMRVRHRC58bR0E<4=RnMRN8CR8bR0E>2RjRC0EMR
RRPRRN:DR=;R4
CRRMH8RVR;
R0sCkRsMP;ND
8CMR0oC_lMk_;4n
MOF#M0N0kRMlC_ODnD_cRR:HCM0oRCs:o=RCM0_knl_cC58b20E;F
OMN#0MD0RCFV0P_Csd:.RR0HMCsoCRR:=o_C0D0CVFsPC_5d.80CbE
2;O#FM00NMRlMk_DOCD._dRH:RMo0CC:sR=CRo0k_Ml._d5VDC0CFPs._d2O;
F0M#NRM0D0CVFsPC_R4n:MRH0CCos=R:R0oC_VDC0CFPsC5DVP0FCds_.d,R.
2;O#FM00NMRlMk_DOCDn_4RH:RMo0CC:sR=CRo0k_Mln_45VDC0CFPsn_42
;
0C$bR0Fk_#Lk_b0$Cc_n##RHRsNsN5$RM_klODCD_Rnc8MFI0jFR,HRI8-0E4FR8IFM0RRj2F#VR0D8_FOoH;$
0bFCRkL0_k0#_$_bCdR.#HN#Rs$sNRk5MlC_ODdD_.FR8IFM0RRj,I0H8ER-48MFI0jFR2VRFR8#0_oDFH
O;0C$bR0Fk_#Lk_b0$Cn_4##RHRsNsN5$RM_klODCD_R4n8MFI0jFR,HRI8-0E4FR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNR0Fk_#Lk_#ncRF:RkL0_k0#_$_bCn;c#RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$F8VRFRk05bHMk00RFsR0H0-#N#0C2H
#oDMNR0Fk_#Lk_#d.RF:RkL0_k0#_$_bCd;.#RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$F8VRFRk05bHMk00RFsR0H0-#N#0C2H
#oDMNR0Fk_#Lk_#4nRF:RkL0_k0#_$_bC4;n#RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$F8VRFRk05bHMk00RFsR0H0-#N#0C2H
#oDMNR0Fk__CM#RR:#_08DHFoOC_POs0F5lMk_DOCDc_nRI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-C-RMDNLCV#RF0sRs#H-0CN0#H
#oDMNR0Fk__CMd:.RR8#0_oDFH
O;#MHoNFDRkC0_Mn_4R#:R0D8_FOoH;H
#oDMNR0Is__CM#RR:#_08DHFoOC_POs0F5lMk_DOCDc_nRI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-I-RsCH0RNCML#DCRsVFROCNEFRsIVRFRv)qRDOCD##
HNoMDsRI0M_C_Rd.:0R#8F_Do;HO
o#HMRNDI_s0C4M_nRR:#_08DHFoO#;
HNoMDMRH_osC_:#RR8#0_oDFHPO_CFO0sH5I8-0E4FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-#RkC08RFCRso0H#C7sRQ
hR#MHoNFDRks0_C#o_R#:R0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-k-R#RC80sFRC#oH0RCs7amz
o#HMRNDs_N8s_Co#RR:#_08DHFoOC_POs0F58N8s8IH04E-RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RCk#8FR0RosCHC#0s7Rq7#)
HNoMDNRI8C_soR_#:0R#8F_Do_HOP0COFNs58I8sHE80-84RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-k-R#RC80sFRC#oH0RCsq)77
o#HMRNDD_FIs8N8sR_#:0R#8F_Do_HOP0COF6s5RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-R8N8sHRL0H#RM0bkRR0F)RqvODCD#cR5R0LH#CRsJskHC
82#MHoNDDRFII_Ns88_:#RR8#0_oDFHPO_CFO0sR568MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--Ns88R0LH#MRHbRk00)FRqOvRC#DDRR5cL#H0RJsCkCHs8-2
-MRC8CR#D0CORlsNRbHlDCClM00NHRFM#MHoN
D#Ns00H0LkC3R\s_NlF#VVCR0\:0R#soHM;L

CMoH
RRRRR--QNVR8I8sHE80RO<REOFHCH_I8R0ENH##o'MRj0'RFMRkk8#CR0LH#R
RRjRzRRR:H5VRNs88I0H8ERR=4o2RCsMCN
0CSRRRRIDF_8sN8<sR=jR"jjjjjjjjjjjj"RR&s_N8s5Coj
2;SRRRRIDF_8IN8<sR=jR"jjjjjjjjjjjj"RR&I_N8s5Coj
2;S8CMRMoCC0sNCjRz;R
RR4RzRRR:H5VRNs88I0H8ERR=.o2RCsMCN
0CSFSDIN_s8R8s<"=Rjjjjjjjjjjjj"RR&s_N8s5Co4FR8IFM0R;j2
RSRRFRDIN_I8R8s<"=Rjjjjjjjjjjjj"RR&I_N8s5Co4FR8IFM0R;j2
MSC8CRoMNCs0zCR4R;
RzRR.:RRRRHV58N8s8IH0=ERRRd2oCCMsCN0
DSSFsI_Ns88RR<="jjjjjjjjjjj"RR&s_N8s5Co.FR8IFM0R;j2
RSRRFRDIN_I8R8s<"=Rjjjjjjjjj"jjRI&RNs8_C.o5RI8FMR0Fj
2;S8CMRMoCC0sNC.Rz;R
RRdRzRRR:H5VRNs88I0H8ERR=co2RCsMCN
0CSFSDIN_s8R8s<"=RjjjjjjjjjRj"&NRs8C_soR5d8MFI0jFR2S;
RRRRD_FII8N8s=R<Rj"jjjjjjjjj"RR&I_N8s5CodFR8IFM0R;j2
MSC8CRoMNCs0zCRdR;
RzRRc:RRRRHV58N8s8IH0=ERRR62oCCMsCN0
RSRRFRDIN_s8R8s<"=Rjjjjjjjjj&"RR8sN_osC58cRF0IMF2Rj;R
SRDRRFII_Ns88RR<="jjjjjjjjRj"&NRI8C_soR5c8MFI0jFR2S;
CRM8oCCMsCN0R;zc
RRRRRz6RH:RVNR58I8sHE80Rn=R2CRoMNCs0SC
RRRRD_FIs8N8s=R<Rj"jjjjjjRj"&NRs8C_soR568MFI0jFR2S;
SIDF_8IN8<sR=jR"jjjjj"jjRI&RNs8_C6o5RI8FMR0Fj
2;S8CMRMoCC0sNC6Rz;R
RRnRzRRR:H5VRNs88I0H8ERR=(o2RCsMCN
0CSRRRRIDF_8sN8<sR=jR"jjjjjRj"&NRs8C_soR5n8MFI0jFR2S;
SIDF_8IN8<sR=jR"jjjjjRj"&NRI8C_soR5n8MFI0jFR2S;
CRM8oCCMsCN0R;zn
RRRRRz(RH:RVNR58I8sHE80RU=R2CRoMNCs0SC
RRRRD_FIs8N8s=R<Rj"jjjjj"RR&s_N8s5Co(FR8IFM0R;j2
DSSFII_Ns88RR<="jjjj"jjRI&RNs8_C(o5RI8FMR0Fj
2;S8CMRMoCC0sNC(Rz;R
RRURzRRR:H5VRNs88I0H8ERR=go2RCsMCN
0CSRRRRIDF_8sN8<sR=jR"jjjj"RR&s_N8s5CoUFR8IFM0R;j2
DSSFII_Ns88RR<="jjjjRj"&NRI8C_soR5U8MFI0jFR2S;
CRM8oCCMsCN0R;zU
RRRRRzgRH:RVNR58I8sHE80R4=Rjo2RCsMCN
0CSRRRRIDF_8sN8<sR=jR"j"jjRs&RNs8_Cgo5RI8FMR0Fj
2;SFSDIN_I8R8s<"=Rjjjj"RR&I_N8s5CogFR8IFM0R;j2
MSC8CRoMNCs0zCRgR;
RzRR4RjR:VRHR85N8HsI8R0E=4R42CRoMNCs0SC
RRRRD_FIs8N8s=R<Rj"jj&"RR8sN_osC5R4j8MFI0jFR2S;
SIDF_8IN8<sR=jR"jRj"&NRI8C_soj54RI8FMR0Fj
2;S8CMRMoCC0sNC4RzjR;
RzRR4R4R:VRHR85N8HsI8R0E=.R42CRoMNCs0SC
RRRRD_FIs8N8s=R<Rj"j"RR&s_N8s5Co484RF0IMF2Rj;S
SD_FII8N8s=R<Rj"j"RR&I_N8s5Co484RF0IMF2Rj;C
SMo8RCsMCNR0Cz;44
RRRR.z4RRR:H5VRNs88I0H8ERR=4Rd2oCCMsCN0
RSRRFRDIN_s8R8s<'=Rj&'RR8sN_osC5R4.8MFI0jFR2S;
SIDF_8IN8<sR=jR''RR&I_N8s5Co48.RF0IMF2Rj;C
SMo8RCsMCNR0Cz;4.
RRRRdz4RRR:H5VRNs88I0H8ERR>4Rd2oCCMsCN0
RSRRFRDIN_s8R8s<s=RNs8_C4o5dFR8IFM0R;j2
RSRRFRDIN_I8R8s<I=RNs8_C4o5dFR8IFM0R;j2
MSC8CRoMNCs0zCR4
d;
RRRRR--Q5VR8_HMs2CoRosCHC#0sQR7h#RkHRMoB
piRRRRzR4cRH:RV8R5HsM_CRo2oCCMsCN0
RRRRRRRRFbsO#C#Rp5Bi7,RQRh2LHCoMR
RRRRRRRRRRVRHRp5BiRR='R4'NRM8B'piCMPC002RE
CMRRRRRRRRRRRRRRRRHsM_C<oR="R5jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"RR&72Qh;R
RRRRRRRRRRMRC8VRH;R
RRRRRRMRC8sRbF#OC#S;
CRM8oCCMsCN0Rcz4;R
RR4Rz6:RRRRHV50MFRM8H_osC2CRoMNCs0RC
RRRRRRRRRHRRMC_so=R<Rj5"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jjR7&RQ;h2
MSC8CRoMNCs0zCR4
6;
RRRRz7ma=R<R0Fk_osC58IH04E-RI8FMR0Fj
2;
RRRRR--Q5VRs8N8sC_sos2RC#oH0RCs)7q7)#RkHRMomiBp
RRRRnz4s:RRRRHV58sN8ss_CRo2oCCMsCN0
R--RRRRRbRRsCFO#5#RmiBp,qR)727)RoLCH-M
-RRRRRRRRRRRRRHV5pmBiRR='R4'NRM8miBp'CCPMR020MEC
R--RRRRRRRRRRRRRsRRNs8_C<oR=qR)757)Ns88I0H8ER-48MFI0jFR2-;
-RRRRRRRRRRRR8CMR;HV
R--RRRRRCRRMb8RsCFO#
#;-C-SMo8RCsMCNR0Czs4n;-
-RRRRzs4(RH:RVMR5Fs0RNs88_osC2CRoMNCs0RC
RRRRRRRRRsRRNs8_C<oR=qR)7;7)
MSC8CRoMNCs0zCR4;ns
-
S-VRQRN5I8_8ss2CoRosCHC#0sqRW7R7)kM#Ho_RWmiBp
RRRRnz4I:RRRRHV58IN8ss_CRo2oCCMsCN0
RRRRRRRRFbsO#C#Rp5BiW,Rq)772CRLo
HMRRRRRRRRRRRRH5VRBRpi=4R''MRN8pRBiP'CC2M0RC0EMR
RRRRRRRRRRRRRRNRI8C_so=R<R7Wq7N)58I8sHE80-84RF0IMF2Rj;R
RRRRRRRRRRMRC8VRH;R
RRRRRRMRC8sRbF#OC#S;
CRM8oCCMsCN0Rnz4IR;
RzRR4R(I:VRHRF5M0NRI8_8ss2CoRMoCC0sNCR
RRRRRRRRRRNRI8C_so=R<R7Wq7
);S8CMRMoCC0sNC4Rz(
I;
RRRRR--tCCMsCN0RC0ERv)qRDOCDN#RM#8RCODC0FRDoRHOVRFs)Aqv41n_44_1
4SzURR:H5VROHEFOIC_HE80R4=R2CRoMNCs0RC
RSRRzR4g:FRVsRRHH5MR80CbEk_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0SC
-Q-RVNR58I8sHE80R4>RcM2RCRC80OFRs0CNCsRIHR0CCLMNDNCRMF8Rkk0b0MRCNCLDRD#CCRO0DHFoOR
RRRRRRzRS.:jRRRHV58N8s8IH0>ERR24cRMoCC0sNC-
S-HRVGFRVsNROD4DRd(UU,CR#D0CORRFV0#sH0CN0R0MFRHLCMsoRC#oH0CCs8S
SSkSF0M_C5RH2<'=R4I'RERCM58sN_osC58N8s8IH04E-RI8FMR0F4Rc2=2RHR#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=WI RERCM58IN_osC58N8s8IH04E-RI8FMR0F4Rc2=2RHR#CDCjR''R;
RRRRRSRRCRM8oCCMsCN0Rjz.;-
S-VRQR85N8HsI8R0E<4=RcM2RFsRIHR0CCLMNDFCRskRF00bkRNCMLRDC#CCDOD0RFOoHRCMC8
C8RRSRRzRS.:4RRRHV58N8s8IH0<ER=cR42CRoMNCs0SC
SFSSkC0_M25HRR<=';4'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RW;R
RRRRRRCRSMo8RCsMCNR0Cz;.4
-S-RMtCC0sNCER0CqR)vCRODRD#NRM80-sH#00NCR#
RRRRRSRRzR..:FRVsRR[H5MRI0H8Ek_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0SC
S0SN0LsHkR0CGbO_s#FbRRFVAv)q_d4nU4cX7RR:DCNLD#RHR)"WQ_a v m7_)q= _q7w1Q)a1,R)peq_"A=R#&RsDPN54[+2RR&"W,R) Qa_7vm =_A"RR&Ils_F;8C
RRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVAv)q_d4nU4cX7RR:DCNLD#RHR7"Aa&"RR0HMCsoC'NHloIC5HE802RR&"R7"&MRH0CCosl'HN5oCHn*4d2UcR"&RW&"RR0HMCsoC'NHlo[C52RR&"R "&MRH0CCosl'HN5oCo_C0C_M880CbEH55R4+R2n*4d,UcRb8C02E2R"&RX&"RR0HMCsoC'NHlo[C5+;42
SSSLHCoMR
RRRRRRRRRRARS)_qv4Undc7X4R):Rq4vAn4_1_
14SRRRRRRRRRRRRsbF0NRlb7R5Qjq52>R=R_HMs5Co[R2,q)77q>R=RIDF_8IN84s5dFR8IFM0R,j2RA7QRR=>",j"R7q7)=AR>FRDIN_s858s48dRF0IMF2Rj,S
SShS q>R=R W_h1,R1R)q='>RjR',WR q=I>RsC0_M25H,pRBi=qR>pRBi ,Rh=AR>hR ,1R1)=AR>1R)aW,R =AR>jR''B,RpRiA=m>RB,pi
SSSRRRR7Rmq=F>Rb,CMRA7m5Rj2=F>RkL0_k5#4H2,[2
;
RRRRRRRRRRRRRRRRF_k0s5Co[<2R=kRF0k_L#H45,R[2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRMSC8CRoMNCs0zCR.
.;RRRRRMSC8CRoMNCs0zCR4
g;RRRRCRM8oCCMsCN0RUz4;RRRRR
RRRRR
RRRRR--tCCMsCN0RC0ERv)qRDOCDN#RM#8RCODC0FRDoRHOVRFs)Aqv41n_.._1
.SzdRR:H5VROHEFOIC_HE80R.=R2CRoMNCs0RC
RSRRzR.c:FRVsRRHH5MR80CbEk_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0SC
-Q-RVNR58I8sHE80R4>RdM2RCRC80OFRs0CNCsRIHR0CCLMNDNCRMF8Rkk0b0MRCNCLDRD#CCRO0DHFoOR
RRRRRRzRS.:6RRRHV58N8s8IH0>ERR24dRMoCC0sNC-
S-HRVGFRVsNROD4DRd(UU,CR#D0CORRFV0#sH0CN0R0MFRHLCMsoRC#oH0CCs8R
RRRRRRRRRRRRRRkRF0M_C5RH2<'=R4I'RERCM58sN_osC58N8s8IH04E-RI8FMR0F4Rd2=2RHR#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=WI RERCM58IN_osC58N8s8IH04E-RI8FMR0F4Rd2=2RHR#CDCjR''R;
RRRRRSRRCRM8oCCMsCN0R6z.;-
S-VRQR85N8HsI8R0E<4=RdM2RFsRIHR0CCLMNDFCRskRF00bkRNCMLRDC#CCDOD0RFOoHRCMC8
C8RRSRRzRS.:nRRRHV58N8s8IH0<ER=dR42CRoMNCs0SC
RRRRRRRRRRRRF_k0CHM52=R<R''4;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R R;
RRRRRSRRCRM8oCCMsCN0Rnz.;-
S-CRtMNCs00CRE)CRqOvRC#DDR8NMRH0s-N#00
C#RRRRRRRRS(z.RV:RF[sRRRHM58IH0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CSNSS0H0sLCk0R_GObbsF#VRFRqA)v4_Ug..X7RR:DCNLD#RHR)"WQ_a v m7_)q= _q7w1Q)a1,R)peq_"A=R#&RsDPN5[.*+8.RF0IMF*R.[2+4R"&R,)RWQ_a v m7_"A=RI&RsF_l8
C;RRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FAVR)_qvU.4gXR.7:NRDLRCDH"#RA"7aRH&RMo0CCHs'lCNo58IH0RE2&7R""RR&HCM0o'CsHolNC*5HU.4g2RR&"RW"&MRH0CCosl'HN5oC[2*.R"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05R5H+2R4*gU4.8,RCEb02&2RR""XRH&RMo0CCHs'lCNo5+5[4.2*2S;
SCSLo
HMRRRRRRRRRRRRSqA)v4_Ug..X7RR:)Aqv41n_.._1
RSRRRRRRRRRRFRbsl0RN5bR7RQq=H>RMC_so*5.[R+48MFI0.FR*,[2R7q7)=qR>FRDIN_I858s48.RF0IMF2Rj,QR7A>R=Rj"j"q,R7A7)RR=>D_FIs8N8s.54RI8FMR0Fj
2,SRSSR RRh=qR>_RW Rh,1q1)RR=>',j'RqW RR=>I_s0CHM52B,RpRiq=B>RpRi, RhA= >Rh1,R1R)A=)>R1Ra,WR A='>RjR',BApiRR=>miBp,S
SSRRRRq7mRR=>FMbC,mR7A254RR=>F_k0L.k#5.H,*4[+27,RmjA52>R=R0Fk_#Lk.,5HR[.*2
2;RRRRRRRRRRRRRRRRF_k0s5Co.2*[RR<=F_k0L.k#5.H,*R[2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5[.*+R42<F=RkL0_k5#.H*,.[2+4RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRCRSMo8RCsMCNR0Cz;.(
RRRRCRSMo8RCsMCNR0Cz;.c
RRRR8CMRMoCC0sNC.RzdR;R
R
SR-RR-CRtMNCs00CRE)CRqOvRC#DDR8NMRD#CCRO0DHFoOFRVsqR)vnA4__1c1Sc
zR.U:VRHRE5OFCHO_8IH0=ERRRc2oCCMsCN0
RRRR.SzgRR:VRFsHMRHRC58b_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
-S-RRQV58N8s8IH0>ERR24.RCMC8FR0RCOsNR0CI0sHCMRCNCLDR8NMR0FkbRk0CLMND#CRCODC0FRDo
HORRRRRRRRSjzdRH:RVNR58I8sHE80R4>R.o2RCsMCN
0CSR--VRHGVRFsODNDRU4dUR(,#CCDOF0RVsR0HN#00MCRFL0RCoHMRosCHC#0s
C8RRRRRRRRRRRRRRRRF_k0CHM52=R<R''4RCIEMsR5Ns8_CNo58I8sHE80-84RF0IMF.R42RR=HC2RDR#C';j'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RWRCIEMIR5Ns8_CNo58I8sHE80-84RF0IMF.R42RR=HC2RDR#C';j'
RRRRRRRRMSC8CRoMNCs0zCRd
j;SR--Q5VRNs88I0H8E=R<R24.RRMFI0sHCMRCNCLDRRFsFbk0kC0RMDNLCCR#D0CORoDFHMORCCC88S
RRRRRS4zdRH:RVNR58I8sHE80RR<=4R.2oCCMsCN0
SSSS0Fk_5CMH<2R=4R''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=W
 ;RRRRRRRRS8CMRMoCC0sNCdRz4S;
-t-RCsMCNR0C0REC)RqvODCD#MRN8sR0H0-#N#0C
RRRRRRRRdSz.RR:VRFs[MRHRH5I8_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
SSSNs00H0LkCORG_FbsbF#RV)RAqcv_jXgnc:7RRLDNCHDR#WR") Qa_7vm =_q)7 q_)wQ1Ra,1q)ep=_A"RR&#NsPD*5c[R+c8MFI0cFR*4[+2RR&"W,R) Qa_7vm =_A"RR&Ils_F;8C
RRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVAv)q_gcjn7XcRD:RNDLCRRH#"aA7"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloHC5*gcjn&2RR""WRH&RMo0CCHs'lCNo5c[*2RR&"R "&MRH0CCosl'HN5oCo_C0C_M880CbEH55R4+R2j*cgRn,80CbER22&XR""RR&HCM0o'CsHolNC[55+*42c
2;SLSSCMoH
RRRRRRRRRRRR)SAqcv_jXgnc:7RRv)qA_4n11c_cR
SRRRRRRRRRbRRFRs0lRNb5q7QRR=>HsM_Cco5*d[+RI8FMR0Fc2*[,7Rq7R)q=D>RFII_Ns885R448MFI0jFR27,RQ=AR>jR"j"jj,7Rq7R)A=D>RFsI_Ns885R448MFI0jFR2S,
S SSh=qR>_RW Rh,1q1)RR=>',j'RqW RR=>I_s0CHM52B,RpRiq=B>RpRi, RhA= >Rh1,R1R)A=)>R1Ra,WR A='>RjR',BApiRR=>miBp,S
SSmS7q>R=RCFbM7,RmdA52>R=R0Fk_#Lkc,5HR[c*+,d2RA7m5R.2=F>RkL0_k5#cH*,c[2+.,SR
S7SSm4A52>R=R0Fk_#Lkc,5Hc+*[4R2,75mAj=2R>kRF0k_L#Hc5,*Rc[;22
RRRRRRRRRRRRRRRR0Fk_osC5[c*2=R<R0Fk_#Lkc,5Hc2*[RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so*5c[2+4RR<=F_k0Lck#5cH,*4[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cco5*.[+2=R<R0Fk_#Lkc,5Hc+*[.I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Coc+*[d<2R=kRF0k_L#Hc5,[c*+Rd2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
R
RRRRRRCRSMo8RCsMCNR0Cz;d.
RRRRCRSMo8RCsMCNR0Cz;.g
RRRR8CMRMoCC0sNC.RzU
;
SRRRRR--tCCMsCN0RC0ERv)qRDOCDN#RM#8RCODC0FRDoRHOVRFs)Aqv41n_gg_1
dSzdRR:H5VROHEFOIC_HE80Rg=R2CRoMNCs0RC
RSRRzRdc:FRVsRRHH5MR80CbEk_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0SC
-Q-RVNR58I8sHE80R4>R4M2RCRC80OFRs0CNCsRIHR0CCLMNDNCRMF8Rkk0b0MRCNCLDRD#CCRO0DHFoOR
RRRRRRzRSd:6RRRHV58N8s8IH0>ERR244RMoCC0sNC-
S-HRVGFRVsNROD4DRd(UU,CR#D0CORRFV0#sH0CN0R0MFRHLCMsoRC#oH0CCs8R
RRRRRRRRRRRRRRkRF0M_C5RH2<'=R4I'RERCM58sN_osC58N8s8IH04E-RI8FMR0F4R42=2RHR#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=WI RERCM58IN_osC58N8s8IH04E-RI8FMR0F4R42=2RHR#CDCjR''R;
RRRRRSRRCRM8oCCMsCN0R6zd;-
S-VRQR85N8HsI8R0E<4=R4M2RFsRIHR0CCLMNDFCRskRF00bkRNCMLRDC#CCDOD0RFOoHRCMC8
C8RRSRRzRSd:nRRRHV58N8s8IH0<ER=4R42CRoMNCs0SC
RRRRRRRRRRRRF_k0CHM52=R<R''4;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R R;
RRRRRSRRCRM8oCCMsCN0Rnzd;-
S-CRtMNCs00CRE)CRqOvRC#DDR8NMRH0s-N#00
C#RRRRRRRRS(zdRV:RF[sRRRHM58IH0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CSNSS0H0sLCk0R_GObbsF#VRFRqA)vj_.cUUX7RR:DCNLD#RHR)"WQ_a v m7_)q= _q7w1Q)a1,R)peq_"A=R#&RsDPN5[g*+8gRF0IMF*Rg[2+4R"&R,)RWQ_a v m7_"A=RI&RsF_l8
C;RRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FAVR)_qv.UjcXRU7:NRDLRCDH"#RA"7aRH&RMo0CCHs'lCNo58IH0RE2&7R""RR&HCM0o'CsHolNC*5H.Ujc2RR&"RW"&MRH0CCosl'HN5oC[2*gR"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05R5H+2R4*c.jU8,RCEb02&2RR""XRH&RMo0CCHs'lCNo5+5[4g2*2S;
SCSLo
HMRRRRRRRRRRRRSqA)vj_.cUUX7RR:)Aqv41n_gg_1
RRRRRRRRRRRRRRRRbRRFRs0lRNb5q7QRR=>HsM_Cgo5*([+RI8FMR0Fg2*[,7Rq7R)q=D>RFII_Ns885R4j8MFI0jFR27,RQ=AR>jR"jjjjj"jj,7Rq7R)A=D>RFsI_Ns885R4j8MFI0jFR2S,
S SSh=qR>_RW Rh,1q1)RR=>',j'RqW RR=>I_s0CHM52B,RpRiq=B>RpRi, RhA= >Rh1,R1R)A=)>R1Ra,WR A='>RjR',BApiRR=>miBp,SR
S7SSm=qR>bRFCRM,75mA(=2R>kRF0k_L#HU5,[U*+,(2RA7m5Rn2=F>RkL0_k5#UH*,U[2+n,SR
S7SSm6A52>R=R0Fk_#LkU,5HU+*[6R2,75mAc=2R>kRF0k_L#HU5,[U*+,c2RA7m5Rd2=F>RkL0_k5#UH*,U[2+d,SR
S7SSm.A52>R=R0Fk_#LkU,5HU+*[.R2,75mA4=2R>kRF0k_L#HU5,[U*+,42RA7m5Rj2=F>RkL0_k5#UH*,U[R2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRu7Qq25jRR=>HsM_Cgo5*U[+27,RQRuA=">Rj
",RRRRRRRRRRRRRRRRRRRRRRRRRRRR7qmuRR=>FMbC,mR7ujA52>R=RsbNH_0$LUk#5[H,2
2;RRRRRRRRRRRRRRRRF_k0s5Cog2*[RR<=F_k0LUk#5UH,*R[2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5[g*+R42<F=RkL0_k5#UH*,U[2+4RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so*5g[2+.RR<=F_k0LUk#5UH,*.[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cgo5*d[+2=R<R0Fk_#LkU,5HU+*[dI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cog+*[c<2R=kRF0k_L#HU5,[U*+Rc2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5[g*+R62<F=RkL0_k5#UH*,U[2+6RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so*5g[2+nRR<=F_k0LUk#5UH,*n[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cgo5*([+2=R<R0Fk_#LkU,5HU+*[(I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cog+*[U<2R=NRbs$H0_#LkU,5H[I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRS8CMRMoCC0sNCdRz(R;
RRRRS8CMRMoCC0sNCdRzcR;
RCRRMo8RCsMCNR0Cz;dd
R
SR-RR-CRtMNCs00CRE)CRqOvRC#DDR8NMRD#CCRO0DHFoOFRVsqR)vnA4_U14_U14
dSzURR:H5VROHEFOIC_HE80R4=RUo2RCsMCN
0CRRRRSgzdRV:RFHsRRRHM5b8C0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CSR--Q5VRNs88I0H8ERR>4Rj2M8CCRR0FONsC0ICRsCH0RNCMLRDCNRM8Fbk0kC0RMDNLCCR#D0CORoDFHRO
RRRRRSRRzRcj:VRHR85N8HsI8R0E>jR42CRoMNCs0SC
-V-RHVGRFOsRNRDD4UdU(#,RCODC0VRFRH0s#00NCFRM0CRLHRMosHCo#s0CCR8
RRRRRRRRRRRRRFRRkC0_M25HRR<='R4'IMECRN5s8C_so85N8HsI8-0E4FR8IFM0R24jRH=R2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0CHM52=R<RRW IMECRN5I8C_so85N8HsI8-0E4FR8IFM0R24jRH=R2DRC#'CRj
';RRRRRRRRS8CMRMoCC0sNCcRzjS;
-Q-RVNR58I8sHE80RR<=4Rj2MIFRsCH0RNCMLRDCFFsRkk0b0MRCNCLDRD#CCRO0DHFoOCRMC88C
RRSRSRRzRc4:VRHR85N8HsI8R0E<4=Rjo2RCsMCN
0CSRRRRRRRRRRRR0Fk_5CMH<2R=4R''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=W
 ;RRRRRRRRS8CMRMoCC0sNCcRz4S;
-t-RCsMCNR0C0REC)RqvODCD#MRN8sR0H0-#N#0C
RRRRRRRRcSz.RR:VRFs[MRHRH5I8_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
SSSNs00H0LkCORG_FbsbF#RV)RAq4v_jX.c4Rn7:NRDLRCDH"#RWa)Q m_v7q _=q) 7Q_w),1aRe1)qAp_=&"RRP#sN4D5U+*[48URF0IMFUR4*4[+2RR&"W,R) Qa_7vm =_A"RR&Ils_F;8C
RRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVAv)q_.4jcnX47RR:DCNLD#RHR7"Aa&"RR0HMCsoC'NHloIC5HE802RR&"R7"&MRH0CCosl'HN5oCHj*4.Rc2&WR""RR&HCM0o'CsHolNC*5[4RU2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50E5+HRR*424cj.,CR8b20E2RR&"RX"&MRH0CCosl'HN5oC54[+2U*42S;
SCSLo
HMRRRRRRRRRRRRSqA)vj_4.4cXn:7RRv)qA_4n1_4U1
4URRRRRRRRRRRRRRRRRFRbsl0RN5bR7RQq=H>RMC_soU54*4[+6FR8IFM0R*4U[R2,q)77q>R=RIDF_8IN8gs5RI8FMR0FjR2,7RQA=">Rjjjjjjjjjjjjjjjj"q,R7A7)RR=>D_FIs8N8sR5g8MFI0jFR2S,
S SSh=qR>_RW Rh,1q1)RR=>',j'RqW RR=>I_s0CHM52B,RpRiq=B>RpRi, RhA= >Rh1,R1R)A=)>R1Ra,WR A='>RjR',BApiRR=>miBp,SR
S7SSm=qR>bRFCRM,75mA4R62=F>RkL0_kn#454H,n+*[4,62RA7m524cRR=>F_k0L4k#n,5H4[n*+24c,SR
S7SSm4A5d=2R>kRF0k_L#54nHn,4*4[+dR2,75mA4R.2=F>RkL0_kn#454H,n+*[4,.2RA7m5244RR=>F_k0L4k#n,5H4[n*+244,SR
S7SSm4A5j=2R>kRF0k_L#54nHn,4*4[+jR2,75mAg=2R>kRF0k_L#54nHn,4*g[+27,RmUA52>R=R0Fk_#Lk4Hn5,*4n[2+U,SR
S7SSm(A52>R=R0Fk_#Lk4Hn5,*4n[2+(,mR7A25nRR=>F_k0L4k#n,5H4[n*+,n2RA7m5R62=F>RkL0_kn#454H,n+*[6R2,
SSSSA7m5Rc2=F>RkL0_kn#454H,n+*[cR2,75mAd=2R>kRF0k_L#54nHn,4*d[+27,Rm.A52>R=R0Fk_#Lk4Hn5,*4n[2+.,SR
S7SSm4A52>R=R0Fk_#Lk4Hn5,*4n[2+4,mR7A25jRR=>F_k0L4k#n,5H4[n*2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRR7qQuRR=>HsM_C4o5U+*[48(RF0IMFUR4*4[+nR2,7AQuRR=>""jj,mR7u=qR>bRFC
M,RRRRRRRRRRRRRRRRRRRRRRRRRRRR7Amu5R42=b>RN0sH$k_L#54nH*,.[2+4,mR7ujA52>R=RsbNH_0$L4k#n,5H.2*[2R;
RRRRRRRRRRRRRFRRks0_C4o5U2*[RR<=F_k0L4k#n,5H4[n*2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[4<2R=kRF0k_L#54nHn,4*4[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[.<2R=kRF0k_L#54nHn,4*.[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[d<2R=kRF0k_L#54nHn,4*d[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[c<2R=kRF0k_L#54nHn,4*c[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[6<2R=kRF0k_L#54nHn,4*6[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[n<2R=kRF0k_L#54nHn,4*n[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[(<2R=kRF0k_L#54nHn,4*([+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[U<2R=kRF0k_L#54nHn,4*U[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[g<2R=kRF0k_L#54nHn,4*g[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[4Rj2<F=RkL0_kn#454H,n+*[4Rj2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[4+42=R<R0Fk_#Lk4Hn5,*4n[4+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[4R.2<F=RkL0_kn#454H,n+*[4R.2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[d+42=R<R0Fk_#Lk4Hn5,*4n[d+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[4Rc2<F=RkL0_kn#454H,n+*[4Rc2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[6+42=R<R0Fk_#Lk4Hn5,*4n[6+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[4Rn2<b=RN0sH$k_L#54nH*,.[I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+24(RR<=bHNs0L$_kn#45.H,*4[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''
;
RRRRRRRRS8CMRMoCC0sNCcRz.R;
RRRRS8CMRMoCC0sNCdRzgR;
RCRRMo8RCsMCNR0Cz;dU
R
SR-RR-CRtMNCs00CRE)CRqOvRC#DDR8NMRD#CCRO0DHFoOFRVsqR)vnA4_n1d_n1d
dSzU:NRRRHV5FOEH_OCI0H8ERR=dRn2oCCMsCN0
RSRRdRzg:NRRsVFRHHRM8R5CEb0_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNC-
S-VRQR85N8HsI8R0E>2RgRCMC8FR0RCOsNR0CI0sHCMRCNCLDR8NMR0FkbRk0CLMND#CRCODC0FRDo
HOSzSScRjN:VRHR85N8HsI8R0E>2RgRMoCC0sNC-
S-HRVGFRVsNROD4DRd(UU,CR#D0CORRFV0#sH0CN0R0MFRHLCMsoRC#oH0CCs8S
SSkSF0M_C5RH2<'=R4I'RERCM58sN_osC58N8s8IH04E-RI8FMR0Fg=2RRRH2CCD#R''j;S
SSsSI0M_C5RH2<W=R ERIC5MRI_N8s5CoNs88I0H8ER-48MFI0gFR2RR=HC2RDR#C';j'
SSSCRM8oCCMsCN0RjzcNS;
-Q-RVNR58I8sHE80RR<=gM2RFsRIHR0CCLMNDFCRskRF00bkRNCMLRDC#CCDOD0RFOoHRCMC8
C8SzSScR4N:VRHR85N8HsI8R0E<g=R2CRoMNCs0SC
SFSSkC0_M25HRR<=';4'
SSSS0Is_5CMH<2R= RW;S
SS8CMRMoCC0sNCcRz4
N;SR--tCCMsCN0RC0ERv)qRDOCDN#RM08Rs#H-0CN0#S
SS.zcNRR:VRFs[MRHRH5I8_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
SSSNs00H0LkCORG_FbsbF#RV)RAq6v_4d.X.:7RRLDNCHDR#WR") Qa_7vm =_q)7 q_)wQ1Ra,1q)ep=_A"RR&#NsPDn5d*d[+nFR8IFM0R*dn[2+4R"&R,)RWQ_a v m7_"A=RI&RsF_l8
C;RRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FAVR)_qv6X4.dR.7:NRDLRCDH"#RA"7aRH&RMo0CCHs'lCNo58IH0RE2&7R""RR&HCM0o'CsHolNC*5H624.R"&RW&"RR0HMCsoC'NHlo[C5*2dnR"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05R5H+2R4*.64,CR8b20E2RR&"RX"&MRH0CCosl'HN5oC54[+2n*d2S;
SCSLo
HMSSSSAv)q_.64X7d.R):Rq4vAnd_1nd_1nR
RRRRRRRRRRRRRRRRRRRRRRRRRRFRbsl0RN5bR7RQq=H>RMC_son5d*d[+4FR8IFM0R*dn[R2,q)77q>R=RIDF_8IN8Us5RI8FMR0FjR2,7RQA=">Rjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"q,R7A7)RR=>D_FIs8N8sR5U8MFI0jFR2S,
S SSh=qR>_RW Rh,1q1)RR=>',j'RqW RR=>I_s0CHM52B,RpRiq=B>RpRi, RhA= >Rh1,R1R)A=)>R1Ra,WR A='>RjR',BApiRR=>miBp,S
SSmS7q>R=RCFbM7,RmdA54=2R>kRF0k_L#5d.H.,d*d[+4R2,75mAdRj2=F>RkL0_k.#d5dH,.+*[d,j2
SSSSA7m52.gRR=>F_k0Ldk#.,5Hd[.*+2.g,mR7AU5.2>R=R0Fk_#LkdH.5,*d.[U+.27,Rm.A5(=2R>kRF0k_L#5d.H.,d*.[+(
2,SSSS75mA.Rn2=F>RkL0_k.#d5dH,.+*[.,n2RA7m52.6RR=>F_k0Ldk#.,5Hd[.*+2.6,mR7Ac5.2>R=R0Fk_#LkdH.5,*d.[c+.2S,
S7SSm.A5d=2R>kRF0k_L#5d.H.,d*.[+dR2,75mA.R.2=F>RkL0_k.#d5dH,.+*[.,.2RA7m52.4RR=>F_k0Ldk#.,5Hd[.*+2.4,S
SSmS7Aj5.2>R=R0Fk_#LkdH.5,*d.[j+.27,Rm4A5g=2R>kRF0k_L#5d.H.,d*4[+gR2,75mA4RU2=F>RkL0_k.#d5dH,.+*[4,U2
SSSSA7m524(RR=>F_k0Ldk#.,5Hd[.*+24(,mR7An542>R=R0Fk_#LkdH.5,*d.[n+427,Rm4A56=2R>kRF0k_L#5d.H.,d*4[+6
2,SSSS75mA4Rc2=F>RkL0_k.#d5dH,.+*[4,c2RA7m524dRR=>F_k0Ldk#.,5Hd[.*+24d,mR7A.542>R=R0Fk_#LkdH.5,*d.[.+42S,
S7SSm4A54=2R>kRF0k_L#5d.H.,d*4[+4R2,75mA4Rj2=F>RkL0_k.#d5dH,.+*[4,j2RA7m5Rg2=F>RkL0_k.#d5dH,.+*[g
2,SSSS75mAU=2R>kRF0k_L#5d.H.,d*U[+27,Rm(A52>R=R0Fk_#LkdH.5,*d.[2+(,mR7A25nRR=>F_k0Ldk#.,5Hd[.*+,n2
SSSSA7m5R62=F>RkL0_k.#d5dH,.+*[6R2,75mAc=2R>kRF0k_L#5d.H.,d*c[+27,RmdA52>R=R0Fk_#LkdH.5,*d.[2+d,S
SSmS7A25.RR=>F_k0Ldk#.,5Hd[.*+,.2RA7m5R42=F>RkL0_k.#d5dH,.+*[4R2,75mAj=2R>kRF0k_L#5d.H.,d*,[2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRQRuq=H>RMC_son5d*d[+6FR8IFM0R*dn[.+d27,RQRuA=">Rjjjj"7,RmRuq=F>Rb,CM
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRm5uAd=2R>NRbs$H0_#LkdH.5,[c*+,d2Ru7mA25.RR=>bHNs0L$_k.#d5cH,*.[+2R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRu7mA254RR=>bHNs0L$_k.#d5cH,*4[+27,Rm5uAj=2R>NRbs$H0_#LkdH.5,[c*2
2;RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*R[2<F=RkL0_k.#d5dH,.2*[RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*+R42<F=RkL0_k.#d5dH,.+*[4I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*.[+2=R<R0Fk_#LkdH.5,*d.[2+.RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*+Rd2<F=RkL0_k.#d5dH,.+*[dI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*c[+2=R<R0Fk_#LkdH.5,*d.[2+cRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*+R62<F=RkL0_k.#d5dH,.+*[6I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*n[+2=R<R0Fk_#LkdH.5,*d.[2+nRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*+R(2<F=RkL0_k.#d5dH,.+*[(I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*U[+2=R<R0Fk_#LkdH.5,*d.[2+URCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*+Rg2<F=RkL0_k.#d5dH,.+*[gI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*4[+j<2R=kRF0k_L#5d.H.,d*4[+jI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*4[+4<2R=kRF0k_L#5d.H.,d*4[+4I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*4[+.<2R=kRF0k_L#5d.H.,d*4[+.I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*4[+d<2R=kRF0k_L#5d.H.,d*4[+dI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*4[+c<2R=kRF0k_L#5d.H.,d*4[+cI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*4[+6<2R=kRF0k_L#5d.H.,d*4[+6I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*4[+n<2R=kRF0k_L#5d.H.,d*4[+nI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*4[+(<2R=kRF0k_L#5d.H.,d*4[+(I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*4[+U<2R=kRF0k_L#5d.H.,d*4[+UI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*4[+g<2R=kRF0k_L#5d.H.,d*4[+gI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*.[+j<2R=kRF0k_L#5d.H.,d*.[+jI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*.[+4<2R=kRF0k_L#5d.H.,d*.[+4I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*.[+.<2R=kRF0k_L#5d.H.,d*.[+.I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*.[+d<2R=kRF0k_L#5d.H.,d*.[+dI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*.[+c<2R=kRF0k_L#5d.H.,d*.[+cI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*.[+6<2R=kRF0k_L#5d.H.,d*.[+6I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*.[+n<2R=kRF0k_L#5d.H.,d*.[+nI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*.[+(<2R=kRF0k_L#5d.H.,d*.[+(I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*.[+U<2R=kRF0k_L#5d.H.,d*.[+UI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*.[+g<2R=kRF0k_L#5d.H.,d*.[+gI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*d[+j<2R=kRF0k_L#5d.H.,d*d[+jI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*d[+4<2R=kRF0k_L#5d.H.,d*d[+4I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*d[+.<2R=NRbs$H0_#LkdH.5,[c*2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[d+d2=R<RsbNH_0$Ldk#.,5Hc+*[4I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*d[+c<2R=NRbs$H0_#LkdH.5,[c*+R.2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[dR62<b=RN0sH$k_L#5d.H*,c[2+dRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;S

SMSC8CRoMNCs0zCRc;.N
CSSMo8RCsMCNR0CzNdg;C
SMo8RCsMCNR0CzNdU;C

MN8RsHOE00COkRsCMsF_IE_OC;O	
-
-

---p-RNR#0HDlbCMlC0HN0FHMR#CR8VDNk0-
-
ONsECH0Os0kCCR#D0CO_lsNRRFV)hqv_W)_R
H#VOkM0MHFR0oC_8CM_b8C0#E5HRxC:MRH0CCosRR;80CbERR:HCM0o2CsR0sCkRsMHCM0oRCsHP#
NNsHLRDCl_HM#CHxRH:RMo0CC:sR=;Rj
oLCHRM
RMlH_x#HC=R:Rb8C0
E;RVRHRH5#x<CRRb8C0RE20MEC
RRRRMlH_x#HC=R:Rx#HCR;
R8CMR;HV
sRRCs0kMHRlMH_#x
C;CRM8o_C0C_M880CbEO;
F0M#NRM0M_klODCD#RR:HCM0oRCs:5=R5b8C0-ERR/424;n2RRRRRRRRRRRR-y-RRRFV)4qvn7X4RDOCDM#RCCC88$
0bFCRkL0_k0#_$RbCHN#Rs$sNRk5MlC_ODRD#8MFI0jFR,HRI8-0E4FR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNR0Fk_#LkRF:RkL0_k0#_$;bCRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RVFR8k50RHkMb0FR0RH0s-N#002C#
o#HMRNDF_k0C:MRR8#0_oDFHPO_CFO0sk5MlC_ODRD#8MFI0jFR2R;RRRRRR-R-RNCML#DCRsVFRH0s-N#00
C##MHoNIDRsC0_MRR:#_08DHFoOC_POs0F5lMk_DOCD8#RF0IMF2Rj;RRRRRRRRR--I0sHCMRCNCLD#FRVsNRCOsERFFIRVqR)vCROD
D##MHoNHDRMC_soRR:#_08DHFoOC_POs0F58IH04E-RI8FMR0FjR2;RRRRRRRRRR--k8#CRR0FsHCo#s0CRh7QRH
#oDMNR0Fk_osCR#:R0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2R;RRRRRR-RR-#RkC08RFCRso0H#C7sRm
za#MHoNsDRNs8_C:oRR8#0_oDFHPO_CFO0s85N8HsI8-0E4FR8IFM0R;j2RRRRRR--k8#CRR0FsHCo#s0CR7)q7#)
HNoMDNRI8C_soRR:#_08DHFoOC_POs0F58N8s8IH04E-RI8FMR0FjR2;RRRR-k-R#RC80sFRC#oH0RCsW7q7)H
#oDMNRIDF_8sN8:sRR8#0_oDFHPO_CFO0sR5d8MFI0jFR2R;RRRRRRRRRR-RR-NRs8R8sL#H0RbHMk00RFqR)vCRODRD#5LcRHR0#skCJH8sC2H
#oDMNRIDF_8IN8:sRR8#0_oDFHPO_CFO0sR5d8MFI0jFR2R;RRRRRRRRRR-RR-NRI8R8sL#H0RbHMk00RFqR)vCRODRD#5LcRHR0#skCJH8sC20
N0LsHkR0C\N3slV_FV0#C\RR:#H0sM
o;
oLCH
M
RRRR-Q-RV8RN8HsI8R0E<RRcNH##o'MRj0'RFMRkk8#CR0LH#R
RR4RzRRR:H5VRNs88I0H8ERR=4o2RCsMCN
0CRRRRRRRRD_FIs8N8s=R<Rj"jj&"RR8sN_osC5;j2
RRRRRRRRIDF_8IN8<sR=jR"jRj"&NRI8C_so25j;R
RRMRC8CRoMNCs0zCR4R;
RzRR.:RRRRHV58N8s8IH0=ERRR.2oCCMsCN0
RRRRRRRRIDF_8sN8<sR=jR"j&"RR8sN_osC584RF0IMF2Rj;R
RRRRRRFRDIN_I8R8s<"=RjRj"&NRI8C_soR548MFI0jFR2R;
RCRRMo8RCsMCNR0Cz
.;RRRRzRdR:VRHR85N8HsI8R0E=2RdRMoCC0sNCR
RRRRRRFRDIN_s8R8s<'=Rj&'RR8sN_osC58.RF0IMF2Rj;R
RRRRRRFRDIN_I8R8s<'=Rj&'RR8IN_osC58.RF0IMF2Rj;R
RRMRC8CRoMNCs0zCRdR;
RzRRc:RRRRHV58N8s8IH0>ERRRd2oCCMsCN0
RRRRRRRRIDF_8sN8<sR=NRs8C_soR5d8MFI0jFR2R;
RRRRRDRRFII_Ns88RR<=I_N8s5CodFR8IFM0R;j2
RRRR8CMRMoCC0sNCcRz;R

R-RR-VRQRH58MC_sos2RC#oH0RCs7RQhkM#HopRBiR
RR6RzRRR:H5VR8_HMs2CoRMoCC0sNCR
RRRRRRsRbF#OC#BR5pRi,72QhRoLCHRM
RRRRRRRRRHRRVBR5p=iRR''4R8NMRiBp'CCPMR020MEC
RRRRRRRRRRRRRRRR_HMsRCo<7=RQ
h;RRRRRRRRRRRRCRM8H
V;RRRRRRRRCRM8bOsFC;##
RRRR8CMRMoCC0sNC6Rz;R
RRnRzRRR:H5VRMRF08_HMs2CoRMoCC0sNCR
RRRRRRRRRRMRH_osCRR<=7;Qh
RRRR8CMRMoCC0sNCnRz;R

R-RR-VRQRF58ks0_CRo2sHCo#s0CRz7ma#RkHRMomiBp
RRRRRz(RH:RV8R5F_k0s2CoRMoCC0sNCR
RRRRRRsRbF#OC#mR5B,piR0Fk_osC2CRLo
HMRRRRRRRRRRRRH5VRmiBpR'=R4N'RMm8RB'piCMPC002RE
CMRRRRRRRRRRRRRRRR7amzRR<=F_k0s;Co
RRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMRFbsO#C#;R
RRMRC8CRoMNCs0zCR(R;
RzRRU:RRRRHV50MFRk8F0C_soo2RCsMCN
0CRRRRRRRRRRRR7amzRR<=F_k0s;Co
RRRR8CMRMoCC0sNCURz;R

R-RR-VRQRN5s8_8ss2CoRosCHC#0sqR)7R7)kM#HoBRmpRi
RzRRg:RRRRHV58sN8ss_CRo2oCCMsCN0
RRRRRRRRFbsO#C#RB5mpRi,)7q7)L2RCMoH
RRRRRRRRRRRRRHV5pmBiRR='R4'NRM8miBp'CCPMR020MEC
RRRRRRRRRRRRRRRR8sN_osCRR<=)7q7)85N8HsI8-0E4FR8IFM0R;j2
RRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMRFbsO#C#;R
RRMRC8CRoMNCs0zCRgR;
RzRR4:jRRRHV50MFR8sN8ss_CRo2oCCMsCN0
RRRRRRRRRRRR8sN_osCRR<=)7q7)R;
RCRRMo8RCsMCNR0Cz;4j
RRRRRRRRR
RR-R-RRQV58IN8ss_CRo2sHCo#s0CR7Wq7k)R#oHMRiBp
RRRR6z4RRR:H5VRI8N8sC_soo2RCsMCN
0CRRRRRRRRbOsFCR##5iBp,qRW727)RoLCHRM
RRRRRRRRRHRRVBR5p=iRR''4R8NMRiBp'CCPMR020MEC
RRRRRRRRRRRRRRRR8IN_osCRR<=W7q7)85N8HsI8-0E4FR8IFM0R;j2
RRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMRFbsO#C#;R
RRMRC8CRoMNCs0zCR4
6;RRRRzR4n:VRHRF5M0NRI8_8ss2CoRMoCC0sNCR
RRRRRRRRRRNRI8C_so=R<R7Wq7
);RRRRCRM8oCCMsCN0Rnz4;R

R-RR-CRtMNCs00CRE)CRqOvRC#DDR8NMRD#CCRO0DHFoOR
RR4Rz4RR:VRFsHMRHRlMk_DOCD8#RF0IMFRRjoCCMsCN0
RRRRRRRRR--Q5VRNs88I0H8ERR>cM2RCRC80OFRs0CNCsRIHR0CCLMNDNCRMF8Rkk0b0MRCNCLDRD#CCRO0DHFoOR
RRRRRR4Rz.RR:H5VRNs88I0H8ERR>co2RCsMCN
0CRRRRRRRRRRRRRRRRF_k0CHM52=R<R''4RCIEMsR5Ns8_CNo58I8sHE80-84RF0IMF2RcRH=R2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0CHM52=R<RRW IMECRN5I8C_so85N8HsI8-0E4FR8IFM0RRc2=2RHR#CDCjR''R;
RRRRRCRRMo8RCsMCNR0Cz;4.
RRRRRRRRR--Q5VRNs88I0H8E=R<RRc2MIFRsCH0RNCMLRDCFFsRkk0b0MRCNCLDRD#CCRO0DHFoOCRMC88C
RRRRRRRRdz4RH:RVNR58I8sHE80RR<=co2RCsMCN
0CRRRRRRRRRRRRRRRRF_k0CHM52=R<R''4;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R R;
RRRRRRRRRCRRMo8RCsMCNR0Cz;4d
RRRRR--tsMCNR0C0REC)RqvODCD#MRN8sR0H0-#N#0C
RRRRRRRRcz4RV:RF[sRRRHM58IH0-ERRR428MFI0jFRRMoCC0sNCR
RRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqz)vRR:DCNLD#RHR7"1a&"RR0HMCsoC'NHloIC5HE802RR&"R7"&MRH0CCosl'HN5oCHn*42RR&"RW"&MRH0CCosl'HN5oC[&2RR"" RH&RMo0CCHs'lCNo50oC_8CM_b8C05E5H2+4*,4nRb8C02E2R"&RX&"RR0HMCsoC'NHlo[C5+;42
RRRRRRRRRRRRoLCHRM
RRRRRRRRRzRR):qvRv)q44nX7RR
RRRRRRRRRRRRRbRRFRs0lRNb5=7R>MRH_osC5,[2RRqj=D>RFII_Ns885,j2RRq4=D>RFII_Ns885,42RRq.=D>RFII_Ns885,.2
RRRRRRRRRRRRRRRRRRRRRRRRqRRd>R=RIDF_8IN8ds527,Ruj)qRR=>D_FIs8N8s25j,uR7)Rq4=D>RFsI_Ns885,42RR
RRRRRRRRRRRRRRRRRRRRRRRRR7qu).>R=RIDF_8sN8.s527,Rud)qRR=>D_FIs8N8s25d, RWRR=>I_s0CHM52
,RRRRRRRRRRRRRRRRRRRRRRRRRRBRWp=iR>pRBi7,Ru=mR>kRF0k_L#,5H[;22
RRRRRRRRRRRR0Fk_osC5R[2<F=RkL0_kH#5,R[2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRR8CMRMoCC0sNC4RzcR;
RRRRRCRRMo8RCsMCNR0Cz;44
RRRRRRRRRRRRRRRRRRRRRRRRRRRRCR
MN8RsHOE00COkRsC#CCDOs0_N
l;
