--
@ER--B$FbsEHo0OR52gR4g-cRRj.jd$R1MHbDO$H0ROQM
R--fN]C8:CsR#//$DMbH0OH$N/lb0DN.Uj4J4.b/blNb#Cs/0N0/LDH/MoC_OFsN/.Ns_Nls3_IPyE84
Rf-
-


---1-RHDlbCqR)vHRI0#ERCsbCNR0Cq)77 R11VRFss8CNR8NMRHIs0-C
-NRas0oCRp:RkMOC0RR-mq)BR
.q---
-D

HNLssH$RC;CC
Ck#RCHCC03#8F_Do_HO4c4n3DND;#
kCCRHC#C30D8_FOoH_o#HM3C8N;DD
LDHs$NsROFsN
.;kR#CFNsO.s3FOFNOlNb3D
D;CHM00)$Rq)v__HWR#R
RRCRoMHCsO
R5RRRRRRRRVHNlDR$:#H0sM:oR=MR"F"MC;R
RRRRRRHRI8R0E:MRH0CCos=R:RR4;
RRRRRRRR8N8s8IH0:ERR0HMCsoCRR:=cR;RRRRRR-R-RoLHRFCMkRoEVRFs80CbER
RRRRRRCR8bR0E:MRH0CCos=R:RnR4;R
RRRRRRFR8ks0_C:oRRFLFDMCNRR:=V#NDCR;RR-RR-NRE#kRF00bkRosC
RRRRRRRRM8H_osCRL:RFCFDN:MR=NRVD;#CRRRRR-R-R#ENR08NNMRHbRk0s
CoRRRRRRRRs8N8sC_soRR:LDFFCRNM:V=RNCD#;RRRRR--ERN8s8CNR8N8s#C#RosC
RRRRRRRR8IN8ss_C:oRRFLFDMCNRR:=V#NDCRRRR-R-R8ENRHIs0NCR8C8s#s#RCRo
RRRRR2RR;R
RRFRbs50R
RRRRRRRRz7ma:RRR0FkR8#0_oDFHPO_CFO0sH5I8-0E4FR8IFM0R;j2
RRRRRRRR7)q7:)RRRHMR8#0_oDFHPO_CFO0s85N8HsI8-0E4FR8IFM0R;j2
RRRRRRRRh7QR:RRRRHMR8#0_oDFHPO_CFO0sH5I8-0E4FR8IFM0R;j2
RRRRRRRR7Wq7:)RRRHMR8#0_oDFHPO_CFO0s85N8HsI8-0E4FR8IFM0R;j2
RRRRRRRRRW R:RRRRHMR8#0_oDFHRO;RRRRR-R-RHIs0CCRMDNLCFRVsNRslR
RRRRRRpRBiRRR:MRHR0R#8F_Do;HORRRRR-RR-DROFRO	VRFss,NlR8N8s8,RHRM
RRRRRmRRBRpiRH:RM#RR0D8_FOoHRRRRRRRR-F-RbO0RD	FORsVFRk8F0R
RRRRRR;R2
8CMR0CMHR0$)_qv);_W
-
-
R--w#Hs0lRHblDCCNM00MHFR#lk0CRLRDONDRC8NEsOj-
-
ONsECH0Os0kCsRNOREjF)VRq)v__HWR#F
OMN#0MM0RkOl_C#DD_C8CbRR:HCM0oRCs:5=R5b8C0-ERR/424;n2RRRRRRRRRR--yVRFRIsF#VRFRw7B4.nXZCRODRD#M8CCCO8
F0M#NRM0M_klODCD#H_I8:CRR0HMCsoCRR:=5H5I8R0E-2R4/;.2RRRRRRRRR-R-RFyRVFRODMkl#VRFRw7B4.nXZCRODRD#M8CCC#8
HNoMDkRF0M_CRRRR:0R#8F_Do_HOP0COFMs5kOl_C#DD_C8CbFR8IFM0R;j2R-R-RNCML#DCRsVFRH0s-N#00
C##MHoNIDRbCC_MRRRR#:R0D8_FOoH_OPC05FsM_klODCD#C_8C8bRF0IMF2Rj;-RR-sRIHR0CCLMNDRC#VRFsCENORIsFRRFV)RqvODCD#H
#oDMNR_HMsRCoR:RRR8#0_oDFHPO_CFO0sH5I8+0E4FR8IFM0R;j2RRRRRRRRRR--k8#CRR0FsHCo#s0CRh7QRH
#oDMNR0Fk_osCR:RRR8#0_oDFHPO_CFO0sH5I8+0E4FR8IFM0R;j2RRRRRRRRRR--k8#CRR0FsHCo#s0CRz7maH
#oDMNR8sN_osCR:RRR8#0_oDFHPO_CFO0s85N8HsI8-0E4FR8IFM0R;j2RRRRRR--k8#CRR0FsHCo#s0CR7)q7#)
HNoMDNRI8C_soRRR:0R#8F_Do_HOP0COFNs58I8sHE80-84RF0IMF2Rj;RRRR-R-RCk#8FR0RosCHC#0sqRW7
7)#MHoNDDRFsI_Ns88R#:R0D8_FOoH_OPC05FsdFR8IFM0R;j2RRRRRRRRRRRRR-RR-NRs8R8sL#H0RbHMk00RFqR)vCRODRD#5LcRHR0#skCJH8sC2H
#oDMNRIDF_8IN8:sRR8#0_oDFHPO_CFO0sR5d8MFI0jFR2R;RRRRRRRRRRRRRRR--I8N8sHRL0H#RM0bkRR0F)RqvODCD#cR5R0LH#CRsJskHC
82
oLCH
M
RRRR-Q-RV8RN8HsI8R0E<RRcNH##o'MRj0'RFMRkk8#CR0LH#R
RR4RzRRR:H5VRNs88I0H8ERR=4o2RCsMCN
0CRRRRRRRRD_FIs8N8s=R<Rj"jj&"RR8sN_osC5;j2
RRRRRRRRIDF_8IN8<sR=jR"jRj"&NRI8C_so25j;R
RRMRC8CRoMNCs0zCR4R;
RzRR.:RRRRHV58N8s8IH0=ERRR.2oCCMsCN0
RRRRRRRRIDF_8sN8<sR=jR"j&"RR8sN_osC584RF0IMF2Rj;R
RRRRRRFRDIN_I8R8s<"=RjRj"&NRI8C_soR548MFI0jFR2R;
RCRRMo8RCsMCNR0Cz
.;RRRRzRdR:VRHR85N8HsI8R0E=2RdRMoCC0sNCR
RRRRRRFRDIN_s8R8s<'=Rj&'RR8sN_osC58.RF0IMF2Rj;R
RRRRRRFRDIN_I8R8s<'=Rj&'RR8IN_osC58.RF0IMF2Rj;R
RRMRC8CRoMNCs0zCRdR;
RzRRc:RRRRHV58N8s8IH0>ERRRd2oCCMsCN0
RRRRRRRRIDF_8sN8<sR=NRs8C_soR5d8MFI0jFR2R;
RRRRRDRRFII_Ns88RR<=I_N8s5CodFR8IFM0R;j2
RRRR8CMRMoCC0sNCcRz;R

R-RR-VRQRH58MC_sos2RC#oH0RCs7RQhkM#HopRBiR
RR6RzRRR:H5VR8_HMs2CoRMoCC0sNCR
RRRRRRsRbF#OC#BR5pRi,72QhRoLCHRM
RRRRRRRRRHRRVBR5p=iRR''4R8NMRiBp'CCPMR020MEC
RRRRRRRRRRRRRRRR_HMsRCo<5=R""jjR7&RQ;h2
RRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMRFbsO#C#;R
RRMRC8CRoMNCs0zCR6R;
RzRRn:RRRRHV50MFRM8H_osC2CRoMNCs0RC
RRRRRRRRRHRRMC_so=R<Rj5"j&"RRh7Q2R;
RCRRMo8RCsMCNR0Cz
n;
RRRRR--Q5VR80Fk_osC2CRso0H#C7sRmRzakM#HoBRmpRi
RzRR(:RRRRHV5k8F0C_soo2RCsMCN
0CRRRRRRRRbOsFCR##5pmBiF,Rks0_CRo2LHCoMR
RRRRRRRRRRVRHRB5mp=iRR''4R8NMRpmBiP'CC2M0RC0EMR
RRRRRRRRRRRRRRmR7z<aR=kRF0C_soH5I8-0E4FR8IFM0R;j2
RRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMRFbsO#C#;R
RRRRRRMRC8CRoMNCs0zCR(R;
RzRRU:RRRRHV50MFRk8F0C_soo2RCsMCN
0CRRRRRRRRRRRR7amzRR<=F_k0s5CoI0H8ER-48MFI0jFR2R;
RCRRMo8RCsMCNR0Cz
U;
RRRRR--Q5VRs8N8sC_sos2RC#oH0RCs)7q7)#RkHRMoB
piRRRRzRgR:VRHRN5s8_8ss2CoRMoCC0sNCR
RRRRRRsRbF#OC#mR5B,piR7)q7R)2LHCoMR
RRRRRRRRRRVRHRB5mp=iRR''4R8NMRpmBiP'CC2M0RC0EMR
RRRRRRRRRRRRRRNRs8C_so=R<R7)q7N)58I8sHE80-84RF0IMF2Rj;R
RRRRRRRRRRMRC8VRH;R
RRRRRRMRC8sRbF#OC#R;
RCRRMo8RCsMCNR0Cz
g;RRRRzR4j:VRHRF5M0NRs8_8ss2CoRMoCC0sNCR
RRRRRRRRRRNRs8C_so=R<R7)q7
);RRRRCRM8oCCMsCN0Rjz4;R
RRRRRRRR
R-RR-VRQRN5I8_8ss2CoRosCHC#0sqRW7R7)kM#HopRBiR
RR4Rz6:RRRRHV58IN8ss_CRo2oCCMsCN0
RRRRRRRRFbsO#C#Rp5BiW,Rq)772CRLo
HMRRRRRRRRRRRRH5VRBRpi=4R''MRN8pRBiP'CC2M0RC0EMR
RRRRRRRRRRRRRRNRI8C_so=R<R7Wq7N)58I8sHE80-84RF0IMF2Rj;R
RRRRRRRRRRMRC8VRH;R
RRRRRRMRC8sRbF#OC#R;
RCRRMo8RCsMCNR0Cz;46
RRRRnz4RH:RVMR5FI0RNs88_osC2CRoMNCs0RC
RRRRRRRRRIRRNs8_C<oR=qRW7;7)
RRRR8CMRMoCC0sNC4Rzn
;
RRRR-t-RCsMCNR0C0REC)RqvODCD#MRN8CR#D0CORoDFHRO
RzRR4:4RRsVFRHHRMkRMlC_OD_D#8bCCRI8FMR0FjCRoMNCs0RC
R-RR-VRQR85N8HsI8R0E>2RcRCMC8FR0RCOsNR0CI0sHCMRCNCLDR8NMR0FkbRk0CLMND#CRCODC0FRDo
HORRRRRRRRzR4.:VRHR85N8HsI8R0E>2RcRMoCC0sNCR
RRRRRRRRRRRRRRkRF0M_C5RH2<'=RjI'RERCM58sN_osC58N8s8IH04E-RI8FMR0Fc=2RRRH2CCD#R''4;R
RRRRRRRRRRRRRRbRICM_C5RH2<'=R4I'RERCM58IN_osC58N8s8IH04E-RI8FMR0Fc=2RRRH2CCD#R''j;R
RRRRRRRRRRMRC8CRoMNCs0zCR4
.;RRRR-Q-RVNR58I8sHE80RR<=cM2RFsRIHR0CCLMNDFCRskRF00bkRNCMLRDC#CCDOD0RFOoHRCMC8
C8RRRRzR4d:VRHR85N8HsI8R0E<c=R2CRoMNCs0RC
RRRRRRRRRFRRkC0_M25HRR<=';j'
RRRRRRRRRRRRRRRRCIb_5CMH<2R=4R''R;
RRRRRRRRRCRRMo8RCsMCNR0Cz;4d
RRRRR--tsMCNR0C0REC)RqvODCD#HRI00ERs#H-0CN0#R
RRRRRR4RzcRR:VRFs[MRHRlMk_DOCDI#_HR8C8MFI0jFRRMoCC0sNCR
RRRRRRRRRR)RzqRv:74BwnZX.RR
RRRRRRRRRRFRbsl0RN5bRaR)Q=F>RkC0_M25H,QR7j>R=R_HMs5Co5[.*2R2,7RQ4=H>RMC_so.55*+[24R2,
RRRRRRRRRRRRRRRRRRRRRRRRqRR7=jR>FRDIN_I858sjR2,qR74=D>RFII_Ns885,42R.q7RR=>D_FII8N8s25.,7Rqd>R=RIDF_8IN8ds52R,
RRRRRRRRRRRRRRRRRRRRRRRRR7)qj>R=RIDF_8sN8js52),RqR74=D>RFsI_Ns885,42R7)q.>R=RIDF_8sN8.s52),RqR7d=D>RFsI_Ns885,d2
RRRRRRRRRRRRRRRRRRRRRRRRWRR)R h=W>R W,Ru= R>bRICM_C5,H2RRBi=B>RpRi,)j7mRR=>F_k0s5Co5.[*2R2,)47mRR=>F_k0s5Co5.[*22+42R;
RRRRRRRRRCRRMo8RCsMCNR0Cz;4c
RRRRRRRR8CMRMoCC0sNC4Rz4R;
RRRRRRRRRRRRRRRRRRRRRRRRRRRR
8CMRONsECH0Os0kCsRNO;Ej
