-- $Header: //synplicity/maplat2018q2p1/mappers/att/lib/gen_orca5g/cmp_eq.vhd#1 $
@ELDHs$NsRCHCC
;RkR#CHCCC38#0_oDFH4O_43ncN;DD
M
C0$H0R_CJClDCCRM0HR#
RbRRF5s0NRj,LRj,NR4,LR4,N,j4R4Lj,4RN4L,R4R4,DM0HRH:RM0R#8F_Do;HO
RRRRRRRRRRRR0RDF:k0R0FkR8#0_oDFH;O2
8CMR_CJClDCC;M0
N

sHOE00COkRsCCRJMFCVRJD_CCMlC0#RH
HS#oDMNR,04R:0.R8#0_oDFH
O;SO
SFFlbM0CMR7wq7R.
RbRRF5s0
RRRRRRRRqRRj:SSSSHM1_a7ztpmQ
B;RRRRRRRRR4RqSSS:H1MSaz7_pQmtBR;
RRRRRRRRRSAjSH:SMaS17p_zmBtQ;R
RRRRRRRRRAS4S:MSHS71a_mzpt;QB
RRRRRRRRBRRQ:SSSSHM1_a7ztpmQ
B;RRRRRRRRRmRBzSajSF:Sk10Saz7_pQmtBR;
RRRRRRRRRzBmaS4S:kSF0aS17p_zmBtQ;R
RRRRRRRRR1SjS:kSF0aS17p_zmBtQ;R
RRRRRRRRR1S4S:kSF0aS17p_zmBtQ
RRRRRRRR
2;S8CMRlOFbCFMM
0;SN--0H0sLCk0RNLDOL	_FFGRVqRw7R7.:FROlMbFCRM0H0#Rs;kC
oLCHSM
0<4R=NR54MRGFLsR4N2RM58RNGjRMRFsL;j2
.S0RR<=54N4RFGMs4RL4N2RM58RNRj4GsMFR4Lj2R;
RlRRkHG_MR#0:qRw7
7.RRRRRRRRb0FsRblN5R
RRRRRRmRBzRa4=D>R00Fk,R
RRRRRRQRBRR=>DM0H,R
RRRRRRjRqRR=>0
4,RRRRRRRRq=4R>.R0,R
RRRRRRjRARR=>',j'
RRRRRRRRRA4='>Rj2'R;M
C8JRCM
;

H
DLssN$CRHCRC;
Ck#RCHCC03#8F_Do_HO4c4n3DND;C

M00H$vRBuT_ R
H#RRRRoCCMs5HOI0H8ERR:HCM0oRCs:2=n;R
RRFRbsq05:MRHR8#0_oDFHPO_CFO0sH5I8R0E-84RF0IMF2Rj;R
RRRRRRARR:MRHR8#0_oDFHPO_CFO0sH5I8R0E-84RF0IMF2Rj;R
RRRRRR RRTRR:FRk0#_08DHFoO
2;CRM8B_vu 
T;
s
NO0EHCkO0sOCRC_DDDCCPDVRFRuBv_R TH
#
VOkM0MHFRMVkOs_Cs5FsCIJ_HE80RH:RMo0CCRs2skC0s#MR0MsHo#RH
oLCHRM
RRHV5J5C_8IH0>ER=nR42MRN8CR5JH_I8R0E<4=R.2U2RC0EMR
RRCRs0Mks52"";R
RCCD#
RRRR0sCk5sM"sCsF2s";R
RCRM8H
V;CRM8VOkM_sCsF
s;Ns00H0LkCCRoMNCs0_FssFCbs:0RRs#0H;Mo
0N0skHL0oCRCsMCNs0F_bsCFRs0FOVRC_DDDCCPDRR:NEsOHO0C0CksRRH#VOkM_sCsFIs5HE802
;
SMOF#M0N00RHC0sNHRFM:MRH0CCos=R:RH5I820E/
c;SMOF#M0N0CRslMNH8RCs:MRH0CCos=R:RH5I820ER8lFR
c;RRRR#MHoN8DRN_0N0Rlb:0R#8F_Do_HOP0COF5sRI0H8ERR-4FR8IFM0R;j2
R
RRFROlMbFCRM0CCJ_DCClMH0R#R
RRRRRRFRbsN05jL,RjN,R4L,R4N,RjR4,L,j4R4N4,4RL4D,R0:HMRRHM#_08DHFoOR;
RRRRRRRRRRRRRRRRDk0F0RR:FRk0#_08DHFoO
2;RRRRCRM8ObFlFMMC0
;
LHCoMz
SjRR:HRV5I0H8E=R>RRc2oCCMsCN0
CSLo
HMRRRRzRj4:JRC_CCDl0CM
RRRRRRRRRRRRRRRRsbF0NRlbS5
SNSSj>R=Rjq52
,RRRRRRRRRRRRRRRRRL=jR>5RAj
2,SSSSN=4R>5Rq4R2,
RRRRRRRRRRRRRRRRRL4=A>R5,42
SSSS4NjRR=>q25.,RR
RRRRRRRRRRRRRLRRj=4R>5RA.
2,SSSSNR44=q>R5,d2RR
RRRRRRRRRRRRRR4RL4>R=RdA52R,
RRRRRRRRRRRRRDRR0RHM='>R4
',RRRRRRRRRRRRRRRRDk0F0>R=R08NNl_0b25j2S;
CRM8oCCMsCN0;R

RRRRR
RRSRz4:VRH5HRI8R0E=2R4RMoCC0sNCL
SCMoH
 SST=R<Rjq52MRGFAsR5;j2
MSC8CRoMNCs0
C;
RRRRRz.:FRVsHRL0M_H8RCGH4MRRR0F5CH0sHN0F-MRRR42RMoCC0sNCR
RRRRRRCRLo
HMRRRRRRRRRRRRzR.4:JRC_CCDl0CM
RRRRRRRRRRRRRRRRsbF0NRlbS5
SNSSj>R=Rcq5*0LH_8HMC,G2RR
RRRRRRRRRRRRRRjRLRR=>A*5cL_H0HCM8G
2,SSSSN=4R>5RqcH*L0M_H8RCG+2R4,RR
RRRRRRRRRRRRRLRR4>R=RcA5*0LH_8HMC+GRR,42
RRRRRRRRRRRRRRRR4NjRR=>q*5cL_H0HCM8G.R+2
,RRRRRRRRRRRRRRRRRLRj4=A>R5Lc*HH0_MG8CR.+R2S,
SNSS4=4R>5RqcH*L0M_H8RCG+2Rd,RR
RRRRRRRRRRRRRLRR4=4R>5RAcH*L0M_H8RCG+2Rd,R
RRRRRRRRRRRRRR0RDH=MR>NR800N_lLb5HH0_MG8CR4-R2R,
RRRRRRRRRRRRRDRR00FkRR=>8NN0_b0l50LH_8HMC2G2;R
RRRRRRMRC8CRoMNCs0
C;
)Sz4RR:HRV5sNClHCM8sRR=4MRN8HRI8R0E>2RcRMoCC0sNCL
SCMoH
zSS)R44:CRRJD_CCMlC0R
RRRRRRRRRRRRRRFRbsl0RN
b5SSSSN=jR>5RqI0H8ERR-4R2,
RRRRRRRRRRRRRRRRRLj=A>R58IH0-ER4
2,SSSSN=4R>jR''
,RRRRRRRRRRRRRRRRRL=4R>jR''R,
RRRRRRRRRRRRRNRRj=4R>jR''
,RRRRRRRRRRRRRRRRRLRj4='>Rj
',SSSSNR44='>RjR',
RRRRRRRRRRRRRRRR4L4RR=>',j'
RRRRRRRRRRRRRRRRHD0M>R=R08NNl_0b05HC0sNHRFM-2R4,R
RRRRRRRRRRRRRR0RDFRk0= >RT
2;S8CMRMoCC0sNC
;
S.z)RH:RVs5RCHlNMs8CR.=RR8NMR8IH0>ERRRc2oCCMsCN0
CSLo
HMS)Sz.:4RRJRC_CCDl0CM
RRRRRRRRRRRRRRRRsbF0NRlbS5
SNSSj>R=RIq5HE80R4-R2
,RRRRRRRRRRRRRRRRRL=jR>5RAI0H8E4R-2S,
SNSS4>R=RIq5HE80R.-R2
,RRRRRRRRRRRRRRRRRL=4R>5RAI0H8ERR-.
2,RRRRRRRRRRRRRRRRNRj4='>RjR',
RRRRRRRRRRRRRRRR4LjRR=>',j'
SSSS4N4RR=>',j'RR
RRRRRRRRRRRRRR4RL4>R=R''j,R
RRRRRRRRRRRRRR0RDH=MR>NR800N_lHb50NCs0MHFR4-R2R,
RRRRRRRRRRRRRDRR00FkRR=> ;T2
MSC8CRoMNCs0
C;
dSzRH:RVs5RCHlNMs8CRd=RR8NMR8IH0>ERRRc2oCCMsCN0
CSLo
HMSdSz4RR:CCJ_DCClMR0
RRRRRRRRRRRRRbRRFRs0l5Nb
SSSSRNj=q>R58IH0-ERR,42RR
RRRRRRRRRRRRRRjRLRR=>AH5I8R0E-,42
SSSSRN4=q>R58IH0-ERR,.2RR
RRRRRRRRRRRRRR4RLRR=>AH5I8R0E-2R.,R
RRRRRRRRRRRRRRjRN4>R=RIq5HE80Rd-R2
,RRRRRRRRRRRRRRRRRLRj4=A>R58IH0-ERR,d2
SSSS4N4RR=>',j'RR
RRRRRRRRRRRRRR4RL4>R=R''j,R
RRRRRRRRRRRRRR0RDH=MR>NR800N_lHb50NCs0MHFR4-R2R,
RRRRRRRRRRRRRDRR00FkRR=> ;T2
MSC8CRoMNCs0
C;
R
RRRRRRSR
z:cRR5HVsNClHCM8sRR=jMRN8HRI8R0ER4>R2CRoMNCs0SC
LHCoMR
RR RST=R<R08NNl_0b05HC0sNHRFM-2R4;SR
CRM8oCCMsCN0;S


RRRRC

MR8RODCD_PDCC
D;




