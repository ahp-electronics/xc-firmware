--
@ER--B$FbsEHo0OR52gR4g-cRRj.jd$R1MHbDO$H0ROQM
R--fN]C8:CsR#//$DMbH0OH$N/lb0DN.Uj4J4.b/blNb#Cs/DGHH/MGD/HLoCCMs/HOo_CMoCCMs.HO/lsN_3sIPyE84
Rf-
-
DsHLNRs$HCCC;#
kCCRHC#C30D8_FOoH_n44cD3NDk;
#HCRC3CC#_08DHFoOH_#o8MC3DND;H
DLssN$MRkHl#H;#
kCMRkHl#H3FPOlMbFC#M03DND;M
C0$H0RqX)vU4.XR41HR#
RsbF0
R5RRRRRRRRmRRR:kRF00R#8D_kFOoH;R

RRRRRqRRjRRR:MRHR8#0_FkDo;HO
RRRRRRRRRq4RRR:H#MR0k8_DHFoOR;
RRRRRqRR.RRR:MRHR8#0_FkDo;HO
RRRRRRRRRqdRRR:H#MR0k8_DHFoOR;
RRRRRqRRcRRR:MRHR8#0_FkDo;HO
RRRRRRRRRq6RRR:H#MR0k8_DHFoOS;
SRqnRRR:H#MR0k8_DHFoOR;
RRRRR7RRR:RRRRHM#_08koDFH
O;RRRRRRRRWiBpRH:RM0R#8D_kFOoH;R
RRRRRR RWR:RRRRHM#_08koDFHRO
RRRRR;R2
8CMRqX)vU4.X;41
s
NO0EHCkO0s)CRqev_RRFVXv)q4X.U4H1R#H
#oDMNR,0jRR04:0R#8D_kFOoH;H
#oDMNR4IC,CRI.RR:#_08koDFH
O;LHCoMR
RRRRRRRRRRzRX)nqvcRR:)nqvc1X4RR
RRRRRRRRRRRRRRFRbsl0RN5bR7>R=RR7,q=jR>jRq,4RqRR=>qR4,q=.R>.Rq,R
RRRRRRRRRRRRRRRRRRRRRRRRRq=dR>dRq,cRqRR=>qRc,q=6R>6Rq,S
SSSSSR RWRR=>I,C4RpWBi>R=RpWBim,RRR=>0;j2
RRRRRRRRRRRRzX4)nqvcRR:)nqvc1X4RR
RRRRRRRRRRRRRRFRbsl0RN5bR7>R=RR7,q=jR>jRq,4RqRR=>qR4,q=.R>.Rq,R
RRRRRRRRRRRRRRRRRRRRRRRRRq=dR>dRq,cRqRR=>qRc,q=6R>6Rq,S
SSSSSR RWRR=>I,C.RpWBi>R=RpWBim,RRR=>0;42
<mR=jR0RCIEMnRqR'=RjC'RDR#C0
4;IRC4<W=R MRN8FRM0n5q2I;
C<.R= RWR8NMR;qn
M
C8qR)v;_e
D

HNLssH$RC;CC
Ck#RCHCC03#8F_Do_HO4c4n3DND;#
kCCRHC#C30D8_FOoH_o#HM3C8N;DD
LDHs$NsRHkM#;Hl
Ck#RHkM#3HlPlOFbCFMM30#N;DD
0CMHR0$Xv)qn.cX1#RH
bRRFRs05R
RRRRRRjRmR:RRR0FkR8#0_FkDo;HO
RRRRRRRRRm4RRR:FRk0#_08koDFH
O;
RRRRRRRRRqjRRR:H#MR0k8_DHFoOR;
RRRRRqRR4RRR:MRHR8#0_FkDo;HO
RRRRRRRRRq.RRR:H#MR0k8_DHFoOR;
RRRRRqRRdRRR:MRHR8#0_FkDo;HO
RRRRRRRRRqcRRR:H#MR0k8_DHFoOR;
RRRRRqRR6RRR:MRHR8#0_FkDo;HO
RRRRRRRRR7jRRR:H#MR0k8_DHFoOR;
RRRRR7RR4RRR:MRHR8#0_FkDo;HO
RRRRRRRRpWBiRR:H#MR0k8_DHFoOR;
RRRRRWRR RRR:MRHR8#0_FkDo
HORRRRR2RR;M
C8)RXqcvnX;.1
s
NO0EHCkO0s)CRqcvnX_.1eVRFRqX)vXnc.H1R#C
Lo
HMRRRRRRRRRRRRXqz)vRnc:qR)vXnc4
1RRRRRRRRRRRRRRRRRb0FsRblNRR57=7>Rjq,Rj>R=R,qjRRq4=q>R4q,R.>R=R,q.
RRRRRRRRRRRRRRRRRRRRRRRRqRRd>R=R,qdRRqc=q>Rcq,R6>R=R,q6
SSSSRSSRRW =W>R W,RBRpi=W>RB,piR=mR>jRm2R;
RRRRRRRRRXRR4qz)vRnc:qR)vXnc4
1RRRRRRRRRRRRRRRRRb0FsRblNRR57=7>R4q,Rj>R=R,qjRRq4=q>R4q,R.>R=R,q.
RRRRRRRRRRRRRRRRRRRRRRRRqRRd>R=R,qdRRqc=q>Rcq,R6>R=R,q6
SSSSRSSRRW =W>R W,RBRpi=W>RB,piR=mR>4Rm2C;
M)8RqcvnX_.1e
;
DsHLNRs$HCCC;#
kCCRHC#C30D8_FOoH_n44cD3NDk;
#HCRC3CC#_08DHFoOH_#o8MC3DND;H
DLssN$MRkHl#H;#
kCMRkHl#H3FPOlMbFC#M03DND;M
C0$H0RqX)vXd.UH1R#R
Rb0FsRS5
S:mRR0FkR8#0_oDFHPO_CFO0s(5RRI8FMR0Fj
2;RRRRRRRRqRjRRH:RM0R#8D_kFOoH;R
RRRRRR4RqR:RRRRHM#_08koDFH
O;RRRRRRRRqR.RRH:RM0R#8D_kFOoH;R
RRRRRRdRqR:RRRRHM#_08koDFH
O;RRRRRRRRqRcRRH:RM0R#8D_kFOoH;R
RRRRRRRR7R:RRRRHM#_08DHFoOC_POs0FR(5RRI8FMR0Fj
2;RRRRRRRRWiBpRH:RM0R#8D_kFOoH;R
RRRRRR RWR:RRRRHM#_08koDFHRO
RRRRR;R2
8CMRqX)vXd.U
1;
ONsECH0Os0kCqR)vR_eFXVR)dqv.1XUR
H#LHCoMR
RRRRRRRRRRzRX)Rqv:qR)vXd..
1RRRRRRRRRRRRRRRRRb0FsRblNRj57RR=>725j,4R7=7>R5,42RRqj=q>Rjq,R4>R=R,q4RRq.=q>R.R,
RRRRRRRRRRRRRRRRRRRRRRRRRRqd=q>Rdq,Rc>R=R,qcRS
SSSSSR RWRR=>WR ,WiBpRR=>WiBp,jRmRR=>m25j,4RmRR=>m2542R;
RRRRRRRRRXRR4qz)vRR:)dqv.1X.RR
RRRRRRRRRRRRRRFRbsl0RN5bR7=jR>5R7.R2,7>4=Rd752q,Rj>R=R,qjRRq4=q>R4q,R.>R=R,q.
RRRRRRRRRRRRRRRRRRRRRRRRqRRd>R=R,qdRRqc=q>RcS,
SSSSSWRR >R=R,W RpWBi>R=RpWBim,Rj>R=R.m52m,R4>R=Rdm52
2;RRRRRRRRRRRRX).zq:vRRv)qd..X1RR
RRRRRRRRRRRRRbRRFRs0lRNb5R7j=7>R5,c2R=74>5R76R2,q=jR>jRq,4RqRR=>qR4,q=.R>.Rq,R
RRRRRRRRRRRRRRRRRRRRRRRRRq=dR>dRq,cRqRR=>q
c,SSSSSRSRW= R> RW,BRWp=iR>BRWpRi,m=jR>5RmcR2,m=4R>5Rm6;22
RRRRRRRRRRRRzXd)Rqv:qR)vXd..
1RRRRRRRRRRRRRRRRRb0FsRblNRj57RR=>725n,4R7=7>R5,(2RRqj=q>Rjq,R4>R=R,q4RRq.=q>R.R,
RRRRRRRRRRRRRRRRRRRRRRRRRRqd=q>Rdq,Rc>R=R,qc
SSSSRSSRRW =W>R W,RBRpi=W>RB,piRRmj=m>R5,n2RRm4=m>R52(2;M
C8qR)v;_e
LDHs$NsRCHCCk;
#HCRC3CC#_08DHFoO4_4nNc3D
D;kR#CHCCC38#0_oDFH#O_HCoM8D3NDD;
HNLssk$RMHH#lk;
#kCRMHH#lO3PFFlbM0CM#D3ND
;
CHM00X$R)dqv.1XcR
H#RFRbs50R
RRRRjSmRF:Rk#0R0k8_DHFoOR;
RSRRm:4RR0FkR8#0_FkDo;HO
RRRR.SmRF:Rk#0R0k8_DHFoOR;
RSRRm:dRR0FkR8#0_FkDo;HO
R
RRRRRRjRqR:RRRRHM#_08koDFH
O;RRRRRRRRqR4RRH:RM0R#8D_kFOoH;R
RRRRRR.RqR:RRRRHM#_08koDFH
O;RRRRRRRRqRdRRH:RM0R#8D_kFOoH;R
RRRRRRcRqR:RRRRHM#_08koDFH
O;RRRRSR7jRRR:H#MR0k8_DHFoOR;
RSRR7R4RRH:RM0R#8D_kFOoH;R
RR7RS.RRR:MRHR8#0_FkDo;HO
RRRRdS7R:RRRRHM#_08koDFH
O;RRRRRRRRWiBpRH:RM0R#8D_kFOoH;R
RRRRRR RWR:RRRRHM#_08koDFHRO
RRRRR;R2
8CMRqX)vXd.c
1;
ONsECH0Os0kCqR)vR_eFXVR)dqv.1XcR
H#LHCoMR
RRRRRRRRRRzRX)Rqv:qR)vXd..
1RRRRRRRRRRRRRRRRRb0FsRblNRj57RR=>7Rj,7>4=R,74RRqj=q>Rjq,R4>R=R,q4RRq.=q>R.R,
RRRRRRRRRRRRRRRRRRRRRRRRRRqd=q>Rdq,Rc>R=R,qcRS
SSSSSR RWRR=>WR ,WiBpRR=>WiBp,jRmRR=>mRj,m=4R>4Rm2R;
RRRRRRRRRXRR4qz)vRR:)dqv.1X.RR
RRRRRRRRRRRRRRFRbsl0RN5bR7=jR>.R7,4R7=7>Rdq,Rj>R=R,qjRRq4=q>R4q,R.>R=R,q.
RRRRRRRRRRRRRRRRRRRRRRRRqRRd>R=R,qdRRqc=q>RcS,
SSSSSWRR >R=R,W RpWBi>R=RpWBim,Rj>R=R,m.RRm4=m>Rd
2;CRM8)_qveD;
HNLssH$RC;CC
Ck#RCHCC03#8F_Do_HO4c4n3DND;#
kCCRHC#C30D8_FOoH_o#HM3C8N;DD
LDHs$NsRHkM#;Hl
Ck#RHkM#3HlPlOFbCFMM30#N;DD
M
C0$H0RqX)vX4nUH1R#R
Rb0FsRS5
S:mRR0FkR8#0_oDFHPO_CFO0sRR5(FR8IFM0R;j2
RRRRRRRRRqjRRR:H#MR0k8_DHFoOR;
RRRRRqRR4RRR:MRHR8#0_FkDo;HO
RRRRRRRRRq.RRR:H#MR0k8_DHFoOR;
RRRRRqRRdRRR:MRHR8#0_FkDo;HO
RRRRRRRRR7RRRR:H#MR0D8_FOoH_OPC0RFs5RR(8MFI0jFR2R;
RRRRRWRRBRpi:MRHR8#0_FkDo;HO
RRRRRRRRRW RRR:H#MR0k8_DHFoOR
RRRRRR
2;CRM8Xv)q4UnX1
;
NEsOHO0C0CksRv)q_FeRV)RXqnv4XRU1HL#
CMoH
RRRRRRRRRRRR)Xzq:vRRv)q4cnX1RR
RRRRRRRRRRRRRbRRFRs0lRNb5R7j=7>R5,j2R=74>5R74R2,7=.R>5R7.R2,7=dR>5R7dR2,
SSSSRRRRRRRRqRRj>R=R,qjRRq4=q>R4q,R.>R=R,q.RRqd=q>Rd
,RSSSSSRSRW= R> RW,BRWp=iR>BRWpRi,
SSSSRSSRRmj=m>R5,j2RRm4=m>R5,42RRm.=m>R5,.2RRmd=m>R52d2;R
RRRRRRRRRR4RXzv)qR):Rqnv4XRc1
RRRRRRRRRRRRRRRRsbF0NRlb7R5j>R=Rc7527,R4R=>7256,.R7RR=>725n,dR7RR=>725(,SR
SRSSRRRRRRRRRRqj=q>Rjq,R4>R=R,q4RRq.=q>R.q,Rd>R=R,qdRS
SSSSSR RWRR=>WR ,WiBpRR=>WiBp,SR
SSSSSmRRj>R=Rcm52m,R4>R=R6m52m,R.>R=Rnm52m,Rd>R=R(m52
2;CRM8)_qve-;
--
-
R--1bHlD)CRqIvRHR0E#oHMDqCR7 7)1V1RFLsRFR0Es8CNR8NMRHIs0-C
-NRas0oCRX:RHMDHG-
-
LDHs$NsRCHCCk;
#HCRC3CC#_08DHFoO4_4nNc3D
D;kR#CHCCC38#0_oDFH#O_HCoM8D3NDD;
HNLssk$RMHH#lk;
#kCRMHH#lO3PFFlbM0CM#D3NDC;
M00H$qR)vW_)R
H#RRRRoCCMsRHO5R
RRRRRRNRVl$HDR#:R0MsHo=R:RF"MM;C"
RRRRRRRR8IH0:ERR0HMCsoCRR:=U
;RRRRRRRRRNs88I0H8ERR:HCM0oRCs:U=R;RRRRRRRRR--LRHoCkMFoVERF8sRCEb0
RRRRRRRRb8C0:ERR0HMCsoCRR:=.;6n
RRRRRRRRk8F0C_soRR:LDFFCRNM:V=RNCD#;RRRR-R-R#ENR0FkbRk0s
CoRRRRRRRR8_HMsRCo:FRLFNDCM=R:RDVN#RC;RRRRRR--ERN#8NN0RbHMks0RCRo
RRRRRNRR8_8ssRCo:FRLFNDCM=R:RDVN#RCRRRRR-E-RNN8R8C8s#s#RCRo
RRRRR2RR;R
RRFRbs50R
RRRRRRRRz7maF:Rk#0R0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2R;
RRRRR7RRQRhR:MRHR8#0_oDFHPO_CFO0sH5I8-0E4FR8IFM0R;j2
RRRRRRRR7q7)RR:H#MR0D8_FOoH_OPC05FsNs88I0H8ER-48MFI0jFR2R;
RRRRRWRR :RRRRHM#_08DHFoOR;RRRRRRR--I0sHCMRCNCLDRsVFRlsN
RRRRRRRRiBpRH:RM0R#8F_Do;HORRRRR-RR-DROFRO	VRFss,NlR8N8s8,RHRM
RRRRRmRRBRpi:MRHR8#0_oDFHRORRRRRRR--FRb0OODF	FRVsFR8kR0
RRRRR2RR;M
C8MRC0$H0Rv)q_;)W
-
-
R--w#Hs0lRHblDCCNM00MHFR#lk0CRLRDONDRC8NEsOj-
-
ONsECH0Os0kCDRLF_O	sRNlF)VRq)v_W#RH
F
OlMbFCRM0Xv)q4X.U4R1
b0FsRR5
RRRm:kRF00R#8F_Do;HO
RRRq:jRRRHM#_08DHFoOR;
R4RqRH:RM0R#8F_Do;HO
RRRq:.RRRHM#_08DHFoOR;
RdRqRH:RM0R#8F_Do;HO
RRRq:cRRRHM#_08DHFoOR;
R6RqRH:RM0R#8F_Do;HO
RRRq:nRRRHM#_08DHFoOR;
RRR7:MRHR8#0_oDFH
O;RWRRBRpi:MRHR8#0_oDFH
O;RWRR RR:H#MR0D8_FOoH
;R2
8CMRlOFbCFMM
0;
F
OlMbFCRM0Xv)qn.cX1b
RFRs05R
RRRmj:kRF00R#8F_Do;HO
RRRm:4RR0FkR8#0_oDFH
O;RqRRjRR:H#MR0D8_FOoH;R
RRRq4:MRHR8#0_oDFH
O;RqRR.RR:H#MR0D8_FOoH;R
RRRqd:MRHR8#0_oDFH
O;RqRRcRR:H#MR0D8_FOoH;R
RRRq6:MRHR8#0_oDFH
O;R7RRjRR:H#MR0D8_FOoH;R
RRR74:MRHR8#0_oDFH
O;RWRRBRpi:MRHR8#0_oDFH
O;RWRR RR:H#MR0D8_FOoH
;R2
8CMRlOFbCFMM
0;
lOFbCFMMX0R)dqv.1Xc
FRbs50R
RRRm:jRR0FkR8#0_oDFH
O;RmRR4RR:FRk0#_08DHFoOR;
R.RmRF:Rk#0R0D8_FOoH;R
RRRmd:kRF00R#8F_Do;HO
RRRq:jRRRHM#_08DHFoOR;
R4RqRH:RM0R#8F_Do;HO
RRRq:.RRRHM#_08DHFoOR;
RdRqRH:RM0R#8F_Do;HO
RRRq:cRRRHM#_08DHFoOR;
RjR7RH:RM0R#8F_Do;HO
RRR7:4RRRHM#_08DHFoOR;
R.R7RH:RM0R#8F_Do;HO
RRR7:dRRRHM#_08DHFoOR;
RBRWp:iRRRHM#_08DHFoOR;
R RWRH:RM0R#8F_Do
HOR
2;CRM8ObFlFMMC0O;
FFlbM0CMRqX)vXd.U
1
RsbF0
R5RmRRRF:Rk#0R0D8_FOoH_OPC05Fs(FR8IFM0R;j2
RRRq:jRRRHM#_08DHFoOR;
R4RqRH:RM0R#8F_Do;HO
RRRq:.RRRHM#_08DHFoOR;
RdRqRH:RM0R#8F_Do;HO
RRRq:cRRRHM#_08DHFoOR;
RRR7:MRHR8#0_oDFHPO_CFO0sR5(8MFI0jFR2R;
RBRWp:iRRRHM#_08DHFoOR;
R RWRH:RM0R#8F_Do
HOR
2;CRM8ObFlFMMC0
;
ObFlFMMC0)RXqnv4X
U1RsbF0
R5RmRRRF:Rk#0R0D8_FOoH_OPC05Fs(FR8IFM0R;j2
RRRq:jRRRHM#_08DHFoOR;
R4RqRH:RM0R#8F_Do;HO
RRRq:.RRRHM#_08DHFoOR;
RdRqRH:RM0R#8F_Do;HO
RRR7RR:H#MR0D8_FOoH_OPC05Fs(FR8IFM0R;j2
RRRWiBpRH:RM0R#8F_Do;HO
RRRW: RRRHM#_08DHFoO2
R;M
C8FROlMbFC;M0
k
VMHO0FVMRk_MOH0MH5:LRRFLFDMCN2CRs0MksRs#0HRMoHL#
CMoH
HRRVLR52ER0CRM
RsRRCs0kM"5"2R;
R#CDCR
RRCRs0Mks5F"BkRD8MRF0HDlbCMlC0DRAFRO	)3qvRRQ#0RECs8CNR8N8s#C#RosCHC#0sRC8kM#HoER0CNR#lOCRD	FORRN#0REC)?qv"
2;RMRC8VRH;M
C8kRVMHO_M;H0
MVkOF0HMCRo0M_C8C_8b50E#CHxRH:RMo0CC;sRRb8C0:ERR0HMCsoC2CRs0MksR0HMCsoCR
H#PHNsNCLDRMlH_x#HCRR:HCM0oRCs:j=R;C
Lo
HMRHRlMH_#x:CR=CR8b;0E
HRRV#R5HRxC<CR8b20ERC0EMR
RRHRlMH_#x:CR=HR#x
C;RMRC8VRH;R
RskC0slMRH#M_H;xC
8CMR0oC_8CM_b8C0
E;Ns00H0LkCCRoMNCs0_FssFCbs:0RRs#0H;Mo
0N0skHL0oCRCsMCNs0F_bsCFRs0FLVRD	FO_lsNRN:RsHOE00COkRsCHV#Rk_MOH0MH58N8sC_so
2;-L-RCMoHRFLDOs	RNHlRlCbDl0CMNF0HMHR#oDMN#$
0bHCRMN0_s$sNRRH#NNss$jR5RR0F6F2RVMRH0CCosO;
F0M#NRM0I0H8Es_NsRN$:MRH0s_NsRN$:5=R4.,R,,RcRRg,4RU,d;n2
MOF#M0N0CR8b_0ENNss$RR:H_M0NNss$=R:Rn54d,UcRgU4.c,Rj,gnRc.jU4,Rj,.cR.642O;
F0M#NRM08dHP.RR:HCM0oRCs:5=RI0H8E2-4/;dn
MOF#M0N0HR8PR4n:MRH0CCos=R:RH5I8-0E442/UO;
F0M#NRM08UHPRH:RMo0CC:sR=IR5HE80-/42gO;
F0M#NRM08cHPRH:RMo0CC:sR=IR5HE80-/42cO;
F0M#NRM08.HPRH:RMo0CC:sR=IR5HE80-/42.O;
F0M#NRM084HPRH:RMo0CC:sR=IR5HE80-/424
;
O#FM00NMRFLFD:4RRFLFDMCNRR:=5P8H4RR>j
2;O#FM00NMRFLFD:.RRFLFDMCNRR:=5P8H.RR>j
2;O#FM00NMRFLFD:cRRFLFDMCNRR:=5P8HcRR>j
2;O#FM00NMRFLFD:URRFLFDMCNRR:=5P8HURR>j
2;O#FM00NMRFLFDR4n:FRLFNDCM=R:RH58PR4n>2Rj;F
OMN#0ML0RFdFD.RR:LDFFCRNM:5=R8dHP.RR>j
2;
MOF#M0N0HR8Pd4nU:cRR0HMCsoCRR:=5b8C04E-2n/4d;Uc
MOF#M0N0HR8PgU4.RR:HCM0oRCs:5=R80CbE2-4/gU4.O;
F0M#NRM08cHPjRgn:MRH0CCos=R:RC58b-0E4c2/j;gn
MOF#M0N0HR8Pc.jURR:HCM0oRCs:5=R80CbE2-4/c.jUO;
F0M#NRM084HPjR.c:MRH0CCos=R:RC58b-0E442/j;.c
MOF#M0N0HR8P.64RH:RMo0CC:sR=8R5CEb0-/426;4.
F
OMN#0ML0RF6FD4:.RRFLFDMCNRR:=5P8H6R4.>2Rj;F
OMN#0ML0RF4FDjR.c:FRLFNDCM=R:RH58P.4jcRR>j
2;O#FM00NMRFLFDc.jURR:LDFFCRNM:5=R8.HPjRcU>2Rj;F
OMN#0ML0RFcFDjRgn:FRLFNDCM=R:RH58PgcjnRR>j
2;O#FM00NMRFLFDgU4.RR:LDFFCRNM:5=R8UHP4Rg.>2Rj;F
OMN#0ML0RF4FDncdURL:RFCFDN:MR=8R5HnP4dRUc>2Rj;O

F0M#NRM0#_klI0H8ERR:HCM0oRCs:A=Rm mpqbh'FL#5F4FD2RR+Apmm 'qhb5F#LDFF.+2RRmAmph q'#bF5FLFDRc2+mRAmqp hF'b#F5LF2DURA+Rm mpqbh'FL#5F4FDn
2;O#FM00NMRl#k_b8C0:ERR0HMCsoCRR:=6RR-5mAmph q'#bF5FLFD.642RR+Apmm 'qhb5F#LDFF4cj.2RR+Apmm 'qhb5F#LDFF.Ujc2RR+Apmm 'qhb5F#LDFFcnjg2RR+Apmm 'qhb5F#LDFFU.4g2
2;
MOF#M0N0_RIOHEFOIC_HE80RH:RMo0CC:sR=HRI8_0ENNss$k5#lH_I820E;F
OMN#0MI0R_FOEH_OC80CbERR:HCM0oRCs:8=RCEb0_sNsN#$5kIl_HE802O;
F0M#NRM08E_OFCHO_8IH0:ERR0HMCsoCRR:=I0H8Es_Ns5N$#_kl80CbE
2;O#FM00NMRO8_EOFHCC_8bR0E:MRH0CCos=R:Rb8C0NE_s$sN5l#k_b8C0;E2
F
OMN#0MI0R_8IH0ME_kOl_C#DDRH:RMo0CC:sR=IR5HE80-/42IE_OFCHO_8IH0+ERR
4;O#FM00NMR8I_CEb0_lMk_DOCD:#RR0HMCsoCRR:=5b8C04E-2_/IOHEFO8C_CEb0R4+R;O

F0M#NRM08H_I8_0EM_klODCD#RR:HCM0oRCs:5=RI0H8E2-4/O8_EOFHCH_I8R0E+;R4
MOF#M0N0_R880CbEk_MlC_ODRD#:MRH0CCos=R:RC58b-0E482/_FOEH_OC80CbERR+4
;
O#FM00NMR#I_HRxC:MRH0CCos=R:RII_HE80_lMk_DOCD*#RR8I_CEb0_lMk_DOCD
#;O#FM00NMR#8_HRxC:MRH0CCos=R:RI8_HE80_lMk_DOCD*#RR88_CEb0_lMk_DOCD
#;
MOF#M0N0FRLF8D_RL:RFCFDN:MR=8R5_x#HCRR-IH_#x<CR=2Rj;F
OMN#0ML0RF_FDIRR:LDFFCRNM:M=RFL05F_FD8
2;
MOF#M0N0EROFCHO_8IH0:ERR0HMCsoCRR:=5mAmph q'#bF5FLFD2_8R8*R_FOEH_OCI0H8E+2RRm5Amqp hF'b#F5LFID_2RR*IE_OFCHO_8IH0;E2
MOF#M0N0EROFCHO_b8C0:ERR0HMCsoCRR:=5mAmph q'#bF5FLFD2_8R8*R_FOEH_OC80CbE+2RRm5Amqp hF'b#F5LFID_2RR*IE_OFCHO_b8C0;E2
MOF#M0N0HRI8_0EM_klODCD#RR:HCM0oRCs:5=RApmm 'qhb5F#LDFF_R82*H5I8-0E482/_FOEH_OCI0H8E+2RRm5Amqp hF'b#F5LFID_2RR*58IH04E-2_/IOHEFOIC_HE802RR+4O;
F0M#NRM080CbEk_MlC_ODRD#:MRH0CCos=R:Rm5Amqp hF'b#F5LF8D_25R*80CbE2-4/O8_EOFHCC_8b20ER5+RApmm 'qhb5F#LDFF_RI2*8R5CEb0-/42IE_OFCHO_b8C0RE2+;R4
O--F0M#NRM0M_klODCD#RR:HCM0oRCs:5=R5C58bR0E-2R4Rd/R.+2RR55580CbERR-4l2RFd8R./2RR24n2R;RRR--yVRFRv)qd4.X1CRODRD#M8CCC
8R-F-OMN#0MD0RC_V0FsPCRH:RMo0CC:sR=5R55b8C0+ERR246R8lFR2d.R4/RnR2;RRRRRRRRRRRRRRRRRRRRRRRR-y-RRRFV)4qvn1X4RCMC8RC8VRFsD0CVRCFPsFRIs
8#0C$bR0Fk_#Lk4$_0bHCR#sRNsRN$5b8C0ME_kOl_C#DD-84RF0IMF,RjR8IH0ME_kOl_C#DD-84RF0IMF2RjRRFV#_08DHFoO#;
HNoMDkRF0k_L#:4RR0Fk_#Lk4$_0bRC;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RV_Rs80FkRM5HbRk000FRs#H-0CN0#02
$RbCF_k0L.k#_b0$C#RHRsNsN5$R80CbEk_MlC_OD-D#4FR8IFM0RRj,.H*I8_0EM_klODCD#R+48MFI0jFR2VRFR8#0_oDFH
O;#MHoNFDRkL0_kR#.:kRF0k_L#0._$;bCRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$FsVR_k8F0HR5M0bkRR0F0-sH#00NC
#20C$bR0Fk_#Lkc$_0bHCR#sRNsRN$5b8C0ME_kOl_C#DD-84RF0IMF,RjRIc*HE80_lMk_DOCDd#+RI8FMR0FjF2RV0R#8F_Do;HO
o#HMRNDF_k0Lck#RF:RkL0_k_#c0C$b;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFVsF_8k50RHkMb0FR0RH0s-N#002C#
b0$CkRF0k_L#0U_$RbCHN#Rs$sNRC58b_0EM_klODCD#R-48MFI0jFR,*RUI0H8Ek_MlC_OD+D#(FR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNR0Fk_#LkURR:F_k0LUk#_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFR8s_FRk05bHMk00RFsR0H0-#N#0C2$
0bbCRN0sH$k_L#0U_$RbCHN#Rs$sNRC58b_0EM_klODCD#R-48MFI0jFR,HRI8_0EM_klODCD#R-48MFI0jFR2VRFR8#0_oDFH
O;#MHoNbDRN0sH$k_L#:URRsbNH_0$LUk#_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$FsVR_k8F0HR5M0bkRR0F0-sH#00NC
#20C$bR0Fk_#Lk40n_$RbCHN#Rs$sNRC58b_0EM_klODCD#R-48MFI0jFR,nR4*8IH0ME_kOl_C#DD+R468MFI0jFR2VRFR8#0_oDFH
O;#MHoNFDRkL0_kn#4RF:RkL0_kn#4_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFR8s_FRk05bHMk00RFsR0H0-#N#0C2$
0bbCRN0sH$k_L#_4n0C$bRRH#NNss$8R5CEb0_lMk_DOCD4#-RI8FMR0Fj.,R*8IH0ME_kOl_C#DD+84RF0IMF2RjRRFV#_08DHFoO#;
HNoMDNRbs$H0_#Lk4:nRRsbNH_0$L4k#n$_0bRC;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFVsF_8k50RHkMb0FR0RH0s-N#002C#
b0$CkRF0k_L#_d.0C$bRRH#NNss$8R5CEb0_lMk_DOCD4#-RI8FMR0Fjd,R.H*I8_0EM_klODCD#4+dRI8FMR0FjF2RV0R#8F_Do;HO
o#HMRNDF_k0Ldk#.RR:F_k0Ldk#.$_0bRC;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RV_Rs80FkRM5HbRk000FRs#H-0CN0#02
$RbCbHNs0L$_k.#d_b0$C#RHRsNsN5$R80CbEk_MlC_OD-D#4FR8IFM0RRj,cH*I8_0EM_klODCD#R+d8MFI0jFR2VRFR8#0_oDFH
O;#MHoNbDRN0sH$k_L#Rd.:NRbs$H0_#Lkd0._$;bCRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFR8s_FRk05bHMk00RFsR0H0-#N#0C2H
#oDMNR0Fk_RCM:0R#8F_Do_HOP0COF8s5CEb0_lMk_DOCD4#-RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-C-RMDNLCV#RF0sRs#H-0CN0#H
#oDMNR0Is_RCM:0R#8F_Do_HOP0COF8s5CEb0_lMk_DOCD4#-RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-I-RsCH0RNCML#DCRsVFROCNEFRsIVRFRv)qRDOCD##
HNoMDMRH_osCR#:R0D8_FOoH_OPC05FsI0H8E6+dRI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RCk#8FR0RosCHC#0sQR7h#R
HNoMDkRF0C_soRR:#_08DHFoOC_POs0F58IH0dE+6FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RCk#8FR0RosCHC#0smR7z#a
HNoMDkRF0C_so:4RR8#0_oDFHPO_CFO0sH5I8-0E4FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--k8#CRR0FOFEF#LCRCC0IC7MRQNhRMF8Rkk0b0VRFRFADO)	Rq#v
HNoMD8RN_osCR#:R0D8_FOoH_OPC05FsNs88I0H8ER-48MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--k8#CRR0FsHCo#s0CR7q7)FRVssRIH
0C#MHoNDDRFsI_Ns88R#:R0D8_FOoH_OPC05Fs48dRF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-s-RNs88R0LH#MRHbRk00)FRqOvRC#DDRR5cL#H0RJsCkCHs8#2
HNoMDFRDIN_I8R8s:0R#8F_Do_HOP0COF4s5dFR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-NRI8R8sL#H0RbHMk00RFqR)vCRODRD#5LcRHR0#skCJH8sC2H
#oDMNR7)q70)_l:bRR8#0_oDFHPO_CFO0s85N8HsI8-0E4FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-#RkC08RFHRbbHCDM)CRq)77
o#HMRNDW7q7)l_0bRR:#_08DHFoOC_POs0F58N8s8IH04E-RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RCk#8FR0RbbHCMDHCqRW7
7)#MHoN7DRQ0h_l:bRR8#0_oDFHPO_CFO0sH5I8-0E4FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--k8#CRR0FbCHbDCHMRh7Q
o#HMRNDW0 _l:bRR8#0_oDFHRO;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-#RkC08RFHRbbHCDMWCR -
-R8CMRFLDOs	RNHlRlCbDl0CMNF0HMHR#oDMN#-

-CRLoRHM#CCDOs0RNHlRlCbDl0CMNF0HMHR#oDMN#$
0bDCRCFV0P_Cs0#RHRsNsN5$RjFR0RRd2FHVRMo0CC
s;0C$bRVDC0CFPs__0.#RHRsNsN5$RjFR0RR42FHVRMo0CC
s;VOkM0MHFR8bN5:HRR8#0_oDFHPO_CFO0sI;R4I,R.RR:HCM0o2CsR0sCkRsM#_08DHFoOC_POs0FR
H#PHNsNCLDRsPNR#:R0D8_FOoH_OPC05FsI44-RI8FMR0Fj
2;LHCoMR
RVRFs[MRHRsPN'MsNoDCRF
FbRRRRH5VR[=R<R2I.RC0EMSR
RNRPs25[RR:=H'5HD+FI[
2;S#CDCR
SRsPN5R[2:'=Rj
';S8CMR;HV
CRRMD8RF;Fb
sRRCs0kMNRPsC;
Mb8RN
8;VOkM0MHFR0oC_8IH0UE_58IH0RE:HCM0o2CsR0sCkRsMHCM0oRCsHP#
NNsHLRDCPRND:MRH0CCos=R:R
j;LHCoMR
RPRND:I=RHE80/
U;RVRHRI55HE80R8lFRRU2>2RcRC0EMR
RRNRPD=R:RDPNR4+R;R
RCRM8H
V;RCRs0MksRDPN;M
C8CRo0H_I8_0EUV;
k0MOHRFMo_C0I0H8E5_.I0H8EH:RMo0CCRs2skC0sHMRMo0CCHsR#N
PsLHNDPCRN:DRR0HMCsoCRR:=jL;
CMoH
PRRN:DR=HRI8/0E.R;
R0sCkRsMP;ND
8CMR0oC_8IH0.E_;k
VMHO0FoMRCI0_HE8058IH0:ERR0HMCsoC2CRs0MksRVDC0CFPs__0.#RH
sPNHDNLCNRPDRR:D0CVFsPC_.0_;C
Lo
HMRNRPD254RR:=o_C0I0H8E5_.I0H8E
2;RVRHRH5I8R0ElRF8.RR=j02RE
CMRRRRP5NDj:2R=;Rj
CRRD
#CRRRRP5NDj:2R=;R4
CRRMH8RVR;
R0sCkRsMP;ND
8CMR0oC_8IH0
E;VOkM0MHFR0oC_8IH0IE5HE80RH:RMo0CCRs2skC0sDMRCFV0P_Cs0#RH
sPNHDNLCNRPDRR:D0CVFsPC_:0R=jR5,,RjRRj,j
2;LHCoMR
RP5NDd:2R=CRo0H_I8_0EUH5I820E;R
ROCN#RH5I8R0ElRF8UH2R#R
RIMECR|cRR=dR>NRPD25.RR:=4R;
RCIEMRR.=P>RN4D52=R:R
4;RERIC4MRRR=>P5NDj:2R=;R4
IRRERCMFC0Es=#R>kRMD
D;RMRC8NRO#
C;RCRs0MksRDPN;M
C8CRo0H_I8;0E
MOF#M0N0_R#I0H8Es_NsRN$:CRDVP0FC0s_RR:=o_C0I0H8EH5I820E;F
OMN#0M#0R_8IH0NE_s$sN_Rnc:CRDVP0FC0s__:.R=CRo0H_I850EI0H8E
2;VOkM0MHFR0oC_lMk_U4.5b8C0RE:HCM0o2CsR0sCkRsMHCM0oRCsHP#
NNsHLRDCPRND:MRH0CCos=R:R
j;LHCoMR
RPRND:8=RCEb0/U4.;R
RH5VR5b8C0lERF48R.RU2>4R4.02RE
CMRRRRPRND:P=RN+DRR
4;RMRC8VRH;R
RskC0sPMRN
D;CRM8o_C0M_kl4;.U
MVkOF0HMCRo0C_DVP0FCns_cC58bR0E:MRH0CCoss2RCs0kMMRH0CCos#RH
oLCHRM
R0sCk5sM80CbEFRl8.R4U
2;CRM8o_C0D0CVFsPC_;nc
MVkOF0HMCRo0k_Mlc_n5b8C0:ERR0HMCsoC2CRs0MksR0HMCsoCR
H#PHNsNCLDRDPNRH:RMo0CC:sR=;Rj
oLCHRM
RVRHRC58bR0E<4=R4N.RM88RCEb0Rc>RU02RE
CMRRRRRDPNRR:=4R;
R8CMR;HV
sRRCs0kMNRPDC;
Mo8RCM0_knl_cV;
k0MOHRFMo_C0D0CVFsPC5b8C0:ERR0HMCsoC;NRlGRR:HCM0o2CsR0sCkRsMHCM0oRCsHP#
NNsHLRDCPRND:MRH0CCos=R:R
j;LHCoMR
RH5VR80CbERR-lRNG>j=R2ER0CRM
RPRRN:DR=CR8bR0E-NRlGR;
R#CDCR
RRNRPD=R:Rb8C0
E;RMRC8VRH;R
RskC0sPM5N;D2
8CMR0oC_VDC0CFPsV;
k0MOHRFMo_C0M_kld8.5CEb0RH:RMo0CCRs2skC0sHMRMo0CCHsR#N
PsLHNDPCRN:DRR0HMCsoCRR:=jL;
CMoH
HRRV8R5CEb0RR<=cNURM88RCEb0R4>Rn02RE
CMRRRRRDPNRR:=4R;
R8CMR;HV
sRRCs0kMNRPDC;
Mo8RCM0_kdl_.V;
k0MOHRFMo_C0M_kl48n5CEb0RH:RMo0CCRs2skC0sHMRMo0CCHsR#N
PsLHNDPCRN:DRR0HMCsoCRR:=jL;
CMoH
HRRV8R5CEb0RR<=4NnRM88RCEb0Rj>R2ER0CRM
RRRRPRND:4=R;R
RCRM8H
V;RCRs0MksRDPN;M
C8CRo0k_Mln_4;-
-O#FM00NMRlMk_DOCD:#RR0HMCsoCRR:=5855CEb0R4-R2RR/dR.2+5R55b8C0-ERRR42lRF8dR.2/nR42R2;R-R-RFyRVqR)vXd.4O1RC#DDRCMC8RC8
MOF#M0N0kRMlC_OD4D_.:URR0HMCsoCRR:=o_C0M_kl45.U80CbE
2;O#FM00NMRVDC0CFPsc_nRH:RMo0CC:sR=CRo0C_DVP0FCns_cC58b20E;F
OMN#0MM0RkOl_C_DDn:cRR0HMCsoCRR:=o_C0M_klnDc5CFV0P_Csn;c2
MOF#M0N0CRDVP0FCds_.RR:HCM0oRCs:o=RCD0_CFV0P5CsD0CVFsPC_,ncR2nc;F
OMN#0MM0RkOl_C_DDd:.RR0HMCsoCRR:=o_C0M_kldD.5CFV0P_Csd;.2
MOF#M0N0CRDVP0FC4s_nRR:HCM0oRCs:o=RCD0_CFV0P5CsD0CVFsPC_,d.R2d.;F
OMN#0MM0RkOl_C_DD4:nRR0HMCsoCRR:=o_C0M_kl4Dn5CFV0P_Cs4;n2
$
0bFCRkL0_k0#_$_bC4R.UHN#Rs$sNRk5MlC_OD4D_.8URF0IMF,RjR8IH04E-RI8FMR0FjF2RV0R#8F_Do;HO
b0$CkRF0k_L#$_0bnC_c#RHRsNsN5$RM_klODCD_Rnc8MFI0jFR,HRI8-0E4FR8IFM0RRj2F#VR0D8_FOoH;$
0bFCRkL0_k0#_$_bCdH.R#sRNsRN$5lMk_DOCD._dRI8FMR0FjI,RHE80-84RF0IMF2RjRRFV#_08DHFoO0;
$RbCF_k0L_k#0C$b_R4nHN#Rs$sNRk5MlC_OD4D_nFR8IFM0RRj,I0H8ER-48MFI0jFR2VRFR8#0_oDFH
O;#MHoNFDRkL0_k4#_.:URR0Fk_#Lk_b0$C._4UR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFRk8F0HR5M0bkRR0F0-sH#00NC
#2#MHoNFDRkL0_kn#_cRR:F_k0L_k#0C$b_;ncRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$F8VRFRk05bHMk00RFsR0H0-#N#0C2H
#oDMNR0Fk_#Lk_Rd.:kRF0k_L#$_0bdC_.R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFRk8F0HR5M0bkRR0F0-sH#00NC
#2#MHoNFDRkL0_k4#_nRR:F_k0L_k#0C$b_;4nRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$F8VRFRk05bHMk00RFsR0H0-#N#0C2H
#oDMNRF#_kC0_MRR:#_08DHFoOC_POs0F5lMk_DOCD._4UFR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--CLMNDRC#VRFs0-sH#00NC##
HNoMDkRF0M_C_Rnc:0R#8F_Do;HO
o#HMRNDF_k0CdM_.RR:#_08DHFoO#;
HNoMDkRF0M_C_R4n:0R#8F_Do;HO
o#HMRND#s_I0M_CR#:R0D8_FOoH_OPC05FsM_klODCD_U4.RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-I-RsCH0RNCML#DCRsVFROCNEFRsIVRFRv)qRDOCD##
HNoMDsRI0M_C_Rnc:0R#8F_Do;HO
o#HMRNDI_s0CdM_.RR:#_08DHFoO#;
HNoMDsRI0M_C_R4n:0R#8F_Do;HO
o#HMRND#M_H_osCR#:R0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--k8#CRR0FsHCo#s0CRh7QRH
#oDMNRF#_ks0_C:oRR8#0_oDFHPO_CFO0sH5I8-0E4FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RCk#8FR0RosCHC#0smR7z#a
HNoMD_R#Ns8_C:oRR8#0_oDFHPO_CFO0s85N8HsI8-0E4FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-#RkC08RFCRso0H#CqsR7
7)#MHoNDDRFNI_8R8s:0R#8F_Do_HOP0COFns5RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-R8N8sHRL0H#RM0bkRR0F)RqvODCD#cR5R0LH#CRsJskHC
82O#FM00NMRLD#_8IH0:ERR0HMCsoCRR:=I0H8E*-U5I#_HE80_sNsNd$522-4-#c*_8IH0NE_s$sN5-.2._*#I0H8Es_Ns5N$4#2-_8IH0NE_s$sN5;j2
b0$ClR0bs_NsUN$RRH#NNss$#R5_8IH0NE_s$sN5-d24FR8IFM0RRj2F#VR0D8_FOoH_OPC05Fs(FR8IFM0R;j2
o#HMRND0_lbU._d,lR0b__U4:nRRb0l_sNsN;$U
R--CRM8#CCDOs0RNHlRlCbDl0CMNF0HMHR#oDMN#0
N0LsHkR0C\N3slV_FV0#C\RR:#H0sM
o;
oLCHRM
RR
RzRcd:VRHR85N8ss_CRo2oCCMsCN0RR--oCCMsCN0RFLDOs	RNRl
R-RR-VRQR8N8s8IH0<ERRFOEH_OCI0H8E#RN#MHoR''jRR0Fk#MkCL8RH
0#RRRRzRjR:VRHR85N8HsI8R0E=2R4RMoCC0sNCR
RRRRRRFRDIN_s8R8s<"=Rjjjjjjjjjjjjj&"RR7q7)25j;R
RRRRRRFRDIN_I8R8s<"=Rjjjjjjjjjjjjj&"RR_N8s5Coj
2;RRRRCRM8oCCMsCN0R;zj
RRRRRz4RH:RVNR58I8sHE80R.=R2CRoMNCs0RC
RRRRRDRRFsI_Ns88RR<="jjjjjjjjjjjj&"RR7q7)R548MFI0jFR2R;
RRRRRDRRFII_Ns88RR<="jjjjjjjjjjjj&"RR_N8s5Co4FR8IFM0R;j2
RRRR8CMRMoCC0sNC4Rz;R
RR.RzRRR:H5VRNs88I0H8ERR=do2RCsMCN
0CRRRRRRRRD_FIs8N8s=R<Rj"jjjjjjjjjj&"RR7q7)R5.8MFI0jFR2R;
RRRRRDRRFII_Ns88RR<="jjjjjjjjjjj"RR&Ns8_C.o5RI8FMR0Fj
2;RRRRCRM8oCCMsCN0R;z.
RRRRRzdRH:RVNR58I8sHE80Rc=R2CRoMNCs0RC
RRRRRDRRFsI_Ns88RR<="jjjjjjjj"jjRq&R757)dFR8IFM0R;j2
RRRRRRRRIDF_8IN8<sR=jR"jjjjjjjjj&"RR_N8s5CodFR8IFM0R;j2
RRRR8CMRMoCC0sNCdRz;R
RRcRzRRR:H5VRNs88I0H8ERR=6o2RCsMCN
0CRRRRRRRRD_FIs8N8s=R<Rj"jjjjjj"jjRq&R757)cFR8IFM0R;j2
RRRRRRRRIDF_8IN8<sR=jR"jjjjjjjj"RR&Ns8_Cco5RI8FMR0Fj
2;RRRRCRM8oCCMsCN0R;zc
RRRRRz6RH:RVNR58I8sHE80Rn=R2CRoMNCs0RC
RRRRRDRRFsI_Ns88RR<="jjjjjjjj&"RR7q7)R568MFI0jFR2R;
RRRRRDRRFII_Ns88RR<="jjjjjjjj&"RR_N8s5Co6FR8IFM0R;j2
RRRR8CMRMoCC0sNC6Rz;R
RRnRzRRR:H5VRNs88I0H8ERR=(o2RCsMCN
0CRRRRRRRRD_FIs8N8s=R<Rj"jjjjjj&"RR7q7)R5n8MFI0jFR2R;
RRRRRDRRFII_Ns88RR<="jjjjjjj"RR&Ns8_Cno5RI8FMR0Fj
2;RRRRCRM8oCCMsCN0R;zn
RRRRRz(RH:RVNR58I8sHE80RU=R2CRoMNCs0RC
RRRRRDRRFsI_Ns88RR<="jjjj"jjRq&R757)(FR8IFM0R;j2
RRRRRRRRIDF_8IN8<sR=jR"jjjjj&"RR_N8s5Co(FR8IFM0R;j2
RRRR8CMRMoCC0sNC(Rz;R
RRURzRRR:H5VRNs88I0H8ERR=go2RCsMCN
0CRRRRRRRRD_FIs8N8s=R<Rj"jj"jjRq&R757)UFR8IFM0R;j2
RRRRRRRRIDF_8IN8<sR=jR"jjjj"RR&Ns8_CUo5RI8FMR0Fj
2;RRRRCRM8oCCMsCN0R;zU
RRRRRzgRH:RVNR58I8sHE80R4=Rjo2RCsMCN
0CRRRRRRRRD_FIs8N8s=R<Rj"jjRj"&7Rq7g)5RI8FMR0Fj
2;RRRRRRRRD_FII8N8s=R<Rj"jjRj"&8RN_osC58gRF0IMF2Rj;R
RRMRC8CRoMNCs0zCRgR;
RzRR4RjR:VRHR85N8HsI8R0E=4R42CRoMNCs0RC
RRRRRDRRFsI_Ns88RR<="jjj"RR&q)775R4j8MFI0jFR2R;
RRRRRDRRFII_Ns88RR<="jjj"RR&Ns8_C4o5jFR8IFM0R;j2
RRRR8CMRMoCC0sNC4RzjR;
RzRR4R4R:VRHR85N8HsI8R0E=.R42CRoMNCs0RC
RRRRRDRRFsI_Ns88RR<=""jjRq&R757)484RF0IMF2Rj;R
RRRRRRFRDIN_I8R8s<"=RjRj"&8RN_osC5R448MFI0jFR2R;
RCRRMo8RCsMCNR0Cz;44
RRRR.z4RRR:H5VRNs88I0H8ERR=4Rd2oCCMsCN0
RRRRRRRRIDF_8sN8<sR=jR''RR&q)775R4.8MFI0jFR2R;
RRRRRDRRFII_Ns88RR<='Rj'&8RN_osC5R4.8MFI0jFR2R;
RCRRMo8RCsMCNR0Cz;4.
RRRRdz4RRR:H5VRNs88I0H8ERR>4Rd2oCCMsCN0
RRRRRRRRIDF_8sN8<sR=7Rq74)5dFR8IFM0R;j2
RRRRRRRRIDF_8IN8<sR=8RN_osC5R4d8MFI0jFR2R;
RCRRMo8RCsMCNR0Cz;4d
R
RR-R-RRQV5M8H_osC2CRso0H#C7sRQkhR#oHMRiBp
RRRRcz4RRR:H5VR8_HMs2CoRMoCC0sNCR
RRRRRRsRbF#OC#BR5pRi,72QhRoLCHRM
RRRRRRRRRHRRVBR5p=iRR''4R8NMRiBp'CCPMR020MEC
RRRRRRRRRRRRRRRR_HMsRCo<5=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj&"RRh7Q2R;
RRRRRRRRRCRRMH8RVR;
RRRRRCRRMb8RsCFO#
#;RRRRCRM8oCCMsCN0Rcz4;R
RR4Rz6:RRRRHV50MFRM8H_osC2CRoMNCs0RC
RRRRRRRRRHRRMC_so=R<Rj5"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jjR7&RQ;h2
RRRR8CMRMoCC0sNC4Rz6
;
RRRR-Q-RVsR580Fk_osC2CRso0H#C)sR_z7ma#RkHRMo)B_mpRi
RzRR4RnR:VRHRF58ks0_CRo2oCCMsCN0
RRRRRRRRFbsO#C#RB5mpRi,F_k0s4Co2CRLo
HMRRRRRRRRRRRRH5VRmiBpR'=R4N'RMm8RB'piCMPC002RE
CMRRRRRRRRRRRRRRRR7amzRR<=F_k0s4Co;R
RRRRRRRRRRMRC8VRH;R
RRRRRRMRC8sRbF#OC#R;
RRRRRCRRMo8RCsMCNR0Cz;4n
RRRR(z4RRR:H5VRMRF080Fk_osC2CRoMNCs0RC
RRRRRRRRR7RRmRza<F=Rks0_C;o4
RRRR8CMRMoCC0sNC4Rz(
;
RRRR-Q-RVNR58_8ss2CoRosCHC#0s7Rq7V)RFIsRsCH0RHk#MBoRpRi
RzRR4RUIRH:RVNR58_8ss2CoRMoCC0sNCR
RRRRRRsRbF#OC#BR5pRi,q)772CRLo
HMRRRRRRRRRRRRH5VRBRpi=4R''MRN8pRBiP'CC2M0RC0EMR
RRRRRRRRRRRRRR8RN_osCRR<=q)7758N8s8IH04E-RI8FMR0Fj
2;RRRRRRRRRRRRCRM8H
V;RRRRRRRRCRM8bOsFC;##
RRRR8CMRMoCC0sNC4RzU
I;RRRRzI4gRH:RVMR5FN0R8_8ss2CoRMoCC0sNCR
RRRRRRRRRR8RN_osCRR<=q)77;R
RRMRC8CRoMNCs0zCR4;gI
R
RR-R-R0 GsDNRFOoHRsVFRN7kDFRbsO0RN
#CRRRRzosCRb:RsCFO#B#5pRi2LHCoMR
RRRRRH5VRB'pi he aMRN8pRBiRR='24'RC0EMR
RRRRRRh7Q_b0lRR<=7;Qh
RRRRRRR)7q7)l_0b=R<R7q7)R;
RRRRRqRW7_7)0Rlb<N=R8C_soR;
RRRRR RW_b0lRR<=W
 ;RRRRRMRC8VRH;R
RRMRC8sRbF#OC#
;
RRRR-Q-RVCR)Nq8R8C8s#=#RRHWs0qCR8C8s#R#,LN$b#7#RQ0hRFkRF00bkRRHVWH R#MRCNCLD8R
RRlRzk:GRRFbsO#C#5_W 0,lbR7)q70)_lRb,W7q7)l_0b7,RQ0h_lRb,F_k0s2Co
RRRRLRRCMoH
RRRRRRRRRHV57Wq70)_l=bRR7)q70)_lNbRMW8R l_0bRR='24'RC0EMR
RRRRRRRRRF_k0s4CoRR<=7_Qh0;lb
RRRRRRRR#CDCR
RRRRRRRRRF_k0s4CoRR<=F_k0s5CoI0H8ER-48MFI0jFR2R;
RRRRRCRRMH8RVR;
RCRRMb8RsCFO#
#;RRRRRRRR
RRRRR--tCCMsCN0RC0ERv)qRDOCDN#RM#8RCODC0FRDoRHOVRFs)Aqv41n_44_1
RRRRUz4RH:RVOR5EOFHCH_I8R0E=2R4RMoCC0sNCR
RRRRRR4RzgRR:VRFsHMRHRC58b_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
RRRRR--Q5VRNs88I0H8ERR>4Rc2M8CCRR0FONsC0ICRsCH0RNCMLRDCNRM8Fbk0kC0RMDNLCCR#D0CORoDFHRO
RRRRRRRRRzRR.:jRRRHV58N8s8IH0>ERR24cRMoCC0sNCR
RRRRRRRRRRRRRRkRF0M_C5RH2<'=R4I'RERCM57)q70)_lNb58I8sHE80-84RF0IMFcR42RR=HC2RDR#C';j'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RWRCIEMNR58C_so85N8HsI8-0E4FR8IFM0R24cRH=R2DRC#'CRj
';RRRRRRRRRRRRCRM8oCCMsCN0Rjz.;R
RR-R-RRQV58N8s8IH0<ER=.R42FRMRHIs0CCRMDNLCsRFR0FkbRk0CLMND#CRCODC0FRDoRHOM8CCCR8
RRRRRRRRRzRR.:4RRRHV58N8s8IH0<ER=cR42CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_M25HRR<=';4'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RW;R
RRRRRRRRRRMRC8CRoMNCs0zCR.
4;RRRR-t-RCsMCNR0C0REC)RqvODCD#MRN8sR0H0-#N#0C
RRRRRRRRRRRR.z.RV:RF[sRRRHM58IH0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CRRRRRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FAVR)_qv4Undc7X4RD:RNDLCRRH#";W"
RRRRRRRRRRRRRRRRoLCHRM
RRRRRRRRRRRRRARR)_qv4Undc7X4R):Rq4vAn4_1_
14RRRRRRRRRRRRRRRRb0FsRblNRQ57q25jRR=>HsM_C[o52q,R7q7)RR=>D_FII8N8sd54RI8FMR0FjR2,7RQA=">RjR",q)77A>R=RIDF_8sN84s5dFR8IFM0R,j2
RRRRRRRRRRRRRRRRq hRR=>',4'R)11q>R=R''j, RWq>R=R0Is_5CMHR2,BqpiRR=>B,piRA hRR=>',4'R)11A>R=R''j, RWA>R=R''j,pRBi=AR>pRBiR,
RRRRRRRRRRRRR7RRm=qR>bRFCRM,75mAj=2R>kRF0k_L#H45,2[2;R

RRRRRRRRRRRRRFRRks0_C[o52=R<R0Fk_#Lk4,5H[I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRCRM8oCCMsCN0R.z.;R
RRRRRRMRC8CRoMNCs0zCR4
g;RRRRCRM8oCCMsCN0RUz4;RRRRR
RRRRR
RRRRR--tCCMsCN0RC0ERv)qRDOCDN#RM#8RCODC0FRDoRHOVRFs)Aqv41n_.._1
RRRRdz.RH:RVOR5EOFHCH_I8R0E=2R.RMoCC0sNCR
RRRRRR.RzcRR:VRFsHMRHRC58b_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
RRRRR--Q5VRNs88I0H8ERR>4Rd2M8CCRR0FONsC0ICRsCH0RNCMLRDCNRM8Fbk0kC0RMDNLCCR#D0CORoDFHRO
RRRRRRRRRzRR.:6RRRHV58N8s8IH0>ERR24dRMoCC0sNCR
RRRRRRRRRRRRRRkRF0M_C5RH2<'=R4I'RERCM57)q70)_lNb58I8sHE80-84RF0IMFdR42RR=HC2RDR#C';j'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RWRCIEMNR58C_so85N8HsI8-0E4FR8IFM0R24dRH=R2DRC#'CRj
';RRRRRRRRRRRRCRM8oCCMsCN0R6z.;R
RR-R-RRQV58N8s8IH0<ER=dR42FRMRHIs0CCRMDNLCsRFR0FkbRk0CLMND#CRCODC0FRDoRHOM8CCCR8
RRRRRRRRRzRR.:nRRRHV58N8s8IH0<ER=dR42CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_M25HRR<=';4'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RW;R
RRRRRRRRRRMRC8CRoMNCs0zCR.
n;RRRR-t-RCsMCNR0C0REC)RqvODCD#MRN8sR0H0-#N#0C
RRRRRRRRRRRR(z.RV:RF[sRRRHM58IH0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CRRRRRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FAVR)_qvU.4gXR.7:NRDLRCDH"#RW
";RRRRRRRRRRRRRRRRLHCoMR
RRRRRRRRRRRRRR)RAqUv_4Xg..:7RRv)qA_4n11._.R
RRRRRRRRRRRRRRFRbsl0RN5bR7RQq=H>RMC_so*5.[R+48MFI0.FR*,[2R7q7)=qR>FRDIN_I858s48.RF0IMF2Rj,QR7A>R=Rj"j"q,R7A7)RR=>D_FIs8N8s.54RI8FMR0Fj
2,RRRRRRRRRRRRRRRR Rhq='>R4R',1q1)RR=>',j'RqW RR=>I_s0CHM52B,RpRiq=B>RpRi, RhA='>R4R',1A1)RR=>',j'RAW RR=>',j'RiBpA>R=RiBp,R
RRRRRRRRRRRRRRmR7q>R=RCFbM7,Rm4A52>R=R0Fk_#Lk.,5H.+*[4R2,75mAj=2R>kRF0k_L#H.5,*R.[;22
RRRRRRRRRRRRRRRR0Fk_osC5[.*2=R<R0Fk_#Lk.,5H.2*[RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so*5.[2+4RR<=F_k0L.k#5.H,*4[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRCRRMo8RCsMCNR0Cz;.(
RRRRRRRR8CMRMoCC0sNC.RzcR;
RCRRMo8RCsMCNR0Cz;.dR
R
RRRRRRRR-t-RCsMCNR0C0REC)RqvODCD#MRN8CR#D0CORoDFHVORF)sRq4vAnc_1_
1cRRRRzR.U:VRHRE5OFCHO_8IH0=ERRRc2oCCMsCN0
RRRRRRRRgz.RV:RFHsRRRHM5b8C0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CRRRR-Q-RVNR58I8sHE80R4>R.M2RCRC80OFRs0CNCsRIHR0CCLMNDNCRMF8Rkk0b0MRCNCLDRD#CCRO0DHFoOR
RRRRRRRRRRdRzjRR:H5VRNs88I0H8ERR>4R.2oCCMsCN0
RRRRRRRRRRRRRRRR0Fk_5CMH<2R=4R''ERIC5MR)7q7)l_0b85N8HsI8-0E4FR8IFM0R24.RH=R2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0CHM52=R<RRW IMECR85N_osC58N8s8IH04E-RI8FMR0F4R.2=2RHR#CDCjR''R;
RRRRRRRRRCRRMo8RCsMCNR0Cz;dj
RRRRR--Q5VRNs88I0H8E=R<R24.RRMFI0sHCMRCNCLDRRFsFbk0kC0RMDNLCCR#D0CORoDFHMORCCC88R
RRRRRRRRRRdRz4RR:H5VRNs88I0H8E=R<R24.RMoCC0sNCR
RRRRRRRRRRRRRRkRF0M_C5RH2<'=R4
';RRRRRRRRRRRRRRRRI_s0CHM52=R<R;W 
RRRRRRRRRRRR8CMRMoCC0sNCdRz4R;
R-RR-CRtMNCs00CRE)CRqOvRC#DDR8NMRH0s-N#00
C#RRRRRRRRRRRRzRd.:FRVsRR[H5MRI0H8Ek_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0RC
RRRRRRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)RAqcv_jXgnc:7RRLDNCHDR#WR""R;
RRRRRRRRRRRRRLRRCMoH
RRRRRRRRRRRRRRRRqA)vj_cgcnX7RR:)Aqv41n_cc_1
RRRRRRRRRRRRRRRRsbF0NRlb7R5Q=qR>MRH_osC5[c*+8dRF0IMF*Rc[R2,q)77q>R=RIDF_8IN84s54FR8IFM0R,j2RA7QRR=>"jjjjR",q)77A>R=RIDF_8sN84s54FR8IFM0R,j2
RRRRRRRRRRRRRRRRq hRR=>',4'R)11q>R=R''j, RWq>R=R0Is_5CMHR2,BqpiRR=>B,piRA hRR=>',4'R)11A>R=R''j, RWA>R=R''j,pRBi=AR>pRBiR,
RRRRRRRRRRRRR7RRm=qR>bRFCRM,75mAd=2R>kRF0k_L#Hc5,*Rc[2+d,mR7A25.RR=>F_k0Lck#5cH,*.[+2
,RRRRRRRRRRRRRRRRR75mA4=2R>kRF0k_L#Hc5,[c*+,42RA7m5Rj2=F>RkL0_k5#cHc,R*2[2;R
RRRRRRRRRRRRRRkRF0C_so*5c[<2R=kRF0k_L#Hc5,[c*2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cco5*4[+2=R<R0Fk_#Lkc,5Hc+*[4I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Coc+*[.<2R=kRF0k_L#Hc5,[c*+R.2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5[c*+Rd2<F=RkL0_k5#cH*,c[2+dRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R

RRRRRRRRRCRRMo8RCsMCNR0Cz;d.
RRRRRRRR8CMRMoCC0sNC.RzgR;
RCRRMo8RCsMCNR0Cz;.U
R
RRRRRR-R-RMtCC0sNCER0CqR)vCRODRD#NRM8#CCDOD0RFOoHRsVFRv)qA_4n11g_gR
RRdRzdRR:H5VROHEFOIC_HE80Rg=R2CRoMNCs0RC
RRRRRzRRd:cRRsVFRHHRM8R5CEb0_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNCR
RR-R-RRQV58N8s8IH0>ERR244RCMC8FR0RCOsNR0CI0sHCMRCNCLDR8NMR0FkbRk0CLMND#CRCODC0FRDo
HORRRRRRRRRRRRzRd6:VRHR85N8HsI8R0E>4R42CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_M25HRR<='R4'IMECRq5)7_7)05lbNs88I0H8ER-48MFI04FR4=2RRRH2CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R ERIC5MRNs8_CNo58I8sHE80-84RF0IMF4R42RR=HC2RDR#C';j'
RRRRRRRRRRRR8CMRMoCC0sNCdRz6R;
R-RR-VRQR85N8HsI8R0E<4=R4M2RFsRIHR0CCLMNDFCRskRF00bkRNCMLRDC#CCDOD0RFOoHRCMC8
C8RRRRRRRRRRRRzRdn:VRHR85N8HsI8R0E<4=R4o2RCsMCN
0CRRRRRRRRRRRRRRRRF_k0CHM52=R<R''4;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R R;
RRRRRRRRRCRRMo8RCsMCNR0Cz;dn
RRRRR--tCCMsCN0RC0ERv)qRDOCDN#RM08Rs#H-0CN0#R
RRRRRRRRRRdRz(RR:VRFs[MRHRH5I8_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
RRRRRRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVAv)q_c.jU7XURD:RNDLCRRH#";W"
RRRRRRRRRRRRRRRRoLCHRM
RRRRRRRRRRRRRARR)_qv.UjcXRU7:qR)vnA4__1g1Rg
RRRRRRRRRRRRRRRRRsbF0NRlb7R5Q=qR>MRH_osC5[g*+8(RF0IMF*Rg[R2,q)77q>R=RIDF_8IN84s5jFR8IFM0R,j2RA7QRR=>"jjjjjjjjR",q)77A>R=RIDF_8sN84s5jFR8IFM0R,j2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRq hRR=>',4'R)11q>R=R''j, RWq>R=R0Is_5CMHR2,BqpiRR=>B,piRA hRR=>',4'R)11A>R=R''j, RWA>R=R''j,pRBi=AR>pRBi
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRR7Rmq=F>Rb,CMRA7m5R(2=F>RkL0_k5#UH*,U[2+(,mR7A25nRR=>F_k0LUk#5UH,*n[+2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mA6=2R>kRF0k_L#HU5,[U*+,62RA7m5Rc2=F>RkL0_k5#UH*,U[2+c,mR7A25dRR=>F_k0LUk#5UH,*d[+2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mA.=2R>kRF0k_L#HU5,[U*+,.2RA7m5R42=F>RkL0_k5#UH*,U[2+4,mR7A25jRR=>F_k0LUk#5UH,*,[2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRu7Qq25jRR=>HsM_Cgo5*U[+27,RQRuA=">RjR",7qmuRR=>FMbC,mR7ujA52>R=RsbNH_0$LUk#5RH,[;22
RRRRRRRRRRRRRRRR0Fk_osC5[g*2=R<R0Fk_#LkU,5HU2*[RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so*5g[2+4RR<=F_k0LUk#5UH,*4[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cgo5*.[+2=R<R0Fk_#LkU,5HU+*[.I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cog+*[d<2R=kRF0k_L#HU5,[U*+Rd2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5[g*+Rc2<F=RkL0_k5#UH*,U[2+cRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so*5g[2+6RR<=F_k0LUk#5UH,*6[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cgo5*n[+2=R<R0Fk_#LkU,5HU+*[nI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cog+*[(<2R=kRF0k_L#HU5,[U*+R(2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5[g*+RU2<b=RN0sH$k_L#HU5,R[2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRR8CMRMoCC0sNCdRz(R;
RRRRRCRRMo8RCsMCNR0Cz;dc
RRRR8CMRMoCC0sNCdRzd
;
RRRRRRRR-t-RCsMCNR0C0REC)RqvODCD#MRN8CR#D0CORoDFHVORF)sRq4vAn4_1U4_1UR
RRdRzURR:H5VROHEFOIC_HE80R4=RUo2RCsMCN
0CRRRRRRRRzRdg:FRVsRRHH5MR80CbEk_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0RC
R-RR-VRQR85N8HsI8R0E>jR42CRMC08RFsROCCN0RHIs0CCRMDNLCMRN8kRF00bkRNCMLRDC#CCDOD0RFOoH
RRRRRRRRRRRRjzcRH:RVNR58I8sHE80R4>Rjo2RCsMCN
0CRRRRRRRRRRRRRRRRF_k0CHM52=R<R''4RCIEM)R5q)77_b0l58N8s8IH04E-RI8FMR0F4Rj2=2RHR#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=WI RERCM5_N8s5CoNs88I0H8ER-48MFI04FRj=2RRRH2CCD#R''j;R
RRRRRRRRRRMRC8CRoMNCs0zCRc
j;RRRR-Q-RVNR58I8sHE80RR<=4Rj2MIFRsCH0RNCMLRDCFFsRkk0b0MRCNCLDRD#CCRO0DHFoOCRMC88C
RRRRRRRRRRRR4zcRH:RVNR58I8sHE80RR<=4Rj2oCCMsCN0
RRRRRRRRRRRRRRRR0Fk_5CMH<2R=4R''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=W
 ;RRRRRRRRRRRRCRM8oCCMsCN0R4zc;R
RR-R-RMtCC0sNCER0CqR)vCRODRD#NRM80-sH#00NCR#
RRRRRRRRRzRRc:.RRsVFRH[RMIR5HE80_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNCR
RRRRRRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqA)vj_4.4cXn:7RRLDNCHDR#WR""R;
RRRRRRRRRRRRRLRRCMoH
RRRRRRRRRRRRRRRRqA)vj_4.4cXn:7RRv)qA_4n1_4U1
4URRRRRRRRRRRRRRRRRFRbsl0RN5bR7RQq=H>RMC_soU54*4[+6FR8IFM0R*4U[R2,q)77q>R=RIDF_8IN8gs5RI8FMR0FjR2,7RQA=">Rjjjjjjjjjjjjjjjj"q,R7A7)RR=>D_FIs8N8sR5g8MFI0jFR2R,
RRRRRRRRRRRRRRRRRRRRRRRRR RRh=qR>4R''1,R1R)q='>RjR',WR q=I>RsC0_M25H,pRBi=qR>pRBi ,Rh=AR>4R''1,R1R)A='>RjR',WR A='>RjR',BApiRR=>B,piRR
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7q>R=RCFbM7,Rm4A56=2R>kRF0k_L#54nHn,4*4[+6R2,75mA4Rc2=F>RkL0_kn#454H,n+*[4,c2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7Ad542>R=R0Fk_#Lk4Hn5,*4n[d+427,Rm4A5.=2R>kRF0k_L#54nHn,4*4[+.R2,75mA4R42=F>RkL0_kn#454H,n+*[4,42RR
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7Aj542>R=R0Fk_#Lk4Hn5,*4n[j+427,RmgA52>R=R0Fk_#Lk4Hn5,*4n[2+g,mR7A25URR=>F_k0L4k#n,5H4[n*+,U2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7A25(RR=>F_k0L4k#n,5H4[n*+,(2RA7m5Rn2=F>RkL0_kn#454H,n+*[nR2,75mA6=2R>kRF0k_L#54nHn,4*6[+2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mAc=2R>kRF0k_L#54nHn,4*c[+27,RmdA52>R=R0Fk_#Lk4Hn5,*4n[2+d,mR7A25.RR=>F_k0L4k#n,5H4[n*+,.2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7A254RR=>F_k0L4k#n,5H4[n*+,42RA7m5Rj2=F>RkL0_kn#454H,n2*[,RR
RRRRRRRRRRRRRRRRRRRRRRRRR7RRQRuq=H>RMC_soU54*4[+(FR8IFM0R*4U[n+427,RQRuA=">Rj,j"
RRRRRRRRRRRRRRRRRRRRRRRRRRRRu7mq>R=RCFbM7,Rm5uA4=2R>NRbs$H0_#Lk4Hn5,*R.[2+4,mR7ujA52>R=RsbNH_0$L4k#n,5HR[.*2
2;RRRRRRRRRRRRRRRRF_k0s5Co4[U*2=R<R0Fk_#Lk4Hn5,*4n[I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+R42<F=RkL0_kn#454H,n+*[4I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+R.2<F=RkL0_kn#454H,n+*[.I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+Rd2<F=RkL0_kn#454H,n+*[dI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+Rc2<F=RkL0_kn#454H,n+*[cI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+R62<F=RkL0_kn#454H,n+*[6I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+Rn2<F=RkL0_kn#454H,n+*[nI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+R(2<F=RkL0_kn#454H,n+*[(I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+RU2<F=RkL0_kn#454H,n+*[UI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+Rg2<F=RkL0_kn#454H,n+*[gI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+24jRR<=F_k0L4k#n,5H4[n*+24jRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*4[+4<2R=kRF0k_L#54nHn,4*4[+4I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+24.RR<=F_k0L4k#n,5H4[n*+24.RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*4[+d<2R=kRF0k_L#54nHn,4*4[+dI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+24cRR<=F_k0L4k#n,5H4[n*+24cRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*4[+6<2R=kRF0k_L#54nHn,4*4[+6I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+24nRR<=bHNs0L$_kn#45.H,*R[2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[(+42=R<RsbNH_0$L4k#n,5H.+*[4I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRCRM8oCCMsCN0R.zc;R
RRRRRRMRC8CRoMNCs0zCRd
g;RRRRCRM8oCCMsCN0RUzd;R

RRRRR-RR-CRtMNCs00CRE)CRqOvRC#DDR8NMRD#CCRO0DHFoOFRVsqR)vnA4_n1d_n1d
RRRRUzdNRR:H5VROHEFOIC_HE80Rd=Rno2RCsMCN
0CRRRRRRRRzNdgRV:RFHsRRRHM5b8C0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CRRRR-Q-RVNR58I8sHE80Rg>R2CRMC08RFsROCCN0RHIs0CCRMDNLCMRN8kRF00bkRNCMLRDC#CCDOD0RFOoH
RRRRRRRRRRRRjzcNRR:H5VRNs88I0H8ERR>go2RCsMCN
0CRRRRRRRRRRRRRRRRF_k0CHM52=R<R''4RCIEM)R5q)77_b0l58N8s8IH04E-RI8FMR0Fg=2RRRH2CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R ERIC5MRNs8_CNo58I8sHE80-84RF0IMF2RgRH=R2DRC#'CRj
';RRRRRRRRRRRRCRM8oCCMsCN0RjzcNR;
R-RR-VRQR85N8HsI8R0E<g=R2FRMRHIs0CCRMDNLCsRFR0FkbRk0CLMND#CRCODC0FRDoRHOM8CCCR8
RRRRRRRRRzRRcR4N:VRHR85N8HsI8R0E<g=R2CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_M25HRR<=';4'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RW;R
RRRRRRRRRRMRC8CRoMNCs0zCRc;4N
RRRRR--tCCMsCN0RC0ERv)qRDOCDN#RM08Rs#H-0CN0#R
RRRRRRRRRRcRz.:NRRsVFRH[RMIR5HE80_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNCR
RRRRRRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqA)v4_6..Xd7RR:DCNLD#RHR""W;R
RRRRRRRRRRRRRRCRLo
HMRRRRRRRRRRRRRRRRAv)q_.64X7d.R):Rq4vAnd_1nd_1nR
RRRRRRRRRRRRRRRRRb0FsRblNRQ57q>R=R_HMs5Cod[n*+Rd48MFI0dFRn2*[,7Rq7R)q=D>RFII_Ns8858URF0IMF2Rj,RR
RRRRRRRRRRRRRRRRRRRRRRRRR7RRQ=AR>jR"jjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj,7Rq7R)A=D>RFsI_Ns8858URF0IMF2Rj,R
RRRRRRRRRRRRRRRRRRRRRRRRRRhR q>R=R''4,1R1)=qR>jR''W,R =qR>sRI0M_C5,H2RiBpq>R=RiBp,hR A>R=R''4,1R1)=AR>jR''W,R =AR>jR''B,RpRiA=B>RpRi,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRq7mRR=>FMbC,mR7A45d2>R=R0Fk_#LkdH.5,*d.[4+d27,RmdA5j=2R>kRF0k_L#5d.H.,d*d[+jR2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRA7m52.gRR=>F_k0Ldk#.,5Hd[.*+2.g,mR7AU5.2>R=R0Fk_#LkdH.5,*d.[U+.27,Rm.A5(=2R>kRF0k_L#5d.H.,d*.[+(
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRR75mA.Rn2=F>RkL0_k.#d5dH,.+*[.,n2RA7m52.6RR=>F_k0Ldk#.,5Hd[.*+2.6,mR7Ac5.2>R=R0Fk_#LkdH.5,*d.[c+.2R,
RRRRRRRRRRRRRRRRRRRRRRRRR7RRm.A5d=2R>kRF0k_L#5d.H.,d*.[+dR2,75mA.R.2=F>RkL0_k.#d5dH,.+*[.,.2RA7m52.4RR=>F_k0Ldk#.,5Hd[.*+2.4,R
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7Aj5.2>R=R0Fk_#LkdH.5,*d.[j+.27,Rm4A5g=2R>kRF0k_L#5d.H.,d*4[+gR2,75mA4RU2=F>RkL0_k.#d5dH,.+*[4,U2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRA7m524(RR=>F_k0Ldk#.,5Hd[.*+24(,mR7An542>R=R0Fk_#LkdH.5,*d.[n+427,Rm4A56=2R>kRF0k_L#5d.H.,d*4[+6
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRR75mA4Rc2=F>RkL0_k.#d5dH,.+*[4,c2RA7m524dRR=>F_k0Ldk#.,5Hd[.*+24d,mR7A.542>R=R0Fk_#LkdH.5,*d.[.+42
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mA4R42=F>RkL0_k.#d5dH,.+*[4,42RA7m524jRR=>F_k0Ldk#.,5Hd[.*+24j,mR7A25gRR=>F_k0Ldk#.,5Hd[.*+,g2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7A25URR=>F_k0Ldk#.,5Hd[.*+,U2RA7m5R(2=F>RkL0_k.#d5dH,.+*[(R2,75mAn=2R>kRF0k_L#5d.H.,d*n[+2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mA6=2R>kRF0k_L#5d.H.,d*6[+27,RmcA52>R=R0Fk_#LkdH.5,*d.[2+c,mR7A25dRR=>F_k0Ldk#.,5Hd[.*+,d2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7A25.RR=>F_k0Ldk#.,5Hd[.*+,.2RA7m5R42=F>RkL0_k.#d5dH,.+*[4R2,75mAj=2R>kRF0k_L#5d.H.,d*,[2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRQR7u=qR>MRH_osC5*dn[6+dRI8FMR0Fd[n*+2d.,QR7u=AR>jR"j"jj,mR7u=qR>bRFCRM,7Amu5Rd2=b>RN0sH$k_L#5d.H*,c[2+d,RR
RRRRRRRRRRRRRRRRRRRRRRRRR7RRm5uA.=2R>NRbs$H0_#LkdH.5,[c*+,.2Ru7mA254RR=>bHNs0L$_k.#d5cH,*4[+27,Rm5uAj=2R>NRbs$H0_#LkdH.5,[c*2
2;RRRRRRRRRRRRRRRRF_k0s5Cod[n*2=R<R0Fk_#LkdH.5,*d.[I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cod[n*+R42<F=RkL0_k.#d5dH,.+*[4I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cod[n*+R.2<F=RkL0_k.#d5dH,.+*[.I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cod[n*+Rd2<F=RkL0_k.#d5dH,.+*[dI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cod[n*+Rc2<F=RkL0_k.#d5dH,.+*[cI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cod[n*+R62<F=RkL0_k.#d5dH,.+*[6I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cod[n*+Rn2<F=RkL0_k.#d5dH,.+*[nI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cod[n*+R(2<F=RkL0_k.#d5dH,.+*[(I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cod[n*+RU2<F=RkL0_k.#d5dH,.+*[UI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cod[n*+Rg2<F=RkL0_k.#d5dH,.+*[gI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cod[n*+24jRR<=F_k0Ldk#.,5Hd[.*+24jRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_son5d*4[+4<2R=kRF0k_L#5d.H.,d*4[+4I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cod[n*+24.RR<=F_k0Ldk#.,5Hd[.*+24.RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_son5d*4[+d<2R=kRF0k_L#5d.H.,d*4[+dI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cod[n*+24cRR<=F_k0Ldk#.,5Hd[.*+24cRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_son5d*4[+6<2R=kRF0k_L#5d.H.,d*4[+6I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cod[n*+24nRR<=F_k0Ldk#.,5Hd[.*+24nRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_son5d*4[+(<2R=kRF0k_L#5d.H.,d*4[+(I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cod[n*+24URR<=F_k0Ldk#.,5Hd[.*+24URCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_son5d*4[+g<2R=kRF0k_L#5d.H.,d*4[+gI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cod[n*+2.jRR<=F_k0Ldk#.,5Hd[.*+2.jRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_son5d*.[+4<2R=kRF0k_L#5d.H.,d*.[+4I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cod[n*+2..RR<=F_k0Ldk#.,5Hd[.*+2..RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_son5d*.[+d<2R=kRF0k_L#5d.H.,d*.[+dI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cod[n*+2.cRR<=F_k0Ldk#.,5Hd[.*+2.cRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_son5d*.[+6<2R=kRF0k_L#5d.H.,d*.[+6I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cod[n*+2.nRR<=F_k0Ldk#.,5Hd[.*+2.nRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_son5d*.[+(<2R=kRF0k_L#5d.H.,d*.[+(I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cod[n*+2.URR<=F_k0Ldk#.,5Hd[.*+2.URCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_son5d*.[+g<2R=kRF0k_L#5d.H.,d*.[+gI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cod[n*+2djRR<=F_k0Ldk#.,5Hd[.*+2djRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_son5d*d[+4<2R=kRF0k_L#5d.H.,d*d[+4I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cod[n*+2d.RR<=bHNs0L$_k.#d5cH,*R[2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*dn[d+d2=R<RsbNH_0$Ldk#.,5Hc+*[4I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cod[n*+2dcRR<=bHNs0L$_k.#d5cH,*.[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cdo5n+*[dR62<b=RN0sH$k_L#5d.H*,c[2+dRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRMRC8CRoMNCs0zCRc;.N
RRRRRRRR8CMRMoCC0sNCdRzg
N;RRRRCRM8oCCMsCN0RUzdNR;
R8CMRMoCC0sNCcRzdR;
Rczc:VRHRF5M08RN8ss_CRo2oCCMsCN0RR--oCCMsCN0RD#CCRO0s
NlRRRR-Q-RV8RN8HsI8R0E<RR(NH##o'MRj0'RFMRkk8#CR0LH#R
RRjRzRRR:H5VRNs88I0H8ERR=4o2RCsMCN
0CRRRRRRRRD_FINs88RR<="jjjj"jjR#&R__N8s5Coj
2;RRRRCRM8oCCMsCN0R;zj
RRRRRz4RH:RVNR58I8sHE80R.=R2CRoMNCs0RC
RRRRRDRRFNI_8R8s<"=Rjjjjj&"RRN#_8C_soR548MFI0jFR2R;
RCRRMo8RCsMCNR0Cz
4;RRRRzR.R:VRHR85N8HsI8R0E=2RdRMoCC0sNCR
RRRRRRFRDI8_N8<sR=jR"j"jjR#&R__N8s5Co.FR8IFM0R;j2
RRRR8CMRMoCC0sNC.Rz;R
RRdRzRRR:H5VRNs88I0H8ERR=co2RCsMCN
0CRRRRRRRRD_FINs88RR<="jjj"RR&#8_N_osC58dRF0IMF2Rj;R
RRMRC8CRoMNCs0zCRdS;
z:cSRRHV58N8s8IH0=ERRR62oCCMsCN0
DSSFNI_8R8s<"=RjRj"&_R#Ns8_Cco5RI8FMR0Fj
2;S8CMRMoCC0sNCcRz;z
S6RS:H5VRNs88I0H8ERR=no2RCsMCN
0CSFSDI8_N8<sR=jR''RR&#8_N_osC586RF0IMF2Rj;R
RRMRC8CRoMNCs0zCR6R;
RzRRn:RRRRHV58N8s8IH0>ERRRn2oCCMsCN0
RRRRRRRRIDF_8N8s=R<RN#_8C_soR5n8MFI0jFR2R;
RCRRMo8RCsMCNR0Cz
n;
RRRRR--Q5VR8_HMs2CoRosCHC#0sQR7h#RkHRMoB
piRRRRzR(R:VRHRH58MC_soo2RCsMCN
0CRRRRRRRRbOsFCR##5iBp,QR7hL2RCMoH
RRRRRRRRRRRRRHV5iBpR'=R4N'RMB8RpCi'P0CM2ER0CRM
RRRRRRRRRRRRR#RR__HMsRCo<7=RQ
h;RRRRRRRRRRRRCRM8H
V;RRRRRRRRCRM8bOsFC;##
RRRR8CMRMoCC0sNC(Rz;R
RRURzRRR:H5VRMRF08_HMs2CoRMoCC0sNCR
RRRRRRRRRR_R#HsM_C<oR=QR7hR;
RCRRMo8RCsMCNR0Cz
U;
RRRRR--Q5VR80Fk_osC2CRso0H#C7sRmRzakM#HoBRmpRi
RzRRg:RRRRHV5k8F0C_soo2RCsMCN
0CRRRRRRRRbOsFCR##5pmBiF,Rks0_CRo2LHCoMR
RRRRRRRRRRVRHRB5mp=iRR''4R8NMRpmBiP'CC2M0RC0EMR
RRRRRRRRRRRRRRmR7z<aR=_R#F_k0s;Co
RRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMRFbsO#C#;R
RRMRC8CRoMNCs0zCRgR;
RzRR4RjR:VRHRF5M0FR8ks0_CRo2oCCMsCN0
RRRRRRRRRRRRz7ma=R<RF#_ks0_C
o;RRRRCRM8oCCMsCN0Rjz4;R

R-RR-VRQR85N8ss_CRo2sHCo#s0CR7q7)#RkHRMoB
piRRRRzR44RH:RVNR58_8ss2CoRMoCC0sNCR
RRRRRRsRbF#OC#BR5pRi,q)772CRLo
HMRRRRRRRRRRRRH5VRBRpi=4R''MRN8pRBiP'CC2M0RC0EMR
RRRRRRRRRRRRRR_R#Ns8_C<oR=7Rq7N)58I8sHE80-84RF0IMF2Rj;R
RRRRRRRRRRMRC8VRH;R
RRRRRRMRC8sRbF#OC#R;
RCRRMo8RCsMCNR0Cz;44
RRRR.z4RH:RVMR5FN0R8_8ss2CoRMoCC0sNCR
RRRRRRRRRR_R#Ns8_C<oR=7Rq7
);RRRRCRM8oCCMsCN0R.z4;R
RRRRRRRR
R-RR-CRtMNCs00CRE)CRqOvRC#DDR8NMRD#CCRO0DHFoOR
RR4RzdRR:VRFsHMRHRk5MlC_OD4D_.-URRR428MFI0jFRRMoCC0sNCR
RR-R-RRQV58N8s8IH0>ERRR62M8CCRR0FONsC0ICRsCH0RNCMLRDCNRM8Fbk0kC0RMDNLCCR#D0CORoDFHRO
RRRRRzRR4:cRRRHV58N8s8IH0>ERRR(2oCCMsCN0
RRRRRRRRRRRRRRRRF#_kC0_M25HRR<='R4'IMECR_5#Ns8_CNo58I8sHE80-84RF0IMF2R(RH=R2DRC#'CRj
';RRRRRRRRRRRRRRRR#s_I0M_C5RH2<W=R ERIC5MR#8_N_osC58N8s8IH04E-RI8FMR0F(=2RRRH2CCD#R''j;R
RRRRRRMRC8CRoMNCs0zCR4
c;RRRR-Q-RVNR58I8sHE80RR<=6M2RFsRIHR0CCLMNDFCRskRF00bkRNCMLRDC#CCDOD0RFOoHRCMC8
C8RRRRRRRRzR46:VRHR85N8HsI8R0E<(=R2CRoMNCs0RC
RRRRRRRRRRRRR#RR_0Fk_5CMH<2R=4R''R;
RRRRRRRRRRRRR#RR_0Is_5CMH<2R= RW;R
RRRRRRMRC8CRoMNCs0zCR4
6;RRRR-t-RCsMCNR0C0REC)RqvODCD#MRN8sR0H0-#N#0C
RRRRRRRRnz4RV:RF[sRRRHM58IH0-ERRR428MFI0jFRRMoCC0sNCR
RRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqz)vU4.RD:RNDLCRRH#"a11"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloHC5*U4.2RR&"RW"&MRH0CCosl'HN5oC[&2RR"" RH&RMo0CCHs'lCNo50oC_8CM_b8C05E5H2+4*U4.,CR8b20E2RR&"RX"&MRH0CCosl'HN5oC[2+4;R
RRRRRRRRRRCRLo
HMRRRRRRRRRRRRzv)q4R.U:)RXq.v4U1X4RR
RRRRRRRRRRRRRRFRbsl0RN5bR7>R=RH#_MC_so25[,jRqRR=>D_FINs885,j2RRq4=D>RFNI_858s4R2,q=.R>FRDI8_N8.s52R,
RRRRRRRRRRRRRRRRRRRRRRRRRRqd=D>RFNI_858sdR2,q=cR>FRDI8_N8cs52q,R6>R=RIDF_8N8s256,nRqRR=>D_FINs885,n2
SSSSRSSRRW =#>R_0Is_5CMHR2,WiBpRR=>B,piR=mR>kRF0k_L#._4U,5H[;22
RRRRRRRRRRRRRRRRF#_ks0_C[o52=R<R0Fk_#Lk_U4.5[H,2ERIC5MR#k_F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRR8CMRMoCC0sNC4RznR;
RRRRCRM8oCCMsCN0Rdz4;RRRRRRRRRRRRR
RRRRR
RRRRR--tCCMsCN0R4NRnFRIs88RCRCb)RqvODCDRRHVNsbbFHbsNR0CRRRRRRRRRRRRRRR
RzRR4:(RRRHV5lMk_DOCDc_nR4=R2CRoMNCs0RC
R-RR-VRQR85N8HsI8R0E>2R(RCMC8FR0RCOsNR0CI0sHCMRCNCLDR8NMR0FkbRk0CLMND#CRCODC0FRDo
HORRRRRRRRzN4URH:RVNR58I8sHE80R(>R2CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_Mc_nRR<='R4'IMECR#55__N8s5CoNs88I0H8ER-48MFI0(FR2RR=M_klODCD_U4.2MRN8#R5__N8s5Con=2RR''j2C2RDR#C';j'
RRRRRRRRRRRRRRRR0Is__CMn<cR= RWRCIEM5R5#8_N_osC58N8s8IH04E-RI8FMR0F(=2RRlMk_DOCD._4UN2RM58R#8_N_osC5Rn2=jR''R22CCD#R''j;R
RRRRRRMRC8CRoMNCs0zCR4;UN
RRRRRRRRUz4LRR:H5VRNs88I0H8ERR=(MRN8kRMlC_OD4D_.=URRRj2oCCMsCN0
RRRRRRRRRRRRRRRR0Fk__CMn<cR=4R''ERIC5MR5N#_8C_so25nR'=Rj2'2R#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_Mc_nRR<=WI RERCM5_5#Ns8_Cno52RR='2j'2DRC#'CRj
';RRRRRRRRCRM8oCCMsCN0RUz4LR;
R-RR-VRQR85N8HsI8R0E<6=R2FRMRHIs0CCRMDNLCsRFR0FkbRk0CLMND#CRCODC0FRDoRHOM8CCCR8
RRRRRzRR4:gRRRHV58N8s8IH0<ER=2RnRMoCC0sNCR
RRRRRRRRRRRRRRkRF0M_C_Rnc<'=R4
';RRRRRRRRRRRRRRRRI_s0CnM_c=R<R;W 
RRRRRRRR8CMRMoCC0sNC4RzgR;
R-RR-CRtMNCs00CRE)CRqOvRCRDDNRM80-sH#00NCR
SRzRRO_E	.RR:H5VR#H_I8_0ENNss$c_n5R42>2RjRMoCC0sNCR
RRRRRR.RzjRR:VRFs[MRHR_5#I0H8Es_Ns_N$n4c52RR-482RF0IMFRRjoCCMsCN0
RRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVzv)qn:cRRLDNCHDR#1R"1Ra"&MRH0CCosl'HN5oCI0H8E&2RR""7RH&RMo0CCHs'lCNo5lMk_DOCD._4U.*4U&2RR""WRH&RMo0CCHs'lCNo58IH0-ERR[.*R.-R2RR&"R "&MRH0CCosl'HN5oCo_C0C_M880CbEk5MlC_OD4D_.4U*.+URR,ncRb8C02E2R"&RX&"RR0HMCsoC'NHloIC5HE80R.-R*;[2
RRRRRRRRRRRRoLCHRM
RRRRRRRRRzRR)nqvcRR:Xv)qn.cX1RR
RRRRRRRRRRRRRbRRFRs0lRNb5R74=#>R__HMs5CoI0H8E*-.[2-4,jR7RR=>#M_H_osC58IH0.E-*.[-2q,Rj>R=RIDF_8N8s25j,4RqRR=>D_FINs885,42RRq.=D>RFNI_858s.
2,RRRRRRRRRRRRRRRRRRRRRRRRRdRqRR=>D_FINs885,d2RRqc=D>RFNI_858scR2,q=6R>FRDI8_N86s52S,
SSSSSWRR >R=R0Is__CMnRc,WiBpRR=>B,piRRm4=F>RkL0_kn#_ck5MlC_ODnD_cH,I8-0E.-*[4R2,m=jR>kRF0k_L#c_n5lMk_DOCDc_n,8IH0.E-*.[-2
2;RRRRRRRRRRRRRRRR#k_F0C_soH5I8-0E.-*[4<2R=kRF0k_L#c_n5lMk_DOCDc_n,8IH0.E-*4[-2ERIC5MRF_k0CnM_cRR='24'R#CDCZR''R;
RRRRRRRRRRRRR#RR_0Fk_osC58IH0.E-*.[-2=R<R0Fk_#Lk_5ncM_klODCD_,ncI0H8E*-.[2-.RCIEMFR5kC0_Mc_nR'=R4R'2CCD#R''Z;R
RRRRRRCRRMo8RCsMCNR0Cz;.j
RSSCRM8oCCMsCN0REzO	;_.
RSSz	OE_:4RRRHV5I#_HE80_sNsNn$_c25jRj>R2CRoMNCs0RC
RRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)RzqcvnRD:RNDLCRRH#"a11"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloMC5kOl_C_DD4*.U42.UR"&RW&"RR0HMCsoC'NHloIC5HE80R.-R*I#_HE80_sNsNn$_c254R4-R2RR&"R "&MRH0CCosl'HN5oCo_C0C_M880CbEk5MlC_OD4D_.4U*.+URR,ncRb8C02E2R"&RX&"RR0HMCsoC'NHloIC5HE80R.-R*I#_HE80_sNsNn$_c2542R;
RRRRRRRRRLRRCMoH
RRRRRRRRRRRRqz)vRnc:qR)vXnc4
1RRRRRRRRRRRRRRRRRb0FsRblNRR57=#>R__HMs5CoI0H8E*-.#H_I8_0ENNss$c_n5-424R2,q=jR>FRDI8_N8js52q,R4>R=RIDF_8N8s254,.RqRR=>D_FINs885,.2
RRRRRRRRRRRRRRRRRRRRRRRRqRRd>R=RIDF_8N8s25d,cRqRR=>D_FINs885,c2RRq6=D>RFNI_858s6
2,SSSSSRSRW= R>sRI0M_C_,ncRpWBi>R=RiBp,RRm=F>RkL0_kn#_ck5MlC_ODnD_cH,I8-0E._*#I0H8Es_Ns_N$n4c522-42R;
RRRRRRRRRRRRR#RR_0Fk_osC58IH0.E-*I#_HE80_sNsNn$_c254-R42<F=RkL0_kn#_ck5MlC_ODnD_cH,I8-0E._*#I0H8Es_Ns_N$n4c522-4RCIEMFR5kC0_Mc_nR'=R4R'2CCD#R''Z;R
RRRRRRCRRMo8RCsMCNR0Cz	OE_
4;SRRRRMRC8CRoMNCs0zCR4R(;RRRRRRRRRR

R-RR-CRtMNCs0NCRRR4nI8FsRC8CbqR)vCRODHDRVbRNbbsFs0HNCRRRRRRRRRRRRRRR
RRRR4z.RH:RVMR5kOl_C_DDd=.RRR42oCCMsCN0
RRRRR--Q5VRNs88I0H8ERR>6M2RCRC80OFRs0CNCsRIHR0CCLMNDNCRMF8Rkk0b0MRCNCLDRD#CCRO0DHFoOR
RRRRRR.Rz.:NRRRHV58N8s8IH0>ERRN(RMM8RkOl_C_DDn=cRRR42oCCMsCN0
RRRRRRRRRRRRRRRR0Fk__CMd<.R=4R''ERIC5MR5N#_8C_so85N8HsI8-0E4FR8IFM0RR(2=kRMlC_OD4D_.RU2NRM85N#_8C_so25nR'=R4R'2NRM85N#_8C_so256R'=Rj2'2R#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_M._dRR<=WI RERCM5_5#Ns8_CNo58I8sHE80-84RF0IMF2R(RM=RkOl_C_DD42.UR8NMR_5#Ns8_Cno52RR='24'R8NMR_5#Ns8_C6o52RR='2j'2DRC#'CRj
';RRRRRRRRCRM8oCCMsCN0R.z.NR;
RRRRRzRR.R.L:VRHR85N8HsI8R0E>RR(NRM8M_klODCD_Rnc/4=R2CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_M._dRR<='R4'IMECR#55__N8s5CoNs88I0H8ER-48MFI0(FR2RR=M_klODCD_U4.2MRN8#R5__N8s5Con=2RR''j2MRN8#R5__N8s5Co6=2RR''j2C2RDR#C';j'
RRRRRRRRRRRRRRRR0Is__CMd<.R= RWRCIEM5R5#8_N_osC58N8s8IH04E-RI8FMR0F(=2RRlMk_DOCD._4UN2RM58R#8_N_osC5Rn2=jR''N2RM58R#8_N_osC5R62=jR''R22CCD#R''j;R
RRRRRRMRC8CRoMNCs0zCR.;.L
RRRRRRRR.z.ORR:H5VRNs88I0H8ERR=(MRN8kRMlC_ODnD_cRR=4o2RCsMCN
0CRRRRRRRRRRRRRRRRF_k0CdM_.=R<R''4RCIEM5R5#8_N_osC5Rn2=4R''N2RM58R#8_N_osC5R62=jR''R22CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C_Rd.<W=R ERIC5MR5N#_8C_so25nR'=R4R'2NRM85N#_8C_so256R'=Rj2'2R#CDCjR''R;
RRRRRCRRMo8RCsMCNR0CzO..;R
RRRRRR.Rz.:8RRRHV58N8s8IH0=ERRNnRMM8RkOl_C_DDn/cR=2R4RMoCC0sNCR
RRRRRRRRRRRRRRkRF0M_C_Rd.<'=R4I'RERCM5_5#Ns8_CNo58I8sHE80-84RF0IMF2R6RM=RkOl_C_DDn2c2R#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_M._dRR<=WI RERCM5_5#Ns8_CNo58I8sHE80-84RF0IMF2R6RM=RkOl_C_DDn2c2R#CDCjR''R;
RRRRRCRRMo8RCsMCNR0Cz8..;R
RR-R-RRQV58N8s8IH0<ER=2R6RRMFI0sHCMRCNCLDRRFsFbk0kC0RMDNLCCR#D0CORoDFHMORCCC88R
RRRRRR.RzdRR:H5VRNs88I0H8E=R<RR62oCCMsCN0
RRRRRRRRRRRRRRRR0Fk__CMd<.R=4R''R;
RRRRRRRRRRRRRIRRsC0_M._dRR<=W
 ;RRRRRRRRCRM8oCCMsCN0Rdz.;R
RR-R-RMtCC0sNCER0CqR)vCRODNDRM08Rs#H-0CN0
RSRRORzEU	_RH:RV#R5_8IH0NE_s$sN5Rd2>2RjRMoCC0sNCS
Sz	OE_6DCRH:RVIR5HE80RR>=U_*#I0H8Es_Ns5N$dN2RMI8RHE80RR>=Uo2RCsMCN
0CRRRRRRRRRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FzVR)dqv.RR:DCNLD#RHR1"1a&"RR0HMCsoC'NHloIC5HE802RR&"R7"&MRH0CCosl'HN5oCM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*c&2RR""WRH&RMo0CCHs'lCNo58IH0-ERRLD#_8IH0RE2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50EM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*cRR+dR.,80CbER22&XR""RR&HCM0o'CsHolNCH5I8R0E-#RDLH_I8R0E+2RU;R
RRRRRRRRRRRRRRRRRRCRLo
HMSRSRR)Rzq.vdRX:R)dqv.1XU
SSSRRRRb0FsRblNRR57=b>RN#85__HMs5CoI0H8ER-48MFI0IFRHE80-LD#_8IH0,E2RRU,D_#LI0H8E2-4,jRqRR=>D_FINs885,j2
SSSSRSSRRq4=D>RFNI_858s4R2,q=.R>FRDI8_N8.s52q,Rd>R=RIDF_8N8s25d,cRqRR=>D_FINs885,c2RRW =I>RsC0_M._d,BRWp=iR>pRBiS,
SSSSSmRRRR=>0_lbU._d52j2;S
SS#SN#MHoRV:RFHsR[MRHR8IH04E-RI8FMR0FI0H8E#-DLH_I8R0EoCCMsCN0
SSSSFRRkL0_kd#_.k5MlC_ODdD_.[,H2=R<Rb0l_dU_.25j5-H[I0H8E#+DLH_I820E;R
RRRRRRRRRRRRRRRRR#k_F0C_so[5H2=R<R0Fk_#Lk_5d.M_klODCD_,d.HR[2IMECRk5F0M_C_Rd.=4R''C2RDR#C';Z'
SSSS8CMRMoCC0sNC#RN#MHo;R
RRRRRRRRRR.RzURR:VRFs[MRHRI#_HE80_sNsNd$52R-48MFI04FRRMoCC0sNCR
RRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FzVR)dqv.RR:DCNLD#RHR1"1a&"RR0HMCsoC'NHloIC5HE802RR&"R7"&MRH0CCosl'HN5oCM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*c&2RR""WRH&RMo0CCHs'lCNo58IH0-ERRLD#_8IH0-ERRU[*2RR&"R "&MRH0CCosl'HN5oCo_C0C_M880CbEk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*Rnc+.Rd,CR8b20E2RR&"RX"&MRH0CCosl'HN5oCI0H8ERR-D_#LI0H8ERR-54[-22*U;R
RRRRRRRRRRRRRLHCoMR
RRRRRRRRRRRRRzv)qd:.RRqX)vXd.U
1RRRRRRRRRRRRRRRRRb0FsRblNRR57=#>R__HMs5CoI0H8E#-DLH_I8-0EU+*[(FR8IFM0R8IH0DE-#IL_HE80-[U*2q,Rj>R=RIDF_8N8s25j,4RqRR=>D_FINs885,42RRq.=D>RFNI_858s.
2,RRRRRRRRRRRRRRRRRRRRRRRRRdRqRR=>D_FINs885,d2RRqc=D>RFNI_858scR2,W= R>sRI0M_C_,d.RpWBi>R=RiBp,RRm=0>RlUb__5d.[;22
SSSRRRRNH##o:MRRsVFRRH[H(MRRI8FMR0FjCRoMNCs0SC
SRSSR0Fk_#Lk_5d.M_klODCD_,d.I0H8E#-DLH_I8-0EU+*[HR[2<0=RlUb__5d.[H25[
2;RRRRRRRRRRRRRRRRR_R#F_k0s5CoI0H8E#-DLH_I8-0EU+*[HR[2<F=RkL0_kd#_.k5MlC_ODdD_.H,I8-0ED_#LI0H8E*-U[[+H2ERIC5MRF_k0CdM_.RR='24'R#CDCZR''R;
RRRRRRRRRRRRRCRRMo8RCsMCNR0CNH##o
M;RRRRRRRRRRRRCRM8oCCMsCN0RUz.;S
SCRM8oCCMsCN0REzO	C_D6S;
SEzO	0_o6RR:H5VRI0H8E=R>RNURMI8RHE80R8lFR>UR=2R6RMoCC0sNCR
RRRRRRRRRRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqz)vRd.:NRDLRCDH"#R1"1aRH&RMo0CCHs'lCNo58IH0RE2&7R""RR&HCM0o'CsHolNCk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*2ncR"&RW&"RR0HMCsoC'NHloIC5HE80RD-R#IL_HE802RR&"R "&MRH0CCosl'HN5oCo_C0C_M880CbEk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*Rnc+.Rd,CR8b20E2RR&"RX"&MRH0CCosl'HN5oCI0H8ERR-D_#LI0H8ERR+U
2;RRRRRRRRRRRRRRRRRRRRLHCoMS
SRRRRzv)qd:.RRqX)vXd.US1
SRSRRFRbsl0RN5bR7>R=R8bN5H#_MC_soH5I8-0E4FR8IFM0R8IH0DE-#IL_HE802U,R,#RDLH_I8-0E4R2,q=jR>FRDI8_N8js52S,
SSSSSqRR4>R=RIDF_8N8s254,.RqRR=>D_FINs885,.2RRqd=D>RFNI_858sdR2,q=cR>FRDI8_N8cs52W,R >R=R0Is__CMdR.,WiBpRR=>B,pi
SSSSRSSR=mR>lR0b__Ud#.5_8IH0NE_s$sN5-d24;22
SSSS#N#HRoM:FRVs[RHRRHMI0H8ER-48MFI0IFRHE80-LD#_8IH0oERCsMCN
0CSSSSRkRF0k_L#._d5lMk_DOCD._d,2H[RR<=0_lbU._d5I#_HE80_sNsNd$522-45-H[I0H8E#+DLH_I820E;R
RRRRRRRRRRRRRRRRR#k_F0C_so[5H2=R<R0Fk_#Lk_5d.M_klODCD_,d.HR[2IMECRk5F0M_C_Rd.=4R''C2RDR#C';Z'
SSSS8CMRMoCC0sNC#RN#MHo;R
RRRRRRRRRR.RzURR:VRFs[MRHRI#_HE80_sNsNd$52R-.8MFI0jFRRMoCC0sNCR
RRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FzVR)dqv.RR:DCNLD#RHR1"1a&"RR0HMCsoC'NHloIC5HE802RR&"R7"&MRH0CCosl'HN5oCM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*c&2RR""WRH&RMo0CCHs'lCNo5U[*2RR&"R "&MRH0CCosl'HN5oCo_C0C_M880CbEk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*Rnc+.Rd,CR8b20E2RR&"RX"&MRH0CCosl'HN5oC54[+22*U;R
RRRRRRRRRRRRRLHCoMR
RRRRRRRRRRRRRzv)qd:.RRqX)vXd.U
1RRRRRRRRRRRRRRRRRb0FsRblNRR57=#>R__HMs5CoU+*[(FR8IFM0R[U*2q,Rj>R=RIDF_8N8s25j,4RqRR=>D_FINs885,42RRq.=D>RFNI_858s.
2,RRRRRRRRRRRRRRRRRRRRRRRRRdRqRR=>D_FINs885,d2RRqc=D>RFNI_858scR2,W= R>sRI0M_C_,d.RpWBi>R=RiBp,RRm=0>RlUb__5d.[;22
SSSS#N#HRoM:FRVs[RHRRHM(FR8IFM0RojRCsMCN
0CSSSSRkRF0k_L#._d5lMk_DOCD._d,[U*+2H[RR<=0_lbU._d55[2H;[2
RRRRRRRRRRRRRRRR#RR_0Fk_osC5[U*+2H[RR<=F_k0L_k#dM.5kOl_C_DDdU.,*H[+[I2RERCM50Fk__CMd=.RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRCRM8oCCMsCN0R#N#H;oM
RRRRRRRRRRRR8CMRMoCC0sNC.RzUS;
S8CMRMoCC0sNCORzEo	_0
6;SOSzEM	_RH:RVIR5HE80RU<R2CRoMNCs0RC
RRRRRRRRRRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)Rzq.vdRD:RNDLCRRH#"a11"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloMC5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*n2RR&"RW"&MRH0CCosl'HN5oCj&2RR"" RH&RMo0CCHs'lCNo50oC_8CM_b8C0ME5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*nRd+R.8,RCEb02&2RR""XRH&RMo0CCHs'lCNo5;U2
RRRRRRRRRRRRRRRRRRRRoLCHSM
SRRRRqz)vRd.:)RXq.vdX
U1SRSSRbRRFRs0lRNb5=7R>NRb8_5#HsM_CIo5HE80-84RF0IMFHRI8-0ED_#LI0H8ER2,UD,R#IL_HE80-,42RRqj=D>RFNI_858sj
2,SSSSSRSRq=4R>FRDI8_N84s52q,R.>R=RIDF_8N8s25.,dRqRR=>D_FINs885,d2RRqc=D>RFNI_858scR2,W= R>sRI0M_C_,d.RpWBi>R=RiBp,S
SSSSSRRRm=0>RlUb__5d.j;22
SSSS#N#HRoM:FRVs[RHRRHMI0H8ER-48MFI0jFRRMoCC0sNCS
SSRSRF_k0L_k#dM.5kOl_C_DDdH.,[<2R=lR0b__Udj.52[5H2R;
RRRRRRRRRRRRRRRRRF#_ks0_CHo5[<2R=kRF0k_L#._d5lMk_DOCD._d,2H[RCIEMFR5kC0_M._dR'=R4R'2CCD#R''Z;S
SSMSC8CRoMNCs0NCR#o#HMS;
S8CMRMoCC0sNCORzEM	_;S
SCRM8oCCMsCN0REzO	;_U
zSSO_E	cRR:H5VR#H_I8_0ENNss$25.Rj>R2CRoMNCs0RC
RRRRRzRR.cc_RH:RVIR5HE80RR>=co2RCsMCN
0CRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FzVR)dqv.RR:DCNLD#RHR1"1a&"RR0HMCsoC'NHloIC5HE802RR&"R7"&MRH0CCosl'HN5oCM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*c&2RR""WRH&RMo0CCHs'lCNo5Rj2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50EM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*cRR+dR.,80CbER22&XR""RR&HCM0o'CsHolNC25c;R
RRRRRRRRRRCRLo
HMRRRRRRRRRRRRzv)qd:.RRqX)vXd.c
1RRRRRRRRRRRRRRRRRb0FsRblNRd57RR=>#M_H_osC5,d2RR7.=#>R__HMs5Co.R2,7=4R>_R#HsM_C4o527,Rj>R=RH#_MC_so25j,S
SSRRRRRRRRRRRRqRRj>R=RIDF_8N8s25j,4RqRR=>D_FINs885,42RRq.=D>RFNI_858s.
2,RRRRRRRRRRRRRRRRRRRRRRRRRdRqRR=>D_FINs885,d2RRqc=D>RFNI_858scR2,W= R>sRI0M_C_,d.RpWBi>R=RiBp,SR
SSSSSmRRd>R=R0Fk_#Lk_5d.M_klODCD_,d.dR2,m=.R>kRF0k_L#._d5lMk_DOCD._d,,.2
SSSSRSSRRm4=F>RkL0_kd#_.k5MlC_ODdD_.2,4,jRmRR=>F_k0L_k#dM.5kOl_C_DDdj.,2
2;RRRRRRRRRRRRRRRR#k_F0C_so25dRR<=F_k0L_k#dM.5kOl_C_DDdd.,2ERIC5MRF_k0CdM_.RR='24'R#CDCZR''R;
RRRRRRRRRRRRR#RR_0Fk_osC5R.2<F=RkL0_kd#_.k5MlC_ODdD_.2,.RCIEMFR5kC0_M._dR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRR_R#F_k0s5Co4<2R=kRF0k_L#._d5lMk_DOCD._d,R42IMECRk5F0M_C_Rd.=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRF#_ks0_Cjo52=R<R0Fk_#Lk_5d.M_klODCD_,d.jI2RERCM50Fk__CMd=.RR''42DRC#'CRZ
';RRRRRRRRCRM8oCCMsCN0Rcz._
c;RRRRRRRRz_.cdRR:H5VRI0H8ERR=do2RCsMCN
0CRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FzVR)dqv.RR:DCNLD#RHR1"1a&"RR0HMCsoC'NHloIC5HE802RR&"R7"&MRH0CCosl'HN5oCM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*c&2RR""WRH&RMo0CCHs'lCNo5Rj2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50EM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*cRR+dR.,80CbER22&XR""RR&HCM0o'CsHolNC25c;R
RRRRRRRRRRCRLo
HMRRRRRRRRRRRRzv)qd:.RRqX)vXd.c
1RRRRRRRRRRRRRRRRRb0FsRblNRd57RR=>',j'RR7.=#>R__HMs5Co.R2,7=4R>_R#HsM_C4o527,Rj>R=RH#_MC_so25j,S
SSRRRRRRRRRRRRqRRj>R=RIDF_8N8s25j,4RqRR=>D_FINs885,42RRq.=D>RFNI_858s.
2,RRRRRRRRRRRRRRRRRRRRRRRRRdRqRR=>D_FINs885,d2RRqc=D>RFNI_858scR2,W= R>sRI0M_C_,d.RpWBi>R=RiBp,SR
SSSSSmRRd>R=RCFbMm,R.>R=R0Fk_#Lk_5d.M_klODCD_,d..
2,SSSSSRSRm=4R>kRF0k_L#._d5lMk_DOCD._d,,42RRmj=F>RkL0_kd#_.k5MlC_ODdD_.2,j2R;
RRRRRRRRRRRRR#RR_0Fk_osC5R.2<F=RkL0_kd#_.k5MlC_ODdD_.2,.RCIEMFR5kC0_M._dR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRR_R#F_k0s5Co4<2R=kRF0k_L#._d5lMk_DOCD._d,R42IMECRk5F0M_C_Rd.=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRF#_ks0_Cjo52=R<R0Fk_#Lk_5d.M_klODCD_,d.jI2RERCM50Fk__CMd=.RR''42DRC#'CRZ
';RRRRRRRRCRM8oCCMsCN0Rcz._
d;SMSC8CRoMNCs0zCRO_E	cS;
SEzO	R_.:VRHR_5#I0H8Es_Ns5N$4>2RRRj2oCCMsCN0
RRRRRRRRcz.RV:RF[sRRRHM5I#_HE80_sNsN4$52RR-482RF0IMFRRjoCCMsCN0
RRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVzv)qd:.RRLDNCHDR#1R"1Ra"&MRH0CCosl'HN5oCI0H8E&2RR""7RH&RMo0CCHs'lCNo5lMk_DOCD._4U.*4URR+M_klODCD_*ncnRc2&WR""RR&HCM0o'CsHolNCH5I8-0EU_*#I0H8Es_Ns5N$d.2-*.[-2RR&"R "&MRH0CCosl'HN5oCo_C0C_M880CbEk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*Rnc+.Rd,CR8b20E2RR&"RX"&MRH0CCosl'HN5oCI0H8E*-U#H_I8_0ENNss$25d-[.*2R;
RRRRRRRRRLRRCMoH
RRRRRRRRRRRRqz)vRd.:qR)vXd..
1RRRRRRRRRRRRRRRRRb0FsRblNRj57RR=>#M_H_osC58IH0UE-*I#_HE80_sNsNd$52*-.[2-.,4R7RR=>#M_H_osC58IH0UE-*I#_HE80_sNsNd$52*-.[2-4,jRqRR=>D_FINs885,j2RRq4=D>RFNI_858s4R2,q=.R>FRDI8_N8.s52R,
RRRRRRRRRRRRRRRRRRRRRRRRRRqd=D>RFNI_858sdR2,q=cR>FRDI8_N8cs52W,R >R=R0Is__CMdR.,WiBpRR=>B,piRRmj=F>RkL0_kd#_.k5MlC_ODdD_.H,I8-0EU_*#I0H8Es_Ns5N$d.2-*.[-2S,
SSSSSmRR4>R=R0Fk_#Lk_5d.M_klODCD_,d.I0H8E*-U#H_I8_0ENNss$25d-[.*-242;R
RRRRRRRRRRRRRR_R#F_k0s5CoI0H8E*-U#H_I8_0ENNss$25d-[.*-R42<F=RkL0_kd#_.k5MlC_ODdD_.H,I8-0EU_*#I0H8Es_Ns5N$d.2-*4[-2ERIC5MRF_k0CdM_.RR='24'R#CDCZR''R;
RRRRRRRRRRRRR#RR_0Fk_osC58IH0UE-*I#_HE80_sNsNd$52*-.[2-.RR<=F_k0L_k#dM.5kOl_C_DDdI.,HE80-#U*_8IH0NE_s$sN5-d2.-*[.I2RERCM50Fk__CMd=.RR''42DRC#'CRZ
';RRRRRRRRCRM8oCCMsCN0Rcz.;S
SCRM8oCCMsCN0REzO	;_.
zSSO_E	4RR:H5VR#H_I8_0ENNss$25jRj>R2CRoMNCs0RC
RRRRRzRR.:cRRRHV58IH0lERFU8RR4=R2CRoMNCs0RC
RRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)Rzq.vdRD:RNDLCRRH#"a11"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloMC5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*n2RR&"RW"&MRH0CCosl'HN5oCj&2RR"" RH&RMo0CCHs'lCNo50oC_8CM_b8C0ME5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*nRd+R.8,RCEb02&2RR""XRH&RMo0CCHs'lCNo5;42
RRRRRRRRRRRRoLCHRM
RRRRRRRRRzRR)dqv.RR:)dqv.1X4RR
RRRRRRRRRRRRRRFRbsl0RN5bR7>R=RH#_MC_so25j,jRqRR=>D_FINs885,j2RRq4=D>RFNI_858s4R2,q=.R>FRDI8_N8.s52R,
RRRRRRRRRRRRRRRRRRRRRRRRRRqd=D>RFNI_858sdR2,q=cR>FRDI8_N8cs52W,R >R=R0Is__CMdR.,WiBpRR=>B,piR=mR>kRF0k_L#._d5lMk_DOCD._d,2j2;R
RRRRRRRRRRRRRR_R#F_k0s5Coj<2R=kRF0k_L#._d5lMk_DOCD._d,Rj2IMECRk5F0M_C_Rd.=4R''C2RDR#C';Z'
RRRRRRRR8CMRMoCC0sNC.RzcS;
S8CMRMoCC0sNCORzE4	_;R
RRMRC8CRoMNCs0zCR.R4;RRRRRRRRRR

R-RR-CRtMNCs0NCRRR4nI8FsRC8CbqR)vCRODHDRVbRNbbsFs0HNCRRRRRRRRRRRRRRR
RRRR6z.RH:RVMR5kOl_C_DD4=nRRR42oCCMsCN0
RRRRR--Q5VRNs88I0H8ERR>6M2RCRC80OFRs0CNCsRIHR0CCLMNDNCRMF8Rkk0b0MRCNCLDRD#CCRO0DHFoOR
RRRRRR.Rzn:NRRRHV58N8s8IH0>ERRN(RMM8RkOl_C_DDn=cRRN4RMM8RkOl_C_DDd=.RRR42oCCMsCN0
RRRRRRRRRRRRRRRR0Fk__CM4<nR=4R''ERIC5MR5N#_8C_so85N8HsI8-0E4FR8IFM0RR(2=kRMlC_OD4D_.RU2NRM85N#_8C_so25nR'=R4R'2NRM85N#_8C_so256R'=R4R'2NRM85N#_8C_so25cR'=Rj2'2R#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_Mn_4RR<=WI RERCM5_5#Ns8_CNo58I8sHE80-84RF0IMF2R(RM=RkOl_C_DD42.UR8NMR_5#Ns8_Cno52RR='24'R8NMR_5#Ns8_C6o52RR='24'R8NMR_5#Ns8_Cco52RR='2j'2DRC#'CRj
';RRRRRRRRCRM8oCCMsCN0Rnz.NR;
RRRRRzRR.RnL:VRHR85N8HsI8R0E>RR(NRM8M_klODCD_Rnc=RR4NRM8M_klODCD_Rd.=2RjRMoCC0sNCR
RRRRRRRRRRRRRRkRF0M_C_R4n<'=R4I'RERCM5_5#Ns8_CNo58I8sHE80-84RF0IMF2R(RM=RkOl_C_DD42.UR8NMR_5#Ns8_Cno52RR='24'R8NMR_5#Ns8_C6o52RR='2j'R8NMR_5#Ns8_Cco52RR='2j'2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0C4M_n=R<RRW IMECR#55__N8s5CoNs88I0H8ER-48MFI0(FR2RR=M_klODCD_U4.2MRN8#R5__N8s5Con=2RR''42MRN8#R5__N8s5Co6=2RR''j2MRN8#R5__N8s5Coc=2RR''j2C2RDR#C';j'
RRRRRRRR8CMRMoCC0sNC.Rzn
L;RRRRRRRRzO.nRH:RVNR58I8sHE80R(>RR8NMRlMk_DOCDc_nRj=RR8NMRlMk_DOCD._dR4=R2CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_Mn_4RR<='R4'IMECR#55__N8s5CoNs88I0H8ER-48MFI0(FR2RR=M_klODCD_U4.2MRN8#R5__N8s5Con=2RR''j2MRN8#R5__N8s5Co6=2RR''42MRN8#R5__N8s5Coc=2RR''j2C2RDR#C';j'
RRRRRRRRRRRRRRRR0Is__CM4<nR= RWRCIEM5R5#8_N_osC58N8s8IH04E-RI8FMR0F(=2RRlMk_DOCD._4UN2RM58R#8_N_osC5Rn2=jR''N2RM58R#8_N_osC5R62=4R''N2RM58R#8_N_osC5Rc2=jR''R22CCD#R''j;R
RRRRRRMRC8CRoMNCs0zCR.;nO
RRRRRRRRnz.8RR:H5VRNs88I0H8ERR>(MRN8kRMlC_ODnD_cRR=jMRN8kRMlC_ODdD_.RR=jo2RCsMCN
0CRRRRRRRRRRRRRRRRF_k0C4M_n=R<R''4RCIEM5R5#8_N_osC58N8s8IH04E-RI8FMR0F(=2RRlMk_DOCD._4UN2RM58R#8_N_osC5Rn2=jR''N2RM58R#8_N_osC5R62=jR''N2RM58R#8_N_osC5Rc2=jR''R22CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C_R4n<W=R ERIC5MR5N#_8C_so85N8HsI8-0E4FR8IFM0RR(2=kRMlC_OD4D_.RU2NRM85N#_8C_so25nR'=RjR'2NRM85N#_8C_so256R'=RjR'2NRM85N#_8C_so25cR'=Rj2'2R#CDCjR''R;
RRRRRCRRMo8RCsMCNR0Cz8.n;R
RRRRRR.Rzn:CRRRHV58N8s8IH0=ERRN(RMM8RkOl_C_DDn=cRRN4RMM8RkOl_C_DDd=.RRR42oCCMsCN0
RRRRRRRRRRRRRRRR0Fk__CM4<nR=4R''ERIC5MR5N#_8C_so25nR'=R4R'2NRM85N#_8C_so256R'=R4R'2NRM85N#_8C_so25cR'=Rj2'2R#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_Mn_4RR<=WI RERCM5_5#Ns8_Cno52RR='24'R8NMR_5#Ns8_C6o52RR='24'R8NMR#R5__N8s5Coc=2RR''j2C2RDR#C';j'
RRRRRRRR8CMRMoCC0sNC.Rzn
C;RRRRRRRRzV.nRH:RVNR58I8sHE80R(=RR8NMRlMk_DOCDc_nR4=RR8NMRlMk_DOCD._dRj=R2CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_Mn_4RR<='R4'IMECR#55__N8s5Con=2RR''42MRN8#R5__N8s5Co6=2RR''j2MRN8#R5__N8s5Coc=2RR''j2C2RDR#C';j'
RRRRRRRRRRRRRRRR0Is__CM4<nR= RWRCIEM5R5#8_N_osC5Rn2=4R''N2RM58R#8_N_osC5R62=jR''N2RM58R#8_N_osC5Rc2=jR''R22CCD#R''j;R
RRRRRRMRC8CRoMNCs0zCR.;nV
RRRRRRRRnz.oRR:H5VRNs88I0H8ERR=nMRN8kRMlC_ODnD_cRR=jMRN8kRMlC_ODdD_.RR=4o2RCsMCN
0CRRRRRRRRRRRRRRRRF_k0C4M_n=R<R''4RCIEM5R5#8_N_osC5R62=4R''N2RM58R#8_N_osC5Rc2=jR''R22CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C_R4n<W=R ERIC5MR5N#_8C_so256R'=R4R'2NRM85N#_8C_so25cR'=Rj2'2R#CDCjR''R;
RRRRRCRRMo8RCsMCNR0Czo.n;R
RRRRRR.Rzn:ERRRHV58N8s8IH0=ERRN6RMM8RkOl_C_DDd/.R=2R4RMoCC0sNCR
RRRRRRRRRRRRRRkRF0M_C_R4n<'=R4I'RERCM5_5#Ns8_CNo58I8sHE80-84RF0IMF2RcRM=RkOl_C_DDd2.2R#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_Mn_4RR<=WI RERCM5_5#Ns8_CNo58I8sHE80-84RF0IMF2RcRM=RkOl_C_DDd2.2R#CDCjR''R;
RRRRRCRRMo8RCsMCNR0CzE.n;R
RR-R-RRQV58N8s8IH0<ER=2R6RRMFI0sHCMRCNCLDRRFsFbk0kC0RMDNLCCR#D0CORoDFHMORCCC88R
RRRRRR.Rz(RR:H5VRNs88I0H8E=R<RRc2oCCMsCN0
RRRRRRRRRRRRRRRR0Fk__CM4<nR=4R''R;
RRRRRRRRRRRRRIRRsC0_Mn_4RR<=W
 ;RRRRRRRRCRM8oCCMsCN0R(z.;R
RR-R-RMtCC0sNCER0CqR)vCRODNDRM08Rs#H-0CN0
RSRRORzEU	_RH:RV#R5_8IH0NE_s$sN5Rd2>2RjRMoCC0sNCS
Sz	OE_6DCRH:RVIR5HE80RR>=U_*#I0H8Es_Ns5N$dN2RMI8RHE80RR>=Uo2RCsMCN
0CRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FzVR)4qvnRR:DCNLD#RHR1"1a&"RR0HMCsoC'NHloIC5HE802RR&"R7"&MRH0CCosl'HN5oCM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*cRR+M_klODCD_*d.dR.2&WR""RR&HCM0o'CsHolNCH5I8R0E-#RDLH_I820ER"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05lMk_DOCD._4U.*4URR+M_klODCD_*ncn+cRRlMk_DOCD._d*Rd.+nR4,CR8b20E2RR&"RX"&MRH0CCosl'HN5oCI0H8ERR-D_#LI0H8ERR+U
2;RRRRRRRRRRRRLHCoMS
SRRRRzv)q4:nRRqX)vX4nUS1
SRSRRFRbsl0RN5bR7>R=R8bN5H#_MC_soH5I8-0E4FR8IFM0R8IH0DE-#IL_HE802U,R,#RDLH_I8-0E4R2,q=jR>FRDI8_N8js52S,
SSSSSqRR4>R=RIDF_8N8s254,.RqRR=>D_FINs885,.2RRqd=D>RFNI_858sdR2,W= R>sRI0M_C_,4nRpWBi>R=RiBp,S
SSSSSRRRm=0>RlUb__54nj;22
SSSS#N#HRoM:FRVs[RHRRHMI0H8ER-48MFI0IFRHE80-LD#_8IH0oERCsMCN
0CSSSSRkRF0k_L#n_45lMk_DOCDn_4,2H[RR<=0_lbUn_455j2HI[-HE80+LD#_8IH0;E2
RRRRRRRRRRRRRRRR#RR_0Fk_osC52H[RR<=F_k0L_k#4Mn5kOl_C_DD4Hn,[I2RERCM50Fk__CM4=nRR''42DRC#'CRZ
';SSSSCRM8oCCMsCN0R#N#H;oM
RRRRRRRRRRRRUz.RV:RF[sRRRHM#H_I8_0ENNss$25d-84RF0IMFRR4oCCMsCN0
RRRRRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)Rzqnv4RD:RNDLCRRH#"a11"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloMC5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*nRM+RkOl_C_DDdd.*.&2RR""WRH&RMo0CCHs'lCNo58IH0-ERRLD#_8IH0-ERRU[*2RR&"R "&MRH0CCosl'HN5oCo_C0C_M880CbEk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*Rnc+kRMlC_ODdD_..*dR4+Rn8,RCEb02&2RR""XRH&RMo0CCHs'lCNo58IH0-ERRLD#_8IH0-ERR-5[4U2*2R;
RRRRRRRRRRRRRoLCHRM
RRRRRRRRRRRRRqz)vR4n:)RXqnv4XRU1
RRRRRRRRRRRRRRRRsbF0NRlb7R5RR=>#M_H_osC58IH0DE-#IL_HE80-[U*+8(RF0IMFHRI8-0ED_#LI0H8E*-U[R2,q=jR>FRDI8_N8js52q,R4>R=RIDF_8N8s254,.RqRR=>D_FINs885,.2
RRRRRRRRRRRRRRRRRRRRRRRRqRRd>R=RIDF_8N8s25d, RWRR=>I_s0C4M_nW,RBRpi=B>RpRi,m>R=Rb0l_4U_n25[2S;
SRSRR#RN#MHoRV:RFHsR[MRHR8(RF0IMFRRjoCCMsCN0
SSSSFRRkL0_k4#_nk5MlC_OD4D_nH,I8-0ED_#LI0H8E*-U[[+H2=R<Rb0l_4U_n25[52H[;R
RRRRRRRRRRRRRRRRR#k_F0C_soH5I8-0ED_#LI0H8E*-U[[+H2=R<R0Fk_#Lk_54nM_klODCD_,4nI0H8E#-DLH_I8-0EU+*[HR[2IMECRk5F0M_C_R4n=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR8CMRMoCC0sNC#RN#MHo;R
RRRRRRRRRRMRC8CRoMNCs0zCR.
U;SMSC8CRoMNCs0zCRO_E	D;C6
zSSO_E	oR06:VRHRH5I8R0E>U=RR8NMR8IH0lERFU8RRR>=6o2RCsMCN
0CRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FzVR)4qvnRR:DCNLD#RHR1"1a&"RR0HMCsoC'NHloIC5HE802RR&"R7"&MRH0CCosl'HN5oCM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*cRR+M_klODCD_*d.dR.2&WR""RR&HCM0o'CsHolNCH5I8R0E-#RDLH_I820ER"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05lMk_DOCD._4U.*4URR+M_klODCD_*ncn+cRRlMk_DOCD._d*Rd.+nR4,CR8b20E2RR&"RX"&MRH0CCosl'HN5oCI0H8ERR-D_#LI0H8ERR+U
2;RRRRRRRRRRRRLHCoMS
SRRRRzv)q4:nRRqX)vX4nUS1
SRSRRFRbsl0RN5bR7>R=R8bN5H#_MC_soH5I8-0E4FR8IFM0R8IH0DE-#IL_HE802U,R,#RDLH_I8-0E4R2,q=jR>FRDI8_N8js52S,
SSSSSqRR4>R=RIDF_8N8s254,.RqRR=>D_FINs885,.2RRqd=D>RFNI_858sdR2,W= R>sRI0M_C_,4nRpWBi>R=RiBp,S
SSSSSRRRm=0>RlUb__54n#H_I8_0ENNss$25d-242;S
SS#SN#MHoRV:RFHsR[MRHR8IH04E-RI8FMR0FI0H8E#-DLH_I8R0EoCCMsCN0
SSSSFRRkL0_k4#_nk5MlC_OD4D_n[,H2=R<Rb0l_4U_n_5#I0H8Es_Ns5N$d42-2[5H-8IH0DE+#IL_HE802R;
RRRRRRRRRRRRRRRRRF#_ks0_CHo5[<2R=kRF0k_L#n_45lMk_DOCDn_4,2H[RCIEMFR5kC0_Mn_4R'=R4R'2CCD#R''Z;S
SSMSC8CRoMNCs0NCR#o#HMR;
RRRRRRRRRzRR.:URRsVFRH[RM_R#I0H8Es_Ns5N$d.2-RI8FMR0FjCRoMNCs0RC
RRRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVzv)q4:nRRLDNCHDR#1R"1Ra"&MRH0CCosl'HN5oCI0H8E&2RR""7RH&RMo0CCHs'lCNo5lMk_DOCD._4U.*4URR+M_klODCD_*ncn+cRRlMk_DOCD._d*2d.R"&RW&"RR0HMCsoC'NHlo[C5*RU2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50EM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*cRR+M_klODCD_*d.d+.RR,4nRb8C02E2R"&RX&"RR0HMCsoC'NHlo5C5[2+4*;U2
RRRRRRRRRRRRLRRCMoH
RRRRRRRRRRRRzRR)4qvnRR:Xv)q4UnX1RR
RRRRRRRRRRRRRbRRFRs0lRNb5=7R>_R#HsM_CUo5*([+RI8FMR0FU2*[,jRqRR=>D_FINs885,j2RRq4=D>RFNI_858s4R2,q=.R>FRDI8_N8.s52R,
RRRRRRRRRRRRRRRRRRRRRRRRRRqd=D>RFNI_858sdR2,W= R>sRI0M_C_,4nRpWBi>R=RiBp,RRm=0>RlUb__54n[;22
SSSS#N#HRoM:FRVs[RHRRHM(FR8IFM0RojRCsMCN
0CSSSSRkRF0k_L#n_45lMk_DOCDn_4,[U*+2H[RR<=0_lbUn_455[2H;[2
RRRRRRRRRRRRRRRR#RR_0Fk_osC5[U*+2H[RR<=F_k0L_k#4Mn5kOl_C_DD4Un,*H[+[I2RERCM50Fk__CM4=nRR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRCRM8oCCMsCN0R#N#H;oM
RRRRRRRRRRRR8CMRMoCC0sNC.RzUS;
S8CMRMoCC0sNCORzEo	_0
6;SOSzEM	_RH:RVIR5HE80RU<R2CRoMNCs0RC
RRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)Rzqnv4RD:RNDLCRRH#"a11"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloMC5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*nRM+RkOl_C_DDdd.*.&2RR""WRH&RMo0CCHs'lCNo5Rj2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50EM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*cRR+M_klODCD_*d.d+.RR,4nRb8C02E2R"&RX&"RR0HMCsoC'NHloUC52R;
RRRRRRRRRLRRCMoH
RSSRzRR)4qvnRR:Xv)q4UnX1S
SSRRRRsbF0NRlb7R5RR=>b5N8#M_H_osC58IH04E-RI8FMR0FI0H8E#-DLH_I820E,,RURLD#_8IH04E-2q,Rj>R=RIDF_8N8s25j,S
SSSSSR4RqRR=>D_FINs885,42RRq.=D>RFNI_858s.R2,q=dR>FRDI8_N8ds52W,R >R=R0Is__CM4Rn,WiBpRR=>B,pi
SSSSRSSR=mR>lR0b__U4jn52
2;SSSSNH##o:MRRsVFRRH[HIMRHE80-84RF0IMFRRjoCCMsCN0
SSSSFRRkL0_k4#_nk5MlC_OD4D_n[,H2=R<Rb0l_4U_n25j52H[;R
RRRRRRRRRRRRRRRRR#k_F0C_so[5H2=R<R0Fk_#Lk_54nM_klODCD_,4nHR[2IMECRk5F0M_C_R4n=4R''C2RDR#C';Z'
SSSS8CMRMoCC0sNC#RN#MHo;S
SCRM8oCCMsCN0REzO	;_M
CSSMo8RCsMCNR0Cz	OE_
U;SOSzEc	_RH:RV#R5_8IH0NE_s$sN5R.2>2RjRMoCC0sNCR
RRRRRR.RzgR_c:VRHRH5I8R0E>c=R2CRoMNCs0RC
RRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)Rzqnv4RD:RNDLCRRH#"a11"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloMC5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*nRM+RkOl_C_DDdd.*.&2RR""WRH&RMo0CCHs'lCNo5Rj2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50EM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*cRR+M_klODCD_*d.d+.RR,4nRb8C02E2R"&RX&"RR0HMCsoC'NHlocC52R;
RRRRRRRRRLRRCMoH
RRRRRRRRRRRRqz)vR4n:qR)vX4nc
1RRRRRRRRRRRRRRRRRb0FsRblNRd57RR=>#M_H_osC5,d2RR7.=#>R__HMs5Co.R2,7=4R>_R#HsM_C4o527,Rj>R=RH#_MC_so25j,S
SSRRRRRRRRRRRRqRRj>R=RIDF_8N8s25j,4RqRR=>D_FINs885,42RRq.=D>RFNI_858s.
2,RRRRRRRRRRRRRRRRRRRRRRRRRdRqRR=>D_FINs885,d2RRW =I>RsC0_Mn_4,BRWp=iR>pRBi
,RSSSSSRSRm=dR>kRF0k_L#n_45lMk_DOCDn_4,,d2RRm.=F>RkL0_k4#_nk5MlC_OD4D_n2,.,S
SSSSSR4RmRR=>F_k0L_k#4Mn5kOl_C_DD44n,2m,Rj>R=R0Fk_#Lk_54nM_klODCD_,4nj;22
RRRRRRRRRRRRRRRRF#_ks0_Cdo52=R<R0Fk_#Lk_54nM_klODCD_,4ndI2RERCM50Fk__CM4=nRR''42DRC#'CRZ
';RRRRRRRRRRRRRRRR#k_F0C_so25.RR<=F_k0L_k#4Mn5kOl_C_DD4.n,2ERIC5MRF_k0C4M_nRR='24'R#CDCZR''R;
RRRRRRRRRRRRR#RR_0Fk_osC5R42<F=RkL0_k4#_nk5MlC_OD4D_n2,4RCIEMFR5kC0_Mn_4R'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRR_R#F_k0s5Coj<2R=kRF0k_L#n_45lMk_DOCDn_4,Rj2IMECRk5F0M_C_R4n=4R''C2RDR#C';Z'
RRRRRRRR8CMRMoCC0sNC.Rzg;_c
RRRRRRRRgz._:dRRRHV58IH0=ERRRd2oCCMsCN0
RRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVzv)q4:nRRLDNCHDR#1R"1Ra"&MRH0CCosl'HN5oCI0H8E&2RR""7RH&RMo0CCHs'lCNo5lMk_DOCD._4U.*4URR+M_klODCD_*ncn+cRRlMk_DOCD._d*2d.R"&RW&"RR0HMCsoC'NHlojC52RR&"R "&MRH0CCosl'HN5oCo_C0C_M880CbEk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*Rnc+kRMlC_ODdD_..*dR4+Rn8,RCEb02&2RR""XRH&RMo0CCHs'lCNo5;c2
RRRRRRRRRRRRoLCHRM
RRRRRRRRRzRR)4qvnRR:)4qvn1XcRR
RRRRRRRRRRRRRRFRbsl0RN5bR7=dR>jR''7,R.>R=RH#_MC_so25.,4R7RR=>#M_H_osC5,42RR7j=#>R__HMs5Coj
2,SRSSRRRRRRRRRRRRRRqj=D>RFNI_858sjR2,q=4R>FRDI8_N84s52q,R.>R=RIDF_8N8s25.,R
RRRRRRRRRRRRRRRRRRRRRRRRRq=dR>FRDI8_N8ds52W,R >R=R0Is__CM4Rn,WiBpRR=>B,piRS
SSSSSRdRmRR=>FMbC,.RmRR=>F_k0L_k#4Mn5kOl_C_DD4.n,2S,
SSSSSmRR4>R=R0Fk_#Lk_54nM_klODCD_,4n4R2,m=jR>kRF0k_L#n_45lMk_DOCDn_4,2j2;R
RRRRRRRRRRRRRR_R#F_k0s5Co.<2R=kRF0k_L#n_45lMk_DOCDn_4,R.2IMECRk5F0M_C_R4n=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRF#_ks0_C4o52=R<R0Fk_#Lk_54nM_klODCD_,4n4I2RERCM50Fk__CM4=nRR''42DRC#'CRZ
';RRRRRRRRRRRRRRRR#k_F0C_so25jRR<=F_k0L_k#4Mn5kOl_C_DD4jn,2ERIC5MRF_k0C4M_nRR='24'R#CDCZR''R;
RRRRRCRRMo8RCsMCNR0Cz_.gdS;
S8CMRMoCC0sNCORzEc	_;S
Sz	OE_:.RRRHV5I#_HE80_sNsN4$52RR>jo2RCsMCN
0CRRRRRRRRzRdj:FRVsRR[H5MR#H_I8_0ENNss$254R4-R2FR8IFM0RojRCsMCN
0CRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FzVR)4qvnRR:DCNLD#RHR1"1a&"RR0HMCsoC'NHloIC5HE802RR&"R7"&MRH0CCosl'HN5oCM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*cRR+M_klODCD_*d.dR.2&WR""RR&HCM0o'CsHolNCH5I8-0EU_*#I0H8Es_Ns5N$d.2-*.[-2RR&"R "&MRH0CCosl'HN5oCo_C0C_M880CbEk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*Rnc+kRMlC_ODdD_..*dR4+Rn8,RCEb02&2RR""XRH&RMo0CCHs'lCNo58IH0UE-*I#_HE80_sNsNd$52*-.[
2;RRRRRRRRRRRRLHCoMR
RRRRRRRRRR)Rzqnv4R):Rqnv4XR.1
RRRRRRRRRRRRRRRRsbF0NRlb7R5j>R=RH#_MC_soH5I8-0EU_*#I0H8Es_Ns5N$d.2-*.[-27,R4>R=RH#_MC_soH5I8-0EU_*#I0H8Es_Ns5N$d.2-*4[-2q,Rj>R=RIDF_8N8s25j,4RqRR=>D_FINs885,42RRq.=D>RFNI_858s.
2,RRRRRRRRRRRRRRRRRRRRRRRRRdRqRR=>D_FINs885,d2RRW =I>RsC0_Mn_4,BRWp=iR>pRBim,Rj>R=R0Fk_#Lk_54nM_klODCD_,4nI0H8E*-U#H_I8_0ENNss$25d-[.*-,.2
SSSSRSSRRm4=F>RkL0_k4#_nk5MlC_OD4D_nH,I8-0EU_*#I0H8Es_Ns5N$d.2-*4[-2
2;RRRRRRRRRRRRRRRR#k_F0C_soH5I8-0EU_*#I0H8Es_Ns5N$d.2-*4[-2=R<R0Fk_#Lk_54nM_klODCD_,4nI0H8E*-U#H_I8_0ENNss$25d-[.*-R42IMECRk5F0M_C_R4n=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRF#_ks0_CIo5HE80-#U*_8IH0NE_s$sN5-d2.-*[.<2R=kRF0k_L#n_45lMk_DOCDn_4,8IH0UE-*I#_HE80_sNsNd$52*-.[2-.RCIEMFR5kC0_Mn_4R'=R4R'2CCD#R''Z;R
RRRRRRMRC8CRoMNCs0zCRd
j;SMSC8CRoMNCs0zCRO_E	.S;
SEzO	R_4:VRHR_5#I0H8Es_Ns5N$j>2RRRj2oCCMsCN0
RRRRRRRR4zdRH:RVIR5HE80R8lFR=URRR42oCCMsCN0
RRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVzv)q4:nRRLDNCHDR#1R"1Ra"&MRH0CCosl'HN5oCI0H8E&2RR""7RH&RMo0CCHs'lCNo5lMk_DOCD._4U.*4URR+M_klODCD_*ncn+cRRlMk_DOCD._d*2d.R"&RW&"RR0HMCsoC'NHlojC52RR&"R "&MRH0CCosl'HN5oCo_C0C_M880CbEk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*Rnc+kRMlC_ODdD_..*dR4+Rn8,RCEb02&2RR""XRH&RMo0CCHs'lCNo5;42
RRRRRRRRRRRRoLCHRM
RRRRRRRRRzRR)4qvnRR:)4qvn1X4RR
RRRRRRRRRRRRRRFRbsl0RN5bR7>R=RH#_MC_so25j,jRqRR=>D_FINs885,j2RRq4=D>RFNI_858s4R2,q=.R>FRDI8_N8.s52R,
RRRRRRRRRRRRRRRRRRRRRRRRRRqd=D>RFNI_858sdR2,W= R>sRI0M_C_,4nRpWBi>R=RiBp,RRm=F>RkL0_k4#_nk5MlC_OD4D_n2,j2R;
RRRRRRRRRRRRR#RR_0Fk_osC5Rj2<F=RkL0_k4#_nk5MlC_OD4D_n2,jRCIEMFR5kC0_Mn_4R'=R4R'2CCD#R''Z;R
RRRRRRMRC8CRoMNCs0zCRd
4;SMSC8CRoMNCs0zCRO_E	4R;
RRRRCRM8oCCMsCN0R6z.;RRRRRRRR
RRRCRRMo8RCsMCNR0Cz;cc
8CMRONsECH0Os0kCDRLF_O	s;Nl
s
NO0EHCkO0sMCRFI_s_COEOF	RVqR)vW_)R
H#ObFlFMMC0)RXq.v4U1X4
FRbs50R
RRRmRR:FRk0#_08DHFoOR;
RjRqRH:RM0R#8F_Do;HO
RRRq:4RRRHM#_08DHFoOR;
R.RqRH:RM0R#8F_Do;HO
RRRq:dRRRHM#_08DHFoOR;
RcRqRH:RM0R#8F_Do;HO
RRRq:6RRRHM#_08DHFoOR;
RnRqRH:RM0R#8F_Do;HO
RRR7RR:H#MR0D8_FOoH;R
RRpWBiRR:H#MR0D8_FOoH;R
RRRW :MRHR8#0_oDFHRO
2C;
MO8RFFlbM0CM;


ObFlFMMC0)RXqcvnX
.1RsbF0
R5RmRRjRR:FRk0#_08DHFoOR;
R4RmRF:Rk#0R0D8_FOoH;R
RRRqj:MRHR8#0_oDFH
O;RqRR4RR:H#MR0D8_FOoH;R
RRRq.:MRHR8#0_oDFH
O;RqRRdRR:H#MR0D8_FOoH;R
RRRqc:MRHR8#0_oDFH
O;RqRR6RR:H#MR0D8_FOoH;R
RRR7j:MRHR8#0_oDFH
O;R7RR4RR:H#MR0D8_FOoH;R
RRpWBiRR:H#MR0D8_FOoH;R
RRRW :MRHR8#0_oDFHRO
2C;
MO8RFFlbM0CM;O

FFlbM0CMRqX)vXd.cR1
b0FsRR5
RjRmRF:Rk#0R0D8_FOoH;R
RRRm4:kRF00R#8F_Do;HO
RRRm:.RR0FkR8#0_oDFH
O;RmRRdRR:FRk0#_08DHFoOR;
RjRqRH:RM0R#8F_Do;HO
RRRq:4RRRHM#_08DHFoOR;
R.RqRH:RM0R#8F_Do;HO
RRRq:dRRRHM#_08DHFoOR;
RcRqRH:RM0R#8F_Do;HO
RRR7:jRRRHM#_08DHFoOR;
R4R7RH:RM0R#8F_Do;HO
RRR7:.RRRHM#_08DHFoOR;
RdR7RH:RM0R#8F_Do;HO
RRRWiBpRH:RM0R#8F_Do;HO
RRRW: RRRHM#_08DHFoO2
R;M
C8FROlMbFC;M0
lOFbCFMMX0R)dqv.1XU
b
RFRs05R
RR:mRR0FkR8#0_oDFHPO_CFO0sR5(8MFI0jFR2R;
RjRqRH:RM0R#8F_Do;HO
RRRq:4RRRHM#_08DHFoOR;
R.RqRH:RM0R#8F_Do;HO
RRRq:dRRRHM#_08DHFoOR;
RcRqRH:RM0R#8F_Do;HO
RRR7RR:H#MR0D8_FOoH_OPC05Fs(FR8IFM0R;j2
RRRWiBpRH:RM0R#8F_Do;HO
RRRW: RRRHM#_08DHFoO2
R;M
C8FROlMbFC;M0
F
OlMbFCRM0Xv)q4UnX1b
RFRs05R
RR:mRR0FkR8#0_oDFHPO_CFO0sR5(8MFI0jFR2R;
RjRqRH:RM0R#8F_Do;HO
RRRq:4RRRHM#_08DHFoOR;
R.RqRH:RM0R#8F_Do;HO
RRRq:dRRRHM#_08DHFoOR;
RRR7:MRHR8#0_oDFHPO_CFO0sR5(8MFI0jFR2R;
RBRWp:iRRRHM#_08DHFoOR;
R RWRH:RM0R#8F_Do
HOR
2;CRM8ObFlFMMC0V;
k0MOHRFMVOkM_HHM0R5L:FRLFNDCMs2RCs0kM0R#soHMR
H#LHCoMR
RH5VRL02RE
CMRRRRskC0s"M5hsFRC/N8I0sHCFROMHVDOO0RE	CO3HR1lNkD0MHFR#lHlON0EFRb#L#HD!CR!;"2
CRRD
#CRRRRskC0s"M5BDFk8FRM0lRHblDCCRM0AODF	qR)vQ3R#ER0CCRsNN8R8C8s#s#RC#oH0CCs8#RkHRMo0REC#CNlRFODON	R#ER0CqR)v2?";R
RCRM8H
V;CRM8VOkM_HHM0V;
k0MOHRFMo_C0C_M880CbEH5#x:CRR0HMCsoCR8;RCEb0RH:RMo0CCRs2skC0sHMRMo0CCHsR#N
PsLHNDlCRH#M_HRxC:MRH0CCos=R:R
j;LHCoMR
Rl_HM#CHxRR:=80CbER;
RRHV5x#HCRR<80CbE02RE
CMRRRRl_HM#CHxRR:=#CHx;R
RCRM8H
V;RCRs0MksRMlH_x#HCC;
Mo8RCC0_M88_CEb0;0
N0LsHkR0CoCCMsFN0sC_sb0FsR#:R0MsHoN;
0H0sLCk0RMoCC0sNFss_CsbF0VRFR_MFsOI_E	CORN:RsHOE00COkRsCHV#Rk_MOH0MH58N8sC_so
2;-L-RCMoHRFLDOs	RNHlRlCbDl0CMNF0HMHR#oDMN#$
0bHCRMN0_s$sNRRH#NNss$jR5RR0F6F2RVMRH0CCosO;
F0M#NRM0I0H8Es_NsRN$:MRH0s_NsRN$:5=R4.,R,,RcRRg,4RU,d;n2
MOF#M0N0CR8b_0ENNss$RR:H_M0NNss$=R:Rn54d,UcRgU4.c,Rj,gnRc.jU4,Rj,.cR.642O;
F0M#NRM08dHP.RR:HCM0oRCs:5=RI0H8E2-4/;dn
MOF#M0N0HR8PR4n:MRH0CCos=R:RH5I8-0E442/UO;
F0M#NRM08UHPRH:RMo0CC:sR=IR5HE80-/42gO;
F0M#NRM08cHPRH:RMo0CC:sR=IR5HE80-/42cO;
F0M#NRM08.HPRH:RMo0CC:sR=IR5HE80-/42.O;
F0M#NRM084HPRH:RMo0CC:sR=IR5HE80-/424
;
O#FM00NMRFLFD:4RRFLFDMCNRR:=5P8H4RR>j
2;O#FM00NMRFLFD:.RRFLFDMCNRR:=5P8H.RR>j
2;O#FM00NMRFLFD:cRRFLFDMCNRR:=5P8HcRR>j
2;O#FM00NMRFLFD:URRFLFDMCNRR:=5P8HURR>j
2;O#FM00NMRFLFDR4n:FRLFNDCM=R:RH58PR4n>2Rj;F
OMN#0ML0RFdFD.RR:LDFFCRNM:5=R8dHP.RR>j
2;
MOF#M0N0HR8Pd4nU:cRR0HMCsoCRR:=5b8C04E-2n/4d;Uc
MOF#M0N0HR8PgU4.RR:HCM0oRCs:5=R80CbE2-4/gU4.O;
F0M#NRM08cHPjRgn:MRH0CCos=R:RC58b-0E4c2/j;gn
MOF#M0N0HR8Pc.jURR:HCM0oRCs:5=R80CbE2-4/c.jUO;
F0M#NRM084HPjR.c:MRH0CCos=R:RC58b-0E442/j;.c
MOF#M0N0HR8P.64RH:RMo0CC:sR=8R5CEb0-/426;4.
F
OMN#0ML0RF6FD4:.RRFLFDMCNRR:=5P8H6R4.>2Rj;F
OMN#0ML0RF4FDjR.c:FRLFNDCM=R:RH58P.4jcRR>j
2;O#FM00NMRFLFDc.jURR:LDFFCRNM:5=R8.HPjRcU>2Rj;F
OMN#0ML0RFcFDjRgn:FRLFNDCM=R:RH58PgcjnRR>j
2;O#FM00NMRFLFDgU4.RR:LDFFCRNM:5=R8UHP4Rg.>2Rj;F
OMN#0ML0RF4FDncdURL:RFCFDN:MR=8R5HnP4dRUc>2Rj;O

F0M#NRM0#_klI0H8ERR:HCM0oRCs:A=Rm mpqbh'FL#5F4FD2RR+Apmm 'qhb5F#LDFF.+2RRmAmph q'#bF5FLFDRc2+mRAmqp hF'b#F5LF2DURA+Rm mpqbh'FL#5F4FDn
2;O#FM00NMRl#k_b8C0:ERR0HMCsoCRR:=6RR-5mAmph q'#bF5FLFD.642RR+Apmm 'qhb5F#LDFF4cj.2RR+Apmm 'qhb5F#LDFF.Ujc2RR+Apmm 'qhb5F#LDFFcnjg2RR+Apmm 'qhb5F#LDFFU.4g2
2;
MOF#M0N0_RIOHEFOIC_HE80RH:RMo0CC:sR=HRI8_0ENNss$k5#lH_I820E;F
OMN#0MI0R_FOEH_OC80CbERR:HCM0oRCs:8=RCEb0_sNsN#$5kIl_HE802O;
F0M#NRM08E_OFCHO_8IH0:ERR0HMCsoCRR:=I0H8Es_Ns5N$#_kl80CbE
2;O#FM00NMRO8_EOFHCC_8bR0E:MRH0CCos=R:Rb8C0NE_s$sN5l#k_b8C0;E2
F
OMN#0MI0R_8IH0ME_kOl_C#DDRH:RMo0CC:sR=IR5HE80-/42IE_OFCHO_8IH0+ERR
4;O#FM00NMR8I_CEb0_lMk_DOCD:#RR0HMCsoCRR:=5b8C04E-2_/IOHEFO8C_CEb0R4+R;O

F0M#NRM08H_I8_0EM_klODCD#RR:HCM0oRCs:5=RI0H8E2-4/O8_EOFHCH_I8R0E+;R4
MOF#M0N0_R880CbEk_MlC_ODRD#:MRH0CCos=R:RC58b-0E482/_FOEH_OC80CbERR+4
;
O#FM00NMR#I_HRxC:MRH0CCos=R:RII_HE80_lMk_DOCD*#RR8I_CEb0_lMk_DOCD
#;O#FM00NMR#8_HRxC:MRH0CCos=R:RI8_HE80_lMk_DOCD*#RR88_CEb0_lMk_DOCD
#;
MOF#M0N0FRLF8D_RL:RFCFDN:MR=8R5_x#HCRR-IH_#x<CR=2Rj;F
OMN#0ML0RF_FDIRR:LDFFCRNM:M=RFL05F_FD8
2;
MOF#M0N0EROFCHO_8IH0:ERR0HMCsoCRR:=5mAmph q'#bF5FLFD2_8R8*R_FOEH_OCI0H8E+2RRm5Amqp hF'b#F5LFID_2RR*IE_OFCHO_8IH0;E2
MOF#M0N0EROFCHO_b8C0:ERR0HMCsoCRR:=5mAmph q'#bF5FLFD2_8R8*R_FOEH_OC80CbE+2RRm5Amqp hF'b#F5LFID_2RR*IE_OFCHO_b8C0;E2
MOF#M0N0HRI8_0EM_klODCD#RR:HCM0oRCs:5=RApmm 'qhb5F#LDFF_R82*H5I8-0E482/_FOEH_OCI0H8E+2RRm5Amqp hF'b#F5LFID_2RR*58IH04E-2_/IOHEFOIC_HE802RR+4O;
F0M#NRM080CbEk_MlC_ODRD#:MRH0CCos=R:Rm5Amqp hF'b#F5LF8D_25R*80CbE2-4/O8_EOFHCC_8b20ER5+RApmm 'qhb5F#LDFF_RI2*8R5CEb0-/42IE_OFCHO_b8C0RE2+;R4
O--F0M#NRM0M_klODCD#RR:HCM0oRCs:5=R5C58bR0E-2R4Rd/R.+2RR55580CbERR-4l2RFd8R./2RR24n2R;RRR--yVRFRv)qd4.X1CRODRD#M8CCC
8R-F-OMN#0MD0RC_V0FsPCRH:RMo0CC:sR=5R55b8C0+ERR246R8lFR2d.R4/RnR2;RRRRRRRRRRRRRRRRRRRRRRRR-y-RRRFV)4qvn1X4RCMC8RC8VRFsD0CVRCFPsFRIs
8#0C$bR0Fk_#Lk4$_0bHCR#sRNsRN$5b8C0ME_kOl_C#DD-84RF0IMF,RjR8IH0ME_kOl_C#DD-84RF0IMF2RjRRFV#_08DHFoO#;
HNoMDkRF0k_L#:4RR0Fk_#Lk4$_0bRC;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RV_Rs80FkRM5HbRk000FRs#H-0CN0#02
$RbCF_k0L.k#_b0$C#RHRsNsN5$R80CbEk_MlC_OD-D#4FR8IFM0RRj,.H*I8_0EM_klODCD#R+48MFI0jFR2VRFR8#0_oDFH
O;#MHoNFDRkL0_kR#.:kRF0k_L#0._$;bCRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$FsVR_k8F0HR5M0bkRR0F0-sH#00NC
#20C$bR0Fk_#Lkc$_0bHCR#sRNsRN$5b8C0ME_kOl_C#DD-84RF0IMF,RjRIc*HE80_lMk_DOCDd#+RI8FMR0FjF2RV0R#8F_Do;HO
o#HMRNDF_k0Lck#RF:RkL0_k_#c0C$b;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFVsF_8k50RHkMb0FR0RH0s-N#002C#
b0$CkRF0k_L#0U_$RbCHN#Rs$sNRC58b_0EM_klODCD#R-48MFI0jFR,*RUI0H8Ek_MlC_OD+D#(FR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNR0Fk_#LkURR:F_k0LUk#_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFR8s_FRk05bHMk00RFsR0H0-#N#0C2$
0bbCRN0sH$k_L#0U_$RbCHN#Rs$sNRC58b_0EM_klODCD#R-48MFI0jFR,HRI8_0EM_klODCD#R-48MFI0jFR2VRFR8#0_oDFH
O;#MHoNbDRN0sH$k_L#:URRsbNH_0$LUk#_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$FsVR_k8F0HR5M0bkRR0F0-sH#00NC
#20C$bR0Fk_#Lk40n_$RbCHN#Rs$sNRC58b_0EM_klODCD#R-48MFI0jFR,nR4*8IH0ME_kOl_C#DD+R468MFI0jFR2VRFR8#0_oDFH
O;#MHoNFDRkL0_kn#4RF:RkL0_kn#4_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFR8s_FRk05bHMk00RFsR0H0-#N#0C2$
0bbCRN0sH$k_L#_4n0C$bRRH#NNss$8R5CEb0_lMk_DOCD4#-RI8FMR0Fj.,R*8IH0ME_kOl_C#DD+84RF0IMF2RjRRFV#_08DHFoO#;
HNoMDNRbs$H0_#Lk4:nRRsbNH_0$L4k#n$_0bRC;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFVsF_8k50RHkMb0FR0RH0s-N#002C#
b0$CkRF0k_L#_d.0C$bRRH#NNss$8R5CEb0_lMk_DOCD4#-RI8FMR0Fjd,R.H*I8_0EM_klODCD#4+dRI8FMR0FjF2RV0R#8F_Do;HO
o#HMRNDF_k0Ldk#.RR:F_k0Ldk#.$_0bRC;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RV_Rs80FkRM5HbRk000FRs#H-0CN0#02
$RbCbHNs0L$_k.#d_b0$C#RHRsNsN5$R80CbEk_MlC_OD-D#4FR8IFM0RRj,cH*I8_0EM_klODCD#R+d8MFI0jFR2VRFR8#0_oDFH
O;#MHoNbDRN0sH$k_L#Rd.:NRbs$H0_#Lkd0._$;bCRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFR8s_FRk05bHMk00RFsR0H0-#N#0C2H
#oDMNR0Fk_RCM:0R#8F_Do_HOP0COF8s5CEb0_lMk_DOCD4#-RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-C-RMDNLCV#RF0sRs#H-0CN0#H
#oDMNR0Is_RCM:0R#8F_Do_HOP0COF8s5CEb0_lMk_DOCD4#-RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-I-RsCH0RNCML#DCRsVFROCNEFRsIVRFRv)qRDOCD##
HNoMDMRH_osCR#:R0D8_FOoH_OPC05FsI0H8E6+dRI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RCk#8FR0RosCHC#0sQR7h#R
HNoMDkRF0C_soRR:#_08DHFoOC_POs0F58IH0dE+6FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RCk#8FR0RosCHC#0smR7z#a
HNoMDkRF0C_so:4RR8#0_oDFHPO_CFO0sH5I8-0E4FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--k8#CRR0FOFEF#LCRCC0IC7MRQNhRMF8Rkk0b0VRFRFADO)	Rq#v
HNoMD8RN_osCR#:R0D8_FOoH_OPC05FsNs88I0H8ER-48MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--k8#CRR0FsHCo#s0CR7q7)FRVssRIH
0C#MHoNDDRFsI_Ns88R#:R0D8_FOoH_OPC05Fs48dRF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-s-RNs88R0LH#MRHbRk00)FRqOvRC#DDRR5cL#H0RJsCkCHs8#2
HNoMDFRDIN_I8R8s:0R#8F_Do_HOP0COF4s5dFR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-NRI8R8sL#H0RbHMk00RFqR)vCRODRD#5LcRHR0#skCJH8sC2H
#oDMNR8sN8ss_C:oRR8#0_oDFHPO_CFO0s85N8HsI8-0E4FR8IFM0R;j2
R--CRM8LODF	NRsllRHblDCCNM00MHFRo#HM#ND
-
-RoLCH#MRCODC0NRsllRHblDCCNM00MHFRo#HM#ND
b0$CCRDVP0FC0s_RRH#NNss$jR5RR0FdF2RVMRH0CCos0;
$RbCD0CVFsPC_.0_RRH#NNss$jR5RR0F4F2RVMRH0CCosV;
k0MOHRFMb5N8HRR:#_08DHFoOC_POs0F;4RI,.RIRH:RMo0CCRs2skC0s#MR0D8_FOoH_OPC0RFsHP#
NNsHLRDCPRNs:0R#8F_Do_HOP0COFIs54R-48MFI0jFR2L;
CMoH
VRRF[sRRRHMP'NssoNMCFRDFRb
RHRRV[R5RR<=IR.20MECRR
SRsPN5R[2:H=R5DH'F[I+2S;
CCD#
RSRP5Ns[:2R=jR''S;
CRM8H
V;RMRC8FRDF
b;RCRs0MksRsPN;M
C8NRb8V;
k0MOHRFMo_C0I0H8E5_UI0H8EH:RMo0CCRs2skC0sHMRMo0CCHsR#N
PsLHNDPCRN:DRR0HMCsoCRR:=jL;
CMoH
PRRN:DR=HRI8/0EUR;
RRHV5H5I8R0ElRF8U>2RRRc20MEC
RRRRDPNRR:=PRND+;R4
CRRMH8RVR;
R0sCkRsMP;ND
8CMR0oC_8IH0UE_;k
VMHO0FoMRCI0_HE80_I.5HE80:MRH0CCoss2RCs0kMMRH0CCos#RH
sPNHDNLCNRPDRR:HCM0oRCs:j=R;C
Lo
HMRNRPD=R:R8IH0.E/;R
RskC0sPMRN
D;CRM8o_C0I0H8E;_.
MVkOF0HMCRo0H_I850EI0H8ERR:HCM0o2CsR0sCkRsMD0CVFsPC_.0_R
H#PHNsNCLDRDPNRD:RCFV0P_Cs0;_.
oLCHRM
RDPN5R42:o=RCI0_HE80_I.5HE802R;
RRHV58IH0lERF.8RRj=R2ER0CRM
RPRRNjD52=R:R
j;RDRC#RC
RPRRNjD52=R:R
4;RMRC8VRH;R
RskC0sPMRN
D;CRM8o_C0I0H8EV;
k0MOHRFMo_C0I0H8EH5I8R0E:MRH0CCoss2RCs0kMCRDVP0FC0s_R
H#PHNsNCLDRDPNRD:RCFV0P_Cs0=R:R,5jRRj,jj,R2L;
CMoH
PRRNdD52=R:R0oC_8IH0UE_58IH0;E2
ORRNR#C58IH0lERFU8R2#RH
IRRERCMcRR|d>R=RDPN5R.2:4=R;R
RIMECR=.R>NRPD254RR:=4R;
RCIEMRR4=P>RNjD52=R:R
4;RERICFMR0sEC#>R=RDMkDR;
R8CMR#ONCR;
R0sCkRsMP;ND
8CMR0oC_8IH0
E;O#FM00NMRI#_HE80_sNsN:$RRVDC0CFPsR_0:o=RCI0_HE8058IH0;E2
MOF#M0N0_R#I0H8Es_Ns_N$n:cRRVDC0CFPs__0.=R:R0oC_8IH0IE5HE802V;
k0MOHRFMo_C0M_kl45.U80CbEH:RMo0CCRs2skC0sHMRMo0CCHsR#N
PsLHNDPCRN:DRR0HMCsoCRR:=jL;
CMoH
PRRN:DR=CR8b/0E4;.U
HRRV5R580CbEFRl8.R4U>2RR.442ER0CRM
RPRRN:DR=NRPDRR+4R;
R8CMR;HV
sRRCs0kMNRPDC;
Mo8RCM0_k4l_.
U;VOkM0MHFR0oC_VDC0CFPsc_n5b8C0:ERR0HMCsoC2CRs0MksR0HMCsoCR
H#LHCoMR
RskC0s8M5CEb0R8lFRU4.2C;
Mo8RCD0_CFV0P_Csn
c;VOkM0MHFR0oC_lMk_5nc80CbERR:HCM0o2CsR0sCkRsMHCM0oRCsHP#
NNsHLRDCPRND:MRH0CCos=R:R
j;LHCoMR
RH5VR80CbE=R<R.44R8NMRb8C0>ERR2cURC0EMR
RRPRRN:DR=;R4
CRRMH8RVR;
R0sCkRsMP;ND
8CMR0oC_lMk_;nc
MVkOF0HMCRo0C_DVP0FC8s5CEb0RH:RMo0CCRs;lRNG:MRH0CCoss2RCs0kMMRH0CCos#RH
sPNHDNLCNRPDRR:HCM0oRCs:j=R;C
Lo
HMRVRHRC58bR0E-NRlG=R>RRj20MEC
RRRRDPNRR:=80CbERR-l;NG
CRRD
#CRRRRPRND:8=RCEb0;R
RCRM8H
V;RCRs0Mks5DPN2C;
Mo8RCD0_CFV0P;Cs
MVkOF0HMCRo0k_Ml._d5b8C0:ERR0HMCsoC2CRs0MksR0HMCsoCR
H#PHNsNCLDRDPNRH:RMo0CC:sR=;Rj
oLCHRM
RRHV5b8C0<ER=URcR8NMRb8C0>ERR24nRC0EMR
RRPRRN:DR=;R4
CRRMH8RVR;
R0sCkRsMP;ND
8CMR0oC_lMk_;d.
MVkOF0HMCRo0k_Mln_45b8C0:ERR0HMCsoC2CRs0MksR0HMCsoCR
H#PHNsNCLDRDPNRH:RMo0CC:sR=;Rj
oLCHRM
RRHV5b8C0<ER=nR4R8NMRb8C0>ERRRj20MEC
RRRRNRPD=R:R
4;RMRC8VRH;R
RskC0sPMRN
D;CRM8o_C0M_kl4
n;-F-OMN#0MM0RkOl_C#DDRH:RMo0CC:sR=5R55b8C0-ERRR42/.Rd2RR+5855CEb0R4-R2FRl8.Rd2RR/42n2;RRR-y-RRRFV)dqv.1X4RDOCDM#RCCC88OR
F0M#NRM0M_klODCD_U4.RH:RMo0CC:sR=CRo0k_Ml._4UC58b20E;F
OMN#0MD0RCFV0P_Csn:cRR0HMCsoCRR:=o_C0D0CVFsPC_5nc80CbE
2;O#FM00NMRlMk_DOCDc_nRH:RMo0CC:sR=CRo0k_Mlc_n5VDC0CFPsc_n2O;
F0M#NRM0D0CVFsPC_Rd.:MRH0CCos=R:R0oC_VDC0CFPsC5DVP0FCns_cn,Rc
2;O#FM00NMRlMk_DOCD._dRH:RMo0CC:sR=CRo0k_Ml._d5VDC0CFPs._d2O;
F0M#NRM0D0CVFsPC_R4n:MRH0CCos=R:R0oC_VDC0CFPsC5DVP0FCds_.d,R.
2;O#FM00NMRlMk_DOCDn_4RH:RMo0CC:sR=CRo0k_Mln_45VDC0CFPsn_42
;
0C$bR0Fk_#Lk_b0$C._4U#RHRsNsN5$RM_klODCD_U4.RI8FMR0FjI,RHE80-84RF0IMF2RjRRFV#_08DHFoO0;
$RbCF_k0L_k#0C$b_RncHN#Rs$sNRk5MlC_ODnD_cFR8IFM0RRj,I0H8ER-48MFI0jFR2VRFR8#0_oDFH
O;0C$bR0Fk_#Lk_b0$C._dRRH#NNss$MR5kOl_C_DDd8.RF0IMF,RjR8IH04E-RI8FMR0FjF2RV0R#8F_Do;HO
b0$CkRF0k_L#$_0b4C_n#RHRsNsN5$RM_klODCD_R4n8MFI0jFR,HRI8-0E4FR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNR0Fk_#Lk_U4.RF:RkL0_k0#_$_bC4;.URRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$F8VRFRk05bHMk00RFsR0H0-#N#0C2H
#oDMNR0Fk_#Lk_Rnc:kRF0k_L#$_0bnC_cR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFRk8F0HR5M0bkRR0F0-sH#00NC
#2#MHoNFDRkL0_kd#_.RR:F_k0L_k#0C$b_;d.RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$F8VRFRk05bHMk00RFsR0H0-#N#0C2H
#oDMNR0Fk_#Lk_R4n:kRF0k_L#$_0b4C_nR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFRk8F0HR5M0bkRR0F0-sH#00NC
#2#MHoN#DR_0Fk_RCM:0R#8F_Do_HOP0COFMs5kOl_C_DD4R.U8MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-MRCNCLD#FRVssR0H0-#N#0C
o#HMRNDF_k0CnM_cRR:#_08DHFoO#;
HNoMDkRF0M_C_Rd.:0R#8F_Do;HO
o#HMRNDF_k0C4M_nRR:#_08DHFoO#;
HNoMD_R#I_s0C:MRR8#0_oDFHPO_CFO0sk5MlC_OD4D_.8URF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RHIs0CCRMDNLCV#RFCsRNROEsRFIF)VRqOvRC#DD
o#HMRNDI_s0CnM_cRR:#_08DHFoO#;
HNoMDsRI0M_C_Rd.:0R#8F_Do;HO
o#HMRNDI_s0C4M_nRR:#_08DHFoO#;
HNoMD_R#HsM_C:oRR8#0_oDFHPO_CFO0sH5I8-0E4FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-#RkC08RFCRso0H#C7sRQ
hR#MHoN#DR_0Fk_osCR#:R0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-k-R#RC80sFRC#oH0RCs7amz
o#HMRND#8_N_osCR#:R0D8_FOoH_OPC05FsNs88I0H8ER-48MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--k8#CRR0FsHCo#s0CR7q7)H
#oDMNRIDF_8N8sRR:#_08DHFoOC_POs0F58nRF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-N-R8R8sL#H0RbHMk00RFqR)vCRODRD#5LcRHR0#skCJH8sC2F
OMN#0MD0R#IL_HE80RH:RMo0CC:sR=HRI8-0EU#*5_8IH0NE_s$sN5-d24c2-*I#_HE80_sNsN.$52*-.#H_I8_0ENNss$254-I#_HE80_sNsNj$520;
$RbC0_lbNNss$HUR#sRNsRN$5I#_HE80_sNsNd$52R-48MFI0jFR2VRFR8#0_oDFHPO_CFO0sR5(8MFI0jFR2#;
HNoMDlR0b__UdR.,0_lbUn_4R0:RlNb_s$sNU-;
-MRC8CR#D0CORlsNRbHlDCClM00NHRFM#MHoN
D#Ns00H0LkC3R\s_NlF#VVCR0\:0R#soHM;L

CMoH

RRRcRzdRR:H5VRNs88_osC2CRoMNCs0-CR-CRoMNCs0LCRD	FORlsN
RRRRR--QNVR8I8sHE80RO<REOFHCH_I8R0ENH##o'MRj0'RFMRkk8#CR0LH#R
RRjRzRRR:H5VRNs88I0H8ERR=4o2RCsMCN
0CRRRRRRRRD_FIs8N8s=R<Rj"jjjjjjjjjj"jjRq&R757)j
2;RRRRRRRRD_FII8N8s=R<Rj"jjjjjjjjjj"jjRN&R8C_so25j;R
RRMRC8CRoMNCs0zCRjR;
RzRR4:RRRRHV58N8s8IH0=ERRR.2oCCMsCN0
RRRRRRRRIDF_8sN8<sR=jR"jjjjjjjjj"jjRq&R757)4FR8IFM0R;j2
RRRRRRRRIDF_8IN8<sR=jR"jjjjjjjjj"jjRN&R8C_soR548MFI0jFR2R;
RCRRMo8RCsMCNR0Cz
4;RRRRzR.R:VRHR85N8HsI8R0E=2RdRMoCC0sNCR
RRRRRRFRDIN_s8R8s<"=Rjjjjjjjjj"jjRq&R757).FR8IFM0R;j2
RRRRRRRRIDF_8IN8<sR=jR"jjjjjjjjjRj"&8RN_osC58.RF0IMF2Rj;R
RRMRC8CRoMNCs0zCR.R;
RzRRd:RRRRHV58N8s8IH0=ERRRc2oCCMsCN0
RRRRRRRRIDF_8sN8<sR=jR"jjjjjjjjj&"RR7q7)R5d8MFI0jFR2R;
RRRRRDRRFII_Ns88RR<="jjjjjjjj"jjRN&R8C_soR5d8MFI0jFR2R;
RCRRMo8RCsMCNR0Cz
d;RRRRzRcR:VRHR85N8HsI8R0E=2R6RMoCC0sNCR
RRRRRRFRDIN_s8R8s<"=Rjjjjjjjjj&"RR7q7)R5c8MFI0jFR2R;
RRRRRDRRFII_Ns88RR<="jjjjjjjjRj"&8RN_osC58cRF0IMF2Rj;R
RRMRC8CRoMNCs0zCRcR;
RzRR6:RRRRHV58N8s8IH0=ERRRn2oCCMsCN0
RRRRRRRRIDF_8sN8<sR=jR"jjjjj"jjRq&R757)6FR8IFM0R;j2
RRRRRRRRIDF_8IN8<sR=jR"jjjjj"jjRN&R8C_soR568MFI0jFR2R;
RCRRMo8RCsMCNR0Cz
6;RRRRzRnR:VRHR85N8HsI8R0E=2R(RMoCC0sNCR
RRRRRRFRDIN_s8R8s<"=Rjjjjj"jjRq&R757)nFR8IFM0R;j2
RRRRRRRRIDF_8IN8<sR=jR"jjjjjRj"&8RN_osC58nRF0IMF2Rj;R
RRMRC8CRoMNCs0zCRnR;
RzRR(:RRRRHV58N8s8IH0=ERRRU2oCCMsCN0
RRRRRRRRIDF_8sN8<sR=jR"jjjjj&"RR7q7)R5(8MFI0jFR2R;
RRRRRDRRFII_Ns88RR<="jjjj"jjRN&R8C_soR5(8MFI0jFR2R;
RCRRMo8RCsMCNR0Cz
(;RRRRzRUR:VRHR85N8HsI8R0E=2RgRMoCC0sNCR
RRRRRRFRDIN_s8R8s<"=Rjjjjj&"RR7q7)R5U8MFI0jFR2R;
RRRRRDRRFII_Ns88RR<="jjjjRj"&8RN_osC58URF0IMF2Rj;R
RRMRC8CRoMNCs0zCRUR;
RzRRg:RRRRHV58N8s8IH0=ERR24jRMoCC0sNCR
RRRRRRFRDIN_s8R8s<"=Rjjjj"RR&q)7758gRF0IMF2Rj;R
RRRRRRFRDIN_I8R8s<"=Rjjjj"RR&Ns8_Cgo5RI8FMR0Fj
2;RRRRCRM8oCCMsCN0R;zg
RRRRjz4RRR:H5VRNs88I0H8ERR=4R42oCCMsCN0
RRRRRRRRIDF_8sN8<sR=jR"jRj"&7Rq74)5jFR8IFM0R;j2
RRRRRRRRIDF_8IN8<sR=jR"jRj"&8RN_osC5R4j8MFI0jFR2R;
RCRRMo8RCsMCNR0Cz;4j
RRRR4z4RRR:H5VRNs88I0H8ERR=4R.2oCCMsCN0
RRRRRRRRIDF_8sN8<sR=jR"j&"RR7q7)454RI8FMR0Fj
2;RRRRRRRRD_FII8N8s=R<Rj"j"RR&Ns8_C4o54FR8IFM0R;j2
RRRR8CMRMoCC0sNC4Rz4R;
RzRR4R.R:VRHR85N8HsI8R0E=dR42CRoMNCs0RC
RRRRRDRRFsI_Ns88RR<='Rj'&7Rq74)5.FR8IFM0R;j2
RRRRRRRRIDF_8IN8<sR=jR''RR&Ns8_C4o5.FR8IFM0R;j2
RRRR8CMRMoCC0sNC4Rz.R;
RzRR4RdR:VRHR85N8HsI8R0E>dR42CRoMNCs0RC
RRRRRDRRFsI_Ns88RR<=q)775R4d8MFI0jFR2R;
RRRRRDRRFII_Ns88RR<=Ns8_C4o5dFR8IFM0R;j2
RRRR8CMRMoCC0sNC4Rzd
;
RRRR-Q-RV8R5HsM_CRo2sHCo#s0CRh7QRHk#MBoRpRi
RzRR4RcR:VRHRH58MC_soo2RCsMCN
0CRRRRRRRRbOsFCR##5iBp,QR7hL2RCMoH
RRRRRRRRRRRRRHV5iBpR'=R4N'RMB8RpCi'P0CM2ER0CRM
RRRRRRRRRRRRRHRRMC_so=R<Rj5"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jjR7&RQ;h2
RRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMRFbsO#C#;R
RRMRC8CRoMNCs0zCR4
c;RRRRzR46RH:RVMR5F80RHsM_CRo2oCCMsCN0
RRRRRRRRRRRR_HMsRCo<5=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj&"RRh7Q2R;
RCRRMo8RCsMCNR0Cz;46
R
RR-R-RRQV5Fs8ks0_CRo2sHCo#s0CR7)_mRzakM#Ho_R)miBp
RRRRnz4RRR:H5VR80Fk_osC2CRoMNCs0RC
RRRRRbRRsCFO#5#RmiBp,kRF0C_soR42LHCoMR
RRRRRRRRRRVRHRB5mp=iRR''4R8NMRpmBiP'CC2M0RC0EMR
RRRRRRRRRRRRRRmR7z<aR=kRF0C_so
4;RRRRRRRRRRRRCRM8H
V;RRRRRRRRCRM8bOsFC;##
RRRRRRRR8CMRMoCC0sNC4RznR;
RzRR4R(R:VRHRF5M0FR8ks0_CRo2oCCMsCN0
RRRRRRRRRRRRz7ma=R<R0Fk_osC4R;
RCRRMo8RCsMCNR0Cz;4(
R
RR-R-RRQV58N8sC_sos2RC#oH0RCsq)77RsVFRHIs0kCR#oHMRiBp
RRRRUz4I:RRRRHV58N8sC_soo2RCsMCN
0CRRRRRRRRbOsFCR##5iBp,7Rq7R)2LHCoMR
RRRRRRRRRRVRHRp5BiRR='R4'NRM8B'piCMPC002RE
CMRRRRRRRRRRRRRRRRNs8_C<oR=7Rq7N)58I8sHE80-84RF0IMF2Rj;R
RRRRRRRRRRMRC8VRH;R
RRRRRRMRC8sRbF#OC#R;
RCRRMo8RCsMCNR0CzI4U;R
RR4Rzg:IRRRHV50MFR8N8sC_soo2RCsMCN
0CRRRRRRRRRRRRNs8_C<oR=7Rq7
);RRRRCRM8oCCMsCN0Rgz4I
;
RRRR- -RGN0sRoDFHVORF7sRkRNDb0FsR#ONC-
S-FR7R0MFRCMC8ER0HV#RFMsRFDRoFRkCDHFoOFROM08HH
FM-R-RRsRzC:oRRFbsO#C#5iBp2CRLo
HM-R-RRRRRH5VRB'pi he aMRN8pRBiRR='24'RC0EM-
-RRRRR7RRQ0h_l<bR=QR7h-;
-RRRRRRR)7q7)l_0b=R<R7q7)-;
-RRRRRRRW7q7)l_0b=R<R_N8s;Co
R--RRRRR RW_b0lRR<=W
 ;-R-RRRRRCRM8H
V;-R-RRMRC8sRbF#OC#
;
RRRRzGlkRb:RsCFO#F#5ks0_C
o2RRRRRCRLo
HM-R-RRRRRRVRHRq5W7_7)0Rlb=qR)7_7)0RlbNRM8W0 _l=bRR''42ER0C-M
-RRRRRRRRFRRks0_CRo4<7=RQ0h_l
b;-R-RRRRRRDRC#RC
RRRRRRRRR0Fk_osC4=R<R0Fk_osC58IH04E-RI8FMR0Fj
2;-R-RRRRRRMRC8VRH;R
RRMRC8sRbF#OC#R;
RRRRR
RRRRRR-t-RCsMCNR0C0REC)RqvODCD#MRN8CR#D0CORoDFHVORF)sRq4vAn4_1_
14RRRRzR4U:VRHRE5OFCHO_8IH0=ERRR42oCCMsCN0
-S-RGVHRsVFRDONDdR4U,U(RD#CCRO0F0VRs0H#NR0CMRF0LMCHoCRso0H#C8sC
RSRRRRRz	OERH:RVRR5Ns88I0H8ERR>4Rc2oCCMsCN0
RRRRRRRRRRRRDkO	b:RsCFO#B#5p
i2RRRRRRRRRRRRRoLCHRM
RRRRRRRRRRRRRRHV5iBp'CCPMN0RMB8Rp=iRR''42ER0CRM
RRRRRRRRRRRRRsRRNs88_osC58N8s8IH04E-RI8FMR0F4Rc2<q=R757)Ns88I0H8ER-48MFI04FRc
2;RRRRRRRRRRRRRMRC8VRH;R
RRRRRRRRRRMRC8sRbF#OC#S;
SCRRMo8RCsMCNR0Cz	OE;R
RRRRRR4RzgRR:VRFsHMRHRC58b_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
RRRRR--Q5VRNs88I0H8ERR>4Rc2M8CCRR0FONsC0ICRsCH0RNCMLRDCNRM8Fbk0kC0RMDNLCCR#D0CORoDFHRO
RRRRRRRRRzRR.:jRRRHV58N8s8IH0>ERR24cRMoCC0sNC-
S-HRVGFRVsNROD4DRd(UU,CR#D0CORRFV0#sH0CN0R0MFRHLCMsoRC#oH0CCs8R
RRRRRRRRRRRRRRkRF0M_C5RH2<'=R4I'RERCM58sN8ss_CNo58I8sHE80-84RF0IMFcR42RR=HC2RDR#C';j'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RWRCIEMNR58C_so85N8HsI8-0E4FR8IFM0R24cRH=R2DRC#'CRj
';RRRRRRRRRRRRCRM8oCCMsCN0Rjz.;R
RR-R-RRQV58N8s8IH0<ER=cR42FRMRHIs0CCRMDNLCsRFR0FkbRk0CLMND#CRCODC0FRDoRHOM8CCCR8
RRRRRRRRRzRR.:4RRRHV58N8s8IH0<ER=cR42CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_M25HRR<=';4'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RW;R
RRRRRRRRRRMRC8CRoMNCs0zCR.
4;RRRR-t-RCsMCNR0C0REC)RqvODCD#MRN8sR0H0-#N#0C
RRRRRRRRRRRR.z.RV:RF[sRRRHM58IH0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CRRRRRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FAVR)_qv4Undc7X4RD:RNDLCRRH#";W"
RRRRRRRRRRRRRRRRoLCHRM
RRRRRRRRRRRRRARR)_qv4Undc7X4R):Rq4vAn4_1_
14RRRRRRRRRRRRRRRRb0FsRblNRQ57q25jRR=>HsM_C[o52q,R7q7)RR=>D_FII8N8sd54RI8FMR0FjR2,7RQA=">RjR",q)77A>R=RIDF_8sN84s5dFR8IFM0R,j2
RRRRRRRRRRRRRRRRq hRR=>',4'R)11q>R=R''j, RWq>R=R0Is_5CMHR2,BqpiRR=>B,piRA hRR=>',4'R)11A>R=R''j, RWA>R=R''j,pRBi=AR>pRBiR,
RRRRRRRRRRRRR7RRm=qR>bRFCRM,75mAj=2R>kRF0k_L#H45,2[2;R

RRRRRRRRRRRRRFRRks0_C[o52=R<R0Fk_#Lk4,5H[I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRCRM8oCCMsCN0R.z.;R
RRRRRRMRC8CRoMNCs0zCR4
g;RRRRCRM8oCCMsCN0RUz4;RRRRR
RRRRR
RRRRR--tCCMsCN0RC0ERv)qRDOCDN#RM#8RCODC0FRDoRHOVRFs)Aqv41n_.._1
RRRRdz.RH:RVOR5EOFHCH_I8R0E=2R.RMoCC0sNC-
S-HRVGFRVsNROD4DRd(UU,CR#D0CORRFV0#sH0CN0R0MFRHLCMsoRC#oH0CCs8R
SRRRRz	OE:VRHR85N8HsI8R0E>dR42CRoMNCs0RC
RRRRRRRRRkRRO:D	RFbsO#C#5iBp2R
RRRRRRRRRRLRRCMoH
RRRRRRRRRRRRHRRVBR5pCi'P0CMR8NMRiBpR'=R4R'20MEC
RRRRRRRRRRRRRRRR8sN8ss_CNo58I8sHE80-84RF0IMFdR42=R<R7q7)85N8HsI8-0E4FR8IFM0R24d;R
RRRRRRRRRRRRRCRM8H
V;RRRRRRRRRRRRCRM8bOsFC;##
RSSCRM8oCCMsCN0REzO	R;
RRRRRzRR.:cRRsVFRHHRM8R5CEb0_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNCR
RR-R-RRQV58N8s8IH0>ERR24dRCMC8FR0RCOsNR0CI0sHCMRCNCLDR8NMR0FkbRk0CLMND#CRCODC0FRDo
HORRRRRRRRRRRRzR.6:VRHR85N8HsI8R0E>dR42CRoMNCs0SC
-V-RHVGRFOsRNRDD4UdU(#,RCODC0VRFRH0s#00NCFRM0CRLHRMosHCo#s0CCR8
RRRRRRRRRRRRRFRRkC0_M25HRR<='R4'IMECRN5s8_8ss5CoNs88I0H8ER-48MFI04FRd=2RRRH2CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R ERIC5MRNs8_CNo58I8sHE80-84RF0IMFdR42RR=HC2RDR#C';j'
RRRRRRRRRRRR8CMRMoCC0sNC.Rz6R;
R-RR-VRQR85N8HsI8R0E<4=RdM2RFsRIHR0CCLMNDFCRskRF00bkRNCMLRDC#CCDOD0RFOoHRCMC8
C8RRRRRRRRRRRRzR.n:VRHR85N8HsI8R0E<4=Rdo2RCsMCN
0CRRRRRRRRRRRRRRRRF_k0CHM52=R<R''4;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R R;
RRRRRRRRRCRRMo8RCsMCNR0Cz;.n
RRRRR--tCCMsCN0RC0ERv)qRDOCDN#RM08Rs#H-0CN0#R
RRRRRRRRRR.Rz(RR:VRFs[MRHRH5I8_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
RRRRRRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVAv)q_gU4.7X.RD:RNDLCRRH#";W"
RRRRRRRRRRRRRRRRoLCHRM
RRRRRRRRRRRRRARR)_qvU.4gXR.7:qR)vnA4__1.1R.
RRRRRRRRRRRRRbRRFRs0lRNb5q7QRR=>HsM_C.o5*4[+RI8FMR0F.2*[,7Rq7R)q=D>RFII_Ns885R4.8MFI0jFR27,RQ=AR>jR"jR",q)77A>R=RIDF_8sN84s5.FR8IFM0R,j2
RRRRRRRRRRRRRRRRq hRR=>',4'R)11q>R=R''j, RWq>R=R0Is_5CMHR2,BqpiRR=>B,piRA hRR=>',4'R)11A>R=R''j, RWA>R=R''j,pRBi=AR>pRBiR,
RRRRRRRRRRRRR7RRm=qR>bRFCRM,75mA4=2R>kRF0k_L#H.5,[.*+,42RA7m5Rj2=F>RkL0_k5#.H.,R*2[2;R
RRRRRRRRRRRRRRkRF0C_so*5.[<2R=kRF0k_L#H.5,[.*2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C.o5*4[+2=R<R0Fk_#Lk.,5H.+*[4I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRCRM8oCCMsCN0R(z.;R
RRRRRRMRC8CRoMNCs0zCR.
c;RRRRCRM8oCCMsCN0Rdz.;
RR
RRRRRRRRR--tCCMsCN0RC0ERv)qRDOCDN#RM#8RCODC0FRDoRHOVRFs)Aqv41n_cc_1
RRRRUz.RH:RVOR5EOFHCH_I8R0E=2RcRMoCC0sNC-
S-HRVGFRVsNROD4DRd(UU,CR#D0CORRFV0#sH0CN0R0MFRHLCMsoRC#oH0CCs8R
SRRRRREzO	H:RVNR58I8sHE80R4>R.o2RCsMCN
0CRRRRRRRRRRRRk	OD:sRbF#OC#p5BiR2
RRRRRRRRRRRRLHCoMR
RRRRRRRRRRRRRH5VRB'piCMPC0MRN8pRBiRR='24'RC0EMR
RRRRRRRRRRRRRRNRs8_8ss5CoNs88I0H8ER-48MFI04FR.<2R=7Rq7N)58I8sHE80-84RF0IMF.R42R;
RRRRRRRRRRRRR8CMR;HV
RRRRRRRRRRRR8CMRFbsO#C#;S
SRMRC8CRoMNCs0zCRO;E	
RRRRRRRRgz.RV:RFHsRRRHM5b8C0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CRRRR-Q-RVNR58I8sHE80R4>R.M2RCRC80OFRs0CNCsRIHR0CCLMNDNCRMF8Rkk0b0MRCNCLDRD#CCRO0DHFoOR
RRRRRRRRRRdRzjRR:H5VRNs88I0H8ERR>4R.2oCCMsCN0
-S-RGVHRsVFRDONDdR4U,U(RD#CCRO0F0VRs0H#NR0CMRF0LMCHoCRso0H#C8sC
RRRRRRRRRRRRRRRR0Fk_5CMH<2R=4R''ERIC5MRs8N8sC_so85N8HsI8-0E4FR8IFM0R24.RH=R2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0CHM52=R<RRW IMECR85N_osC58N8s8IH04E-RI8FMR0F4R.2=2RHR#CDCjR''R;
RRRRRRRRRCRRMo8RCsMCNR0Cz;dj
RRRRR--Q5VRNs88I0H8E=R<R24.RRMFI0sHCMRCNCLDRRFsFbk0kC0RMDNLCCR#D0CORoDFHMORCCC88R
RRRRRRRRRRdRz4RR:H5VRNs88I0H8E=R<R24.RMoCC0sNCR
RRRRRRRRRRRRRRkRF0M_C5RH2<'=R4
';RRRRRRRRRRRRRRRRI_s0CHM52=R<R;W 
RRRRRRRRRRRR8CMRMoCC0sNCdRz4R;
R-RR-CRtMNCs00CRE)CRqOvRC#DDR8NMRH0s-N#00
C#RRRRRRRRRRRRzRd.:FRVsRR[H5MRI0H8Ek_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0RC
RRRRRRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)RAqcv_jXgnc:7RRLDNCHDR#WR""R;
RRRRRRRRRRRRRLRRCMoH
RRRRRRRRRRRRRRRRqA)vj_cgcnX7RR:)Aqv41n_cc_1
RRRRRRRRRRRRRRRRsbF0NRlb7R5Q=qR>MRH_osC5[c*+8dRF0IMF*Rc[R2,q)77q>R=RIDF_8IN84s54FR8IFM0R,j2RA7QRR=>"jjjjR",q)77A>R=RIDF_8sN84s54FR8IFM0R,j2
RRRRRRRRRRRRRRRRq hRR=>',4'R)11q>R=R''j, RWq>R=R0Is_5CMHR2,BqpiRR=>B,piRA hRR=>',4'R)11A>R=R''j, RWA>R=R''j,pRBi=AR>pRBiR,
RRRRRRRRRRRRR7RRm=qR>bRFCRM,75mAd=2R>kRF0k_L#Hc5,*Rc[2+d,mR7A25.RR=>F_k0Lck#5cH,*.[+2
,RRRRRRRRRRRRRRRRR75mA4=2R>kRF0k_L#Hc5,[c*+,42RA7m5Rj2=F>RkL0_k5#cHc,R*2[2;R
RRRRRRRRRRRRRRkRF0C_so*5c[<2R=kRF0k_L#Hc5,[c*2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cco5*4[+2=R<R0Fk_#Lkc,5Hc+*[4I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Coc+*[.<2R=kRF0k_L#Hc5,[c*+R.2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5[c*+Rd2<F=RkL0_k5#cH*,c[2+dRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R

RRRRRRRRRCRRMo8RCsMCNR0Cz;d.
RRRRRRRR8CMRMoCC0sNC.RzgR;
RCRRMo8RCsMCNR0Cz;.U
R
RRRRRR-R-RMtCC0sNCER0CqR)vCRODRD#NRM8#CCDOD0RFOoHRsVFRv)qA_4n11g_gR
RRdRzdRR:H5VROHEFOIC_HE80Rg=R2CRoMNCs0SC
-V-RHVGRFOsRNRDD4UdU(#,RCODC0VRFRH0s#00NCFRM0CRLHRMosHCo#s0CCS8
RRRRRORzER	:H5VRNs88I0H8ERR>4R42oCCMsCN0
RRRRRRRRRRRRDkO	b:RsCFO#B#5p
i2RRRRRRRRRRRRRoLCHRM
RRRRRRRRRRRRRRHV5iBp'CCPMN0RMB8Rp=iRR''42ER0CRM
RRRRRRRRRRRRRsRRNs88_osC58N8s8IH04E-RI8FMR0F4R42<q=R757)Ns88I0H8ER-48MFI04FR4
2;RRRRRRRRRRRRRMRC8VRH;R
RRRRRRRRRRMRC8sRbF#OC#S;
SCRRMo8RCsMCNR0Cz	OE;R
RRRRRRdRzcRR:VRFsHMRHRC58b_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
RRRRR--Q5VRNs88I0H8ERR>4R42M8CCRR0FONsC0ICRsCH0RNCMLRDCNRM8Fbk0kC0RMDNLCCR#D0CORoDFHRO
RRRRRRRRRzRRd:6RRRHV58N8s8IH0>ERR244RMoCC0sNC-
S-HRVGFRVsNROD4DRd(UU,CR#D0CORRFV0#sH0CN0R0MFRHLCMsoRC#oH0CCs8R
RRRRRRRRRRRRRRkRF0M_C5RH2<'=R4I'RERCM58sN8ss_CNo58I8sHE80-84RF0IMF4R42RR=HC2RDR#C';j'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RWRCIEMNR58C_so85N8HsI8-0E4FR8IFM0R244RH=R2DRC#'CRj
';RRRRRRRRRRRRCRM8oCCMsCN0R6zd;R
RR-R-RRQV58N8s8IH0<ER=4R42FRMRHIs0CCRMDNLCsRFR0FkbRk0CLMND#CRCODC0FRDoRHOM8CCCR8
RRRRRRRRRzRRd:nRRRHV58N8s8IH0<ER=4R42CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_M25HRR<=';4'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RW;R
RRRRRRRRRRMRC8CRoMNCs0zCRd
n;RRRR-t-RCsMCNR0C0REC)RqvODCD#MRN8sR0H0-#N#0C
RRRRRRRRRRRR(zdRV:RF[sRRRHM58IH0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CRRRRRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FAVR)_qv.UjcXRU7:NRDLRCDH"#RW
";RRRRRRRRRRRRRRRRLHCoMR
RRRRRRRRRRRRRR)RAq.v_jXcUU:7RRv)qA_4n11g_gR
RRRRRRRRRRRRRRRRRb0FsRblNRQ57q>R=R_HMs5Cog+*[(FR8IFM0R[g*2q,R7q7)RR=>D_FII8N8sj54RI8FMR0FjR2,7RQA=">Rjjjjjjjj"q,R7A7)RR=>D_FIs8N8sj54RI8FMR0Fj
2,RRRRRRRRRRRRRRRR Rhq='>R4R',1q1)RR=>',j'RqW RR=>I_s0CHM52B,RpRiq=B>RpRi, RhA='>R4R',1A1)RR=>',j'RAW RR=>',j'RiBpA>R=RiBp,RR
RRRRRRRRRRRRR7RRm=qR>bRFCRM,75mA(=2R>kRF0k_L#HU5,[U*+,(2RA7m5Rn2=F>RkL0_k5#UH*,U[2+n,RR
RRRRRRRRRRRRR7RRm6A52>R=R0Fk_#LkU,5HU+*[6R2,75mAc=2R>kRF0k_L#HU5,[U*+,c2RA7m5Rd2=F>RkL0_k5#UH*,U[2+d,RR
RRRRRRRRRRRRR7RRm.A52>R=R0Fk_#LkU,5HU+*[.R2,75mA4=2R>kRF0k_L#HU5,[U*+,42RA7m5Rj2=F>RkL0_k5#UH*,U[
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRR7qQu5Rj2=H>RMC_so*5g[2+U,QR7u=AR>jR""7,RmRuq=F>Rb,CMRu7mA25jRR=>bHNs0L$_k5#UH[,R2
2;RRRRRRRRRRRRRRRRF_k0s5Cog2*[RR<=F_k0LUk#5UH,*R[2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5[g*+R42<F=RkL0_k5#UH*,U[2+4RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so*5g[2+.RR<=F_k0LUk#5UH,*.[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cgo5*d[+2=R<R0Fk_#LkU,5HU+*[dI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cog+*[c<2R=kRF0k_L#HU5,[U*+Rc2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5[g*+R62<F=RkL0_k5#UH*,U[2+6RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so*5g[2+nRR<=F_k0LUk#5UH,*n[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cgo5*([+2=R<R0Fk_#LkU,5HU+*[(I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cog+*[U<2R=NRbs$H0_#LkU,5H[I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRCRM8oCCMsCN0R(zd;R
RRRRRRMRC8CRoMNCs0zCRd
c;RRRRCRM8oCCMsCN0Rdzd;R

RRRRR-RR-CRtMNCs00CRE)CRqOvRC#DDR8NMRD#CCRO0DHFoOFRVsqR)vnA4_U14_U14
RRRRUzdRH:RVOR5EOFHCH_I8R0E=UR42CRoMNCs0SC
-V-RHVGRFOsRNRDD4UdU(#,RCODC0VRFRH0s#00NCFRM0CRLHRMosHCo#s0CCS8
RRRRRORzER	:H5VRNs88I0H8ERR>4Rj2oCCMsCN0
RRRRRRRRRRRRDkO	b:RsCFO#B#5p
i2RRRRRRRRRRRRRoLCHRM
RRRRRRRRRRRRRRHV5iBp'CCPMN0RMB8Rp=iRR''42ER0CRM
RRRRRRRRRRRRRsRRNs88_osC58N8s8IH04E-RI8FMR0F4Rj2<q=R757)Ns88I0H8ER-48MFI04FRj
2;RRRRRRRRRRRRRMRC8VRH;R
RRRRRRRRRRMRC8sRbF#OC#S;
SCRRMo8RCsMCNR0Cz	OE;R
RRRRRRdRzgRR:VRFsHMRHRC58b_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
RRRRR--Q5VRNs88I0H8ERR>4Rj2M8CCRR0FONsC0ICRsCH0RNCMLRDCNRM8Fbk0kC0RMDNLCCR#D0CORoDFHRO
RRRRRRRRRzRRc:jRRRHV58N8s8IH0>ERR24jRMoCC0sNC-
S-HRVGFRVsNROD4DRd(UU,CR#D0CORRFV0#sH0CN0R0MFRHLCMsoRC#oH0CCs8R
RRRRRRRRRRRRRRkRF0M_C5RH2<'=R4I'RERCM58sN8ss_CNo58I8sHE80-84RF0IMFjR42RR=HC2RDR#C';j'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RWRCIEMNR58C_so85N8HsI8-0E4FR8IFM0R24jRH=R2DRC#'CRj
';RRRRRRRRRRRRCRM8oCCMsCN0Rjzc;R
RR-R-RRQV58N8s8IH0<ER=jR42FRMRHIs0CCRMDNLCsRFR0FkbRk0CLMND#CRCODC0FRDoRHOM8CCCR8
RRRRRRRRRzRRc:4RRRHV58N8s8IH0<ER=jR42CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_M25HRR<=';4'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RW;R
RRRRRRRRRRMRC8CRoMNCs0zCRc
4;RRRR-t-RCsMCNR0C0REC)RqvODCD#MRN8sR0H0-#N#0C
RRRRRRRRRRRR.zcRV:RF[sRRRHM58IH0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CRRRRRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FAVR)_qv4cj.X74nRD:RNDLCRRH#";W"
RRRRRRRRRRRRRRRRoLCHRM
RRRRRRRRRRRRRARR)_qv4cj.X74nR):Rq4vAn4_1U4_1UR
RRRRRRRRRRRRRRRRRb0FsRblNRQ57q>R=R_HMs5Co4[U*+R468MFI04FRU2*[,7Rq7R)q=D>RFII_Ns8858gRF0IMF2Rj,QR7A>R=Rj"jjjjjjjjjjjjjj,j"R7q7)=AR>FRDIN_s858sgFR8IFM0R,j2
RRRRRRRRRRRRRRRRq hRR=>',4'R)11q>R=R''j, RWq>R=R0Is_5CMHR2,BqpiRR=>B,piRA hRR=>',4'R)11A>R=R''j, RWA>R=R''j,pRBi=AR>pRBi
,RRRRRRRRRRRRRRRRR7Rmq=F>Rb,CMRA7m5246RR=>F_k0L4k#n,5H4[n*+246,mR7Ac542>R=R0Fk_#Lk4Hn5,*4n[c+42
,RRRRRRRRRRRRRRRRR75mA4Rd2=F>RkL0_kn#454H,n+*[4,d2RA7m524.RR=>F_k0L4k#n,5H4[n*+24.,mR7A4542>R=R0Fk_#Lk4Hn5,*4n[4+42
,RRRRRRRRRRRRRRRRR75mA4Rj2=F>RkL0_kn#454H,n+*[4,j2RA7m5Rg2=F>RkL0_kn#454H,n+*[gR2,75mAU=2R>kRF0k_L#54nHn,4*U[+2
,RRRRRRRRRRRRRRRRR75mA(=2R>kRF0k_L#54nHn,4*([+27,RmnA52>R=R0Fk_#Lk4Hn5,*4n[2+n,mR7A256RR=>F_k0L4k#n,5H4[n*+,62RR
RRRRRRRRRRRRRRmR7A25cRR=>F_k0L4k#n,5H4[n*+,c2RA7m5Rd2=F>RkL0_kn#454H,n+*[dR2,75mA.=2R>kRF0k_L#54nHn,4*.[+2
,RRRRRRRRRRRRRRRRR75mA4=2R>kRF0k_L#54nHn,4*4[+27,RmjA52>R=R0Fk_#Lk4Hn5,*4n[R2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRu7Qq>R=R_HMs5Co4[U*+R4(8MFI04FRU+*[4,n2Ru7QA>R=Rj"j"R,
RRRRRRRRRRRRRRRRRRRRRRRRR7RRmRuq=F>Rb,CMRu7mA254RR=>bHNs0L$_kn#45RH,.+*[4R2,7Amu5Rj2=b>RN0sH$k_L#54nH.,R*2[2;R
RRRRRRRRRRRRRRkRF0C_soU54*R[2<F=RkL0_kn#454H,n2*[RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*4[+2=R<R0Fk_#Lk4Hn5,*4n[2+4RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*.[+2=R<R0Fk_#Lk4Hn5,*4n[2+.RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*d[+2=R<R0Fk_#Lk4Hn5,*4n[2+dRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*c[+2=R<R0Fk_#Lk4Hn5,*4n[2+cRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*6[+2=R<R0Fk_#Lk4Hn5,*4n[2+6RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*n[+2=R<R0Fk_#Lk4Hn5,*4n[2+nRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*([+2=R<R0Fk_#Lk4Hn5,*4n[2+(RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*U[+2=R<R0Fk_#Lk4Hn5,*4n[2+URCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*g[+2=R<R0Fk_#Lk4Hn5,*4n[2+gRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*4[+j<2R=kRF0k_L#54nHn,4*4[+jI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+244RR<=F_k0L4k#n,5H4[n*+244RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*4[+.<2R=kRF0k_L#54nHn,4*4[+.I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+24dRR<=F_k0L4k#n,5H4[n*+24dRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*4[+c<2R=kRF0k_L#54nHn,4*4[+cI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+246RR<=F_k0L4k#n,5H4[n*+246RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*4[+n<2R=NRbs$H0_#Lk4Hn5,[.*2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[4R(2<b=RN0sH$k_L#54nH*,.[2+4RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRMRC8CRoMNCs0zCRc
.;RRRRRRRRCRM8oCCMsCN0Rgzd;R
RRMRC8CRoMNCs0zCRd
U;
RSRR-R-RMtCC0sNCER0CqR)vCRODRD#NRM8#CCDOD0RFOoHRsVFRv)qA_4n1_dn1
dnSUzdNRR:H5VROHEFOIC_HE80Rd=Rno2RCsMCN
0CSR--VRHGVRFsODNDRU4dUR(,#CCDOF0RVsR0HN#00MCRFL0RCoHMRosCHC#0s
C8SRRRRzRRO:E	RRHV58N8s8IH0>ERRRg2oCCMsCN0
RSSRkRRO:D	RFbsO#C#5iBp2S
SSCRLo
HMSRSSRRHV5iBp'CCPMN0RMB8Rp=iRR''42ER0CSM
SRSRRNRs8_8ss5CoNs88I0H8ER-48MFI0gFR2=R<R7q7)85N8HsI8-0E4FR8IFM0R;g2
SSSRMRC8VRH;S
SS8CMRFbsO#C#;S
SRMRC8CRoMNCs0zCRO;E	
RSRRdRzg:NRRsVFRHHRM8R5CEb0_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNC-
S-VRQR85N8HsI8R0E>2RgRCMC8FR0RCOsNR0CI0sHCMRCNCLDR8NMR0FkbRk0CLMND#CRCODC0FRDo
HOSzSScRjN:VRHR85N8HsI8R0E>2RgRMoCC0sNC-
S-HRVGFRVsNROD4DRd(UU,CR#D0CORRFV0#sH0CN0R0MFRHLCMsoRC#oH0CCs8S
SSRRRR0Fk_5CMH<2R=4R''ERIC5MRs8N8sC_so85N8HsI8-0E4FR8IFM0RRg2=2RHR#CDCjR''S;
SISSsC0_M25HRR<=WI RERCM5_N8s5CoNs88I0H8ER-48MFI0gFR2RR=HC2RDR#C';j'
SSSCRM8oCCMsCN0RjzcNS;
-Q-RVNR58I8sHE80RR<=gM2RFsRIHR0CCLMNDFCRskRF00bkRNCMLRDC#CCDOD0RFOoHRCMC8
C8SzSScR4N:VRHR85N8HsI8R0E<g=R2CRoMNCs0SC
SFSSkC0_M25HRR<=';4'
SSSS0Is_5CMH<2R= RW;S
SS8CMRMoCC0sNCcRz4
N;SR--tCCMsCN0RC0ERv)qRDOCDN#RM08Rs#H-0CN0#S
SS.zcNRR:VRFs[MRHRH5I8_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
RRRRRRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVAv)q_.64X7d.RD:RNDLCRRH#";W"
RRRRRRRRRRRRRRRRoLCHSM
SASS)_qv6X4.dR.7:qR)vnA4_n1d_n1d
RRRRRRRRRRRRRRRRbRRFRs0lRNb5q7QRR=>HsM_Cdo5n+*[d84RF0IMFnRd*,[2R7q7)=qR>FRDIN_I858sUFR8IFM0R,j2RS
SSQS7A>R=Rj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjj,j"R7q7)=AR>FRDIN_s858sUFR8IFM0R,j2
SSSSq hRR=>',4'R)11q>R=R''j, RWq>R=R0Is_5CMHR2,BqpiRR=>B,piRA hRR=>',4'R)11A>R=R''j, RWA>R=R''j,pRBi=AR>pRBiS,
S7SSm=qR>bRFCRM,75mAdR42=F>RkL0_k.#d5dH,.+*[d,42RA7m52djRR=>F_k0Ldk#.,5Hd[.*+2dj,S
SSmS7Ag5.2>R=R0Fk_#LkdH.5,*d.[g+.27,Rm.A5U=2R>kRF0k_L#5d.H.,d*.[+UR2,75mA.R(2=F>RkL0_k.#d5dH,.+*[.,(2
SSSSA7m52.nRR=>F_k0Ldk#.,5Hd[.*+2.n,mR7A65.2>R=R0Fk_#LkdH.5,*d.[6+.27,Rm.A5c=2R>kRF0k_L#5d.H.,d*.[+c
2,SSSS75mA.Rd2=F>RkL0_k.#d5dH,.+*[.,d2RA7m52..RR=>F_k0Ldk#.,5Hd[.*+2..,mR7A45.2>R=R0Fk_#LkdH.5,*d.[4+.2S,
S7SSm.A5j=2R>kRF0k_L#5d.H.,d*.[+jR2,75mA4Rg2=F>RkL0_k.#d5dH,.+*[4,g2RA7m524URR=>F_k0Ldk#.,5Hd[.*+24U,S
SSmS7A(542>R=R0Fk_#LkdH.5,*d.[(+427,Rm4A5n=2R>kRF0k_L#5d.H.,d*4[+nR2,75mA4R62=F>RkL0_k.#d5dH,.+*[4,62
SSSSA7m524cRR=>F_k0Ldk#.,5Hd[.*+24c,mR7Ad542>R=R0Fk_#LkdH.5,*d.[d+427,Rm4A5.=2R>kRF0k_L#5d.H.,d*4[+.R2,
SSSSA7m5244RR=>F_k0Ldk#.,5Hd[.*+244,mR7Aj542>R=R0Fk_#LkdH.5,*d.[j+427,RmgA52>R=R0Fk_#LkdH.5,*d.[2+g,SR
S7SSmUA52>R=R0Fk_#LkdH.5,*d.[2+U,mR7A25(RR=>F_k0Ldk#.,5Hd[.*+,(2RA7m5Rn2=F>RkL0_k.#d5dH,.+*[nR2,
SSSSA7m5R62=F>RkL0_k.#d5dH,.+*[6R2,75mAc=2R>kRF0k_L#5d.H.,d*c[+27,RmdA52>R=R0Fk_#LkdH.5,*d.[2+d,SR
S7SSm.A52>R=R0Fk_#LkdH.5,*d.[2+.,mR7A254RR=>F_k0Ldk#.,5Hd[.*+,42RA7m5Rj2=F>RkL0_k.#d5dH,.2*[,RR
RRRRRRRRRRRRRRRRRRRRRRRRR7RRQRuq=H>RMC_son5d*d[+6FR8IFM0R*dn[.+d27,RQRuA=">Rjjjj"7,RmRuq=F>Rb,CMRu7mA25dRR=>bHNs0L$_k.#d5cH,*d[+2R,
RRRRRRRRRRRRRRRRRRRRRRRRR7RRm5uA.=2R>NRbs$H0_#LkdH.5,[c*+,.2Ru7mA254RR=>bHNs0L$_k.#d5cH,*4[+27,Rm5uAj=2R>NRbs$H0_#LkdH.5,[c*2
2;RRRRRRRRRRRRRRRRF_k0s5Cod[n*2=R<R0Fk_#LkdH.5,*d.[I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cod[n*+R42<F=RkL0_k.#d5dH,.+*[4I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cod[n*+R.2<F=RkL0_k.#d5dH,.+*[.I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cod[n*+Rd2<F=RkL0_k.#d5dH,.+*[dI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cod[n*+Rc2<F=RkL0_k.#d5dH,.+*[cI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cod[n*+R62<F=RkL0_k.#d5dH,.+*[6I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cod[n*+Rn2<F=RkL0_k.#d5dH,.+*[nI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cod[n*+R(2<F=RkL0_k.#d5dH,.+*[(I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cod[n*+RU2<F=RkL0_k.#d5dH,.+*[UI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cod[n*+Rg2<F=RkL0_k.#d5dH,.+*[gI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cod[n*+24jRR<=F_k0Ldk#.,5Hd[.*+24jRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_son5d*4[+4<2R=kRF0k_L#5d.H.,d*4[+4I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cod[n*+24.RR<=F_k0Ldk#.,5Hd[.*+24.RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_son5d*4[+d<2R=kRF0k_L#5d.H.,d*4[+dI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cod[n*+24cRR<=F_k0Ldk#.,5Hd[.*+24cRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_son5d*4[+6<2R=kRF0k_L#5d.H.,d*4[+6I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cod[n*+24nRR<=F_k0Ldk#.,5Hd[.*+24nRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_son5d*4[+(<2R=kRF0k_L#5d.H.,d*4[+(I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cod[n*+24URR<=F_k0Ldk#.,5Hd[.*+24URCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_son5d*4[+g<2R=kRF0k_L#5d.H.,d*4[+gI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cod[n*+2.jRR<=F_k0Ldk#.,5Hd[.*+2.jRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_son5d*.[+4<2R=kRF0k_L#5d.H.,d*.[+4I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cod[n*+2..RR<=F_k0Ldk#.,5Hd[.*+2..RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_son5d*.[+d<2R=kRF0k_L#5d.H.,d*.[+dI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cod[n*+2.cRR<=F_k0Ldk#.,5Hd[.*+2.cRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_son5d*.[+6<2R=kRF0k_L#5d.H.,d*.[+6I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cod[n*+2.nRR<=F_k0Ldk#.,5Hd[.*+2.nRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_son5d*.[+(<2R=kRF0k_L#5d.H.,d*.[+(I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cod[n*+2.URR<=F_k0Ldk#.,5Hd[.*+2.URCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_son5d*.[+g<2R=kRF0k_L#5d.H.,d*.[+gI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cod[n*+2djRR<=F_k0Ldk#.,5Hd[.*+2djRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_son5d*d[+4<2R=kRF0k_L#5d.H.,d*d[+4I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cod[n*+2d.RR<=bHNs0L$_k.#d5cH,*R[2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*dn[d+d2=R<RsbNH_0$Ldk#.,5Hc+*[4I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cod[n*+2dcRR<=bHNs0L$_k.#d5cH,*.[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cdo5n+*[dR62<b=RN0sH$k_L#5d.H*,c[2+dRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRMRC8CRoMNCs0zCRc;.N
RRRRRRRR8CMRMoCC0sNCdRzg
N;RRRRCRM8oCCMsCN0RUzdNR;
R8CMRMoCC0sNCcRzdR;
Rczc:VRHRF5M08RN8ss_CRo2oCCMsCN0RR--oCCMsCN0RD#CCRO0s
NlRRRR-Q-RV8RN8HsI8R0E<RR(NH##o'MRj0'RFMRkk8#CR0LH#R
RRjRzRRR:H5VRNs88I0H8ERR=4o2RCsMCN
0CRRRRRRRRD_FINs88RR<="jjjj"jjR#&R__N8s5Coj
2;RRRRCRM8oCCMsCN0R;zj
RRRRRz4RH:RVNR58I8sHE80R.=R2CRoMNCs0RC
RRRRRDRRFNI_8R8s<"=Rjjjjj&"RRN#_8C_soR548MFI0jFR2R;
RCRRMo8RCsMCNR0Cz
4;RRRRzR.R:VRHR85N8HsI8R0E=2RdRMoCC0sNCR
RRRRRRFRDI8_N8<sR=jR"j"jjR#&R__N8s5Co.FR8IFM0R;j2
RRRR8CMRMoCC0sNC.Rz;R
RRdRzRRR:H5VRNs88I0H8ERR=co2RCsMCN
0CRRRRRRRRD_FINs88RR<="jjj"RR&#8_N_osC58dRF0IMF2Rj;R
RRMRC8CRoMNCs0zCRdS;
z:cSRRHV58N8s8IH0=ERRR62oCCMsCN0
DSSFNI_8R8s<"=RjRj"&_R#Ns8_Cco5RI8FMR0Fj
2;S8CMRMoCC0sNCcRz;z
S6RS:H5VRNs88I0H8ERR=no2RCsMCN
0CSFSDI8_N8<sR=jR''RR&#8_N_osC586RF0IMF2Rj;R
RRMRC8CRoMNCs0zCR6R;
RzRRn:RRRRHV58N8s8IH0>ERRRn2oCCMsCN0
RRRRRRRRIDF_8N8s=R<RN#_8C_soR5n8MFI0jFR2R;
RCRRMo8RCsMCNR0Cz
n;
RRRRR--Q5VR8_HMs2CoRosCHC#0sQR7h#RkHRMoB
piRRRRzR(R:VRHRH58MC_soo2RCsMCN
0CRRRRRRRRbOsFCR##5iBp,QR7hL2RCMoH
RRRRRRRRRRRRRHV5iBpR'=R4N'RMB8RpCi'P0CM2ER0CRM
RRRRRRRRRRRRR#RR__HMsRCo<7=RQ
h;RRRRRRRRRRRRCRM8H
V;RRRRRRRRCRM8bOsFC;##
RRRR8CMRMoCC0sNC(Rz;R
RRURzRRR:H5VRMRF08_HMs2CoRMoCC0sNCR
RRRRRRRRRR_R#HsM_C<oR=QR7hR;
RCRRMo8RCsMCNR0Cz
U;
RRRRR--Q5VR80Fk_osC2CRso0H#C7sRmRzakM#HoBRmpRi
RzRRg:RRRRHV5k8F0C_soo2RCsMCN
0CRRRRRRRRbOsFCR##5pmBiF,Rks0_CRo2LHCoMR
RRRRRRRRRRVRHRB5mp=iRR''4R8NMRpmBiP'CC2M0RC0EMR
RRRRRRRRRRRRRRmR7z<aR=_R#F_k0s;Co
RRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMRFbsO#C#;R
RRMRC8CRoMNCs0zCRgR;
RzRR4RjR:VRHRF5M0FR8ks0_CRo2oCCMsCN0
RRRRRRRRRRRRz7ma=R<RF#_ks0_C
o;RRRRCRM8oCCMsCN0Rjz4;R

R-RR-VRQR85N8ss_CRo2sHCo#s0CR7q7)#RkHRMoB
piRRRRzR44RH:RVNR58_8ss2CoRMoCC0sNCR
RRRRRRsRbF#OC#BR5pRi,q)772CRLo
HMRRRRRRRRRRRRH5VRBRpi=4R''MRN8pRBiP'CC2M0RC0EMR
RRRRRRRRRRRRRR_R#Ns8_C<oR=7Rq7N)58I8sHE80-84RF0IMF2Rj;R
RRRRRRRRRRMRC8VRH;R
RRRRRRMRC8sRbF#OC#R;
RCRRMo8RCsMCNR0Cz;44
RRRR.z4RH:RVMR5FN0R8_8ss2CoRMoCC0sNCR
RRRRRRRRRR_R#Ns8_C<oR=7Rq7
);RRRRCRM8oCCMsCN0R.z4;R
RRRRRRRR
R-RR-CRtMNCs00CRE)CRqOvRC#DDR8NMRD#CCRO0DHFoOR
RR4RzdRR:VRFsHMRHRk5MlC_OD4D_.-URRR428MFI0jFRRMoCC0sNCR
RR-R-RRQV58N8s8IH0>ERRR62M8CCRR0FONsC0ICRsCH0RNCMLRDCNRM8Fbk0kC0RMDNLCCR#D0CORoDFHRO
RRRRRzRR4:cRRRHV58N8s8IH0>ERRR(2oCCMsCN0
RRRRRRRRRRRRRRRRF#_kC0_M25HRR<='R4'IMECR_5#Ns8_CNo58I8sHE80-84RF0IMF2R(RH=R2DRC#'CRj
';RRRRRRRRRRRRRRRR#s_I0M_C5RH2<W=R ERIC5MR#8_N_osC58N8s8IH04E-RI8FMR0F(=2RRRH2CCD#R''j;R
RRRRRRMRC8CRoMNCs0zCR4
c;RRRR-Q-RVNR58I8sHE80RR<=6M2RFsRIHR0CCLMNDFCRskRF00bkRNCMLRDC#CCDOD0RFOoHRCMC8
C8RRRRRRRRzR46:VRHR85N8HsI8R0E<(=R2CRoMNCs0RC
RRRRRRRRRRRRR#RR_0Fk_5CMH<2R=4R''R;
RRRRRRRRRRRRR#RR_0Is_5CMH<2R= RW;R
RRRRRRMRC8CRoMNCs0zCR4
6;RRRR-t-RCsMCNR0C0REC)RqvODCD#MRN8sR0H0-#N#0C
RRRRRRRRnz4RV:RF[sRRRHM58IH0-ERRR428MFI0jFRRMoCC0sNCR
RRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqz)vU4.RD:RNDLCRRH#"a11"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloHC5*U4.2RR&"RW"&MRH0CCosl'HN5oC[&2RR"" RH&RMo0CCHs'lCNo50oC_8CM_b8C05E5H2+4*U4.,CR8b20E2RR&"RX"&MRH0CCosl'HN5oC[2+4;R
RRRRRRRRRRCRLo
HMRRRRRRRRRRRRzv)q4R.U:)RXq.v4U1X4RR
RRRRRRRRRRRRRRFRbsl0RN5bR7>R=RH#_MC_so25[,jRqRR=>D_FINs885,j2RRq4=D>RFNI_858s4R2,q=.R>FRDI8_N8.s52R,
RRRRRRRRRRRRRRRRRRRRRRRRRRqd=D>RFNI_858sdR2,q=cR>FRDI8_N8cs52q,R6>R=RIDF_8N8s256,nRqRR=>D_FINs885,n2
SSSSRSSRRW =#>R_0Is_5CMHR2,WiBpRR=>B,piR=mR>kRF0k_L#._4U,5H[;22
RRRRRRRRRRRRRRRRF#_ks0_C[o52=R<R0Fk_#Lk_U4.5[H,2ERIC5MR#k_F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRR8CMRMoCC0sNC4RznR;
RRRRCRM8oCCMsCN0Rdz4;RRRRRRRRRRRRR
RRRRR
RRRRR--tCCMsCN0R4NRnFRIs88RCRCb)RqvODCDRRHVNsbbFHbsNR0CRRRRRRRRRRRRRRR
RzRR4:(RRRHV5lMk_DOCDc_nR4=R2CRoMNCs0RC
R-RR-VRQR85N8HsI8R0E>2R(RCMC8FR0RCOsNR0CI0sHCMRCNCLDR8NMR0FkbRk0CLMND#CRCODC0FRDo
HORRRRRRRRzN4URH:RVNR58I8sHE80R(>R2CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_Mc_nRR<='R4'IMECR#55__N8s5CoNs88I0H8ER-48MFI0(FR2RR=M_klODCD_U4.2MRN8#R5__N8s5Con=2RR''j2C2RDR#C';j'
RRRRRRRRRRRRRRRR0Is__CMn<cR= RWRCIEM5R5#8_N_osC58N8s8IH04E-RI8FMR0F(=2RRlMk_DOCD._4UN2RM58R#8_N_osC5Rn2=jR''R22CCD#R''j;R
RRRRRRMRC8CRoMNCs0zCR4;UN
RRRRRRRRUz4LRR:H5VRNs88I0H8ERR=(MRN8kRMlC_OD4D_.=URRRj2oCCMsCN0
RRRRRRRRRRRRRRRR0Fk__CMn<cR=4R''ERIC5MR5N#_8C_so25nR'=Rj2'2R#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_Mc_nRR<=WI RERCM5_5#Ns8_Cno52RR='2j'2DRC#'CRj
';RRRRRRRRCRM8oCCMsCN0RUz4LR;
R-RR-VRQR85N8HsI8R0E<6=R2FRMRHIs0CCRMDNLCsRFR0FkbRk0CLMND#CRCODC0FRDoRHOM8CCCR8
RRRRRzRR4:gRRRHV58N8s8IH0<ER=2RnRMoCC0sNCR
RRRRRRRRRRRRRRkRF0M_C_Rnc<'=R4
';RRRRRRRRRRRRRRRRI_s0CnM_c=R<R;W 
RRRRRRRR8CMRMoCC0sNC4RzgR;
R-RR-CRtMNCs00CRE)CRqOvRCRDDNRM80-sH#00NCR
SRzRRO_E	.RR:H5VR#H_I8_0ENNss$c_n5R42>2RjRMoCC0sNCR
RRRRRR.RzjRR:VRFs[MRHR_5#I0H8Es_Ns_N$n4c52RR-482RF0IMFRRjoCCMsCN0
RRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVzv)qn:cRRLDNCHDR#1R"1Ra"&MRH0CCosl'HN5oCI0H8E&2RR""7RH&RMo0CCHs'lCNo5lMk_DOCD._4U.*4U&2RR""WRH&RMo0CCHs'lCNo58IH0-ERR[.*R.-R2RR&"R "&MRH0CCosl'HN5oCo_C0C_M880CbEk5MlC_OD4D_.4U*.+URR,ncRb8C02E2R"&RX&"RR0HMCsoC'NHloIC5HE80R.-R*;[2
RRRRRRRRRRRRoLCHRM
RRRRRRRRRzRR)nqvcRR:Xv)qn.cX1RR
RRRRRRRRRRRRRbRRFRs0lRNb5R74=#>R__HMs5CoI0H8E*-.[2-4,jR7RR=>#M_H_osC58IH0.E-*.[-2q,Rj>R=RIDF_8N8s25j,4RqRR=>D_FINs885,42RRq.=D>RFNI_858s.
2,RRRRRRRRRRRRRRRRRRRRRRRRRdRqRR=>D_FINs885,d2RRqc=D>RFNI_858scR2,q=6R>FRDI8_N86s52S,
SSSSSWRR >R=R0Is__CMnRc,WiBpRR=>B,piRRm4=F>RkL0_kn#_ck5MlC_ODnD_cH,I8-0E.-*[4R2,m=jR>kRF0k_L#c_n5lMk_DOCDc_n,8IH0.E-*.[-2
2;RRRRRRRRRRRRRRRR#k_F0C_soH5I8-0E.-*[4<2R=kRF0k_L#c_n5lMk_DOCDc_n,8IH0.E-*4[-2ERIC5MRF_k0CnM_cRR='24'R#CDCZR''R;
RRRRRRRRRRRRR#RR_0Fk_osC58IH0.E-*.[-2=R<R0Fk_#Lk_5ncM_klODCD_,ncI0H8E*-.[2-.RCIEMFR5kC0_Mc_nR'=R4R'2CCD#R''Z;R
RRRRRRCRRMo8RCsMCNR0Cz;.j
RSSCRM8oCCMsCN0REzO	;_.
RSSz	OE_:4RRRHV5I#_HE80_sNsNn$_c25jRj>R2CRoMNCs0RC
RRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)RzqcvnRD:RNDLCRRH#"a11"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloMC5kOl_C_DD4*.U42.UR"&RW&"RR0HMCsoC'NHloIC5HE80R.-R*I#_HE80_sNsNn$_c254R4-R2RR&"R "&MRH0CCosl'HN5oCo_C0C_M880CbEk5MlC_OD4D_.4U*.+URR,ncRb8C02E2R"&RX&"RR0HMCsoC'NHloIC5HE80R.-R*I#_HE80_sNsNn$_c2542R;
RRRRRRRRRLRRCMoH
RRRRRRRRRRRRqz)vRnc:qR)vXnc4
1RRRRRRRRRRRRRRRRRb0FsRblNRR57=#>R__HMs5CoI0H8E*-.#H_I8_0ENNss$c_n5-424R2,q=jR>FRDI8_N8js52q,R4>R=RIDF_8N8s254,.RqRR=>D_FINs885,.2
RRRRRRRRRRRRRRRRRRRRRRRRqRRd>R=RIDF_8N8s25d,cRqRR=>D_FINs885,c2RRq6=D>RFNI_858s6
2,SSSSSRSRW= R>sRI0M_C_,ncRpWBi>R=RiBp,RRm=F>RkL0_kn#_ck5MlC_ODnD_cH,I8-0E._*#I0H8Es_Ns_N$n4c522-42R;
RRRRRRRRRRRRR#RR_0Fk_osC58IH0.E-*I#_HE80_sNsNn$_c254-R42<F=RkL0_kn#_ck5MlC_ODnD_cH,I8-0E._*#I0H8Es_Ns_N$n4c522-4RCIEMFR5kC0_Mc_nR'=R4R'2CCD#R''Z;R
RRRRRRCRRMo8RCsMCNR0Cz	OE_
4;SRRRRMRC8CRoMNCs0zCR4R(;RRRRRRRRRR

R-RR-CRtMNCs0NCRRR4nI8FsRC8CbqR)vCRODHDRVbRNbbsFs0HNCRRRRRRRRRRRRRRR
RRRR4z.RH:RVMR5kOl_C_DDd=.RRR42oCCMsCN0
RRRRR--Q5VRNs88I0H8ERR>6M2RCRC80OFRs0CNCsRIHR0CCLMNDNCRMF8Rkk0b0MRCNCLDRD#CCRO0DHFoOR
RRRRRR.Rz.:NRRRHV58N8s8IH0>ERRN(RMM8RkOl_C_DDn=cRRR42oCCMsCN0
RRRRRRRRRRRRRRRR0Fk__CMd<.R=4R''ERIC5MR5N#_8C_so85N8HsI8-0E4FR8IFM0RR(2=kRMlC_OD4D_.RU2NRM85N#_8C_so25nR'=R4R'2NRM85N#_8C_so256R'=Rj2'2R#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_M._dRR<=WI RERCM5_5#Ns8_CNo58I8sHE80-84RF0IMF2R(RM=RkOl_C_DD42.UR8NMR_5#Ns8_Cno52RR='24'R8NMR_5#Ns8_C6o52RR='2j'2DRC#'CRj
';RRRRRRRRCRM8oCCMsCN0R.z.NR;
RRRRRzRR.R.L:VRHR85N8HsI8R0E>RR(NRM8M_klODCD_Rnc/4=R2CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_M._dRR<='R4'IMECR#55__N8s5CoNs88I0H8ER-48MFI0(FR2RR=M_klODCD_U4.2MRN8#R5__N8s5Con=2RR''j2MRN8#R5__N8s5Co6=2RR''j2C2RDR#C';j'
RRRRRRRRRRRRRRRR0Is__CMd<.R= RWRCIEM5R5#8_N_osC58N8s8IH04E-RI8FMR0F(=2RRlMk_DOCD._4UN2RM58R#8_N_osC5Rn2=jR''N2RM58R#8_N_osC5R62=jR''R22CCD#R''j;R
RRRRRRMRC8CRoMNCs0zCR.;.L
RRRRRRRR.z.ORR:H5VRNs88I0H8ERR=(MRN8kRMlC_ODnD_cRR=4o2RCsMCN
0CRRRRRRRRRRRRRRRRF_k0CdM_.=R<R''4RCIEM5R5#8_N_osC5Rn2=4R''N2RM58R#8_N_osC5R62=jR''R22CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C_Rd.<W=R ERIC5MR5N#_8C_so25nR'=R4R'2NRM85N#_8C_so256R'=Rj2'2R#CDCjR''R;
RRRRRCRRMo8RCsMCNR0CzO..;R
RRRRRR.Rz.:8RRRHV58N8s8IH0=ERRNnRMM8RkOl_C_DDn/cR=2R4RMoCC0sNCR
RRRRRRRRRRRRRRkRF0M_C_Rd.<'=R4I'RERCM5_5#Ns8_CNo58I8sHE80-84RF0IMF2R6RM=RkOl_C_DDn2c2R#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_M._dRR<=WI RERCM5_5#Ns8_CNo58I8sHE80-84RF0IMF2R6RM=RkOl_C_DDn2c2R#CDCjR''R;
RRRRRCRRMo8RCsMCNR0Cz8..;R
RR-R-RRQV58N8s8IH0<ER=2R6RRMFI0sHCMRCNCLDRRFsFbk0kC0RMDNLCCR#D0CORoDFHMORCCC88R
RRRRRR.RzdRR:H5VRNs88I0H8E=R<RR62oCCMsCN0
RRRRRRRRRRRRRRRR0Fk__CMd<.R=4R''R;
RRRRRRRRRRRRRIRRsC0_M._dRR<=W
 ;RRRRRRRRCRM8oCCMsCN0Rdz.;R
RR-R-RMtCC0sNCER0CqR)vCRODNDRM08Rs#H-0CN0
RSRRORzEU	_RH:RV#R5_8IH0NE_s$sN5Rd2>2RjRMoCC0sNCS
Sz	OE_6DCRH:RVIR5HE80RR>=U_*#I0H8Es_Ns5N$dN2RMI8RHE80RR>=Uo2RCsMCN
0CRRRRRRRRRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FzVR)dqv.RR:DCNLD#RHR1"1a&"RR0HMCsoC'NHloIC5HE802RR&"R7"&MRH0CCosl'HN5oCM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*c&2RR""WRH&RMo0CCHs'lCNo58IH0-ERRLD#_8IH0RE2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50EM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*cRR+dR.,80CbER22&XR""RR&HCM0o'CsHolNCH5I8R0E-#RDLH_I8R0E+2RU;R
RRRRRRRRRRRRRRRRRRCRLo
HMSRSRR)Rzq.vdRX:R)dqv.1XU
SSSRRRRb0FsRblNRR57=b>RN#85__HMs5CoI0H8ER-48MFI0IFRHE80-LD#_8IH0,E2RRU,D_#LI0H8E2-4,jRqRR=>D_FINs885,j2
SSSSRSSRRq4=D>RFNI_858s4R2,q=.R>FRDI8_N8.s52q,Rd>R=RIDF_8N8s25d,cRqRR=>D_FINs885,c2RRW =I>RsC0_M._d,BRWp=iR>pRBiS,
SSSSSmRRRR=>0_lbU._d52j2;S
SS#SN#MHoRV:RFHsR[MRHR8IH04E-RI8FMR0FI0H8E#-DLH_I8R0EoCCMsCN0
SSSSFRRkL0_kd#_.k5MlC_ODdD_.[,H2=R<Rb0l_dU_.25j5-H[I0H8E#+DLH_I820E;R
RRRRRRRRRRRRRRRRR#k_F0C_so[5H2=R<R0Fk_#Lk_5d.M_klODCD_,d.HR[2IMECRk5F0M_C_Rd.=4R''C2RDR#C';Z'
SSSS8CMRMoCC0sNC#RN#MHo;R
RRRRRRRRRR.RzURR:VRFs[MRHRI#_HE80_sNsNd$52R-48MFI04FRRMoCC0sNCR
RRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FzVR)dqv.RR:DCNLD#RHR1"1a&"RR0HMCsoC'NHloIC5HE802RR&"R7"&MRH0CCosl'HN5oCM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*c&2RR""WRH&RMo0CCHs'lCNo58IH0-ERRLD#_8IH0-ERRU[*2RR&"R "&MRH0CCosl'HN5oCo_C0C_M880CbEk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*Rnc+.Rd,CR8b20E2RR&"RX"&MRH0CCosl'HN5oCI0H8ERR-D_#LI0H8ERR-54[-22*U;R
RRRRRRRRRRRRRLHCoMR
RRRRRRRRRRRRRzv)qd:.RRqX)vXd.U
1RRRRRRRRRRRRRRRRRb0FsRblNRR57=#>R__HMs5CoI0H8E#-DLH_I8-0EU+*[(FR8IFM0R8IH0DE-#IL_HE80-[U*2q,Rj>R=RIDF_8N8s25j,4RqRR=>D_FINs885,42RRq.=D>RFNI_858s.
2,RRRRRRRRRRRRRRRRRRRRRRRRRdRqRR=>D_FINs885,d2RRqc=D>RFNI_858scR2,W= R>sRI0M_C_,d.RpWBi>R=RiBp,RRm=0>RlUb__5d.[;22
SSSRRRRNH##o:MRRsVFRRH[H(MRRI8FMR0FjCRoMNCs0SC
SRSSR0Fk_#Lk_5d.M_klODCD_,d.I0H8E#-DLH_I8-0EU+*[HR[2<0=RlUb__5d.[H25[
2;RRRRRRRRRRRRRRRRR_R#F_k0s5CoI0H8E#-DLH_I8-0EU+*[HR[2<F=RkL0_kd#_.k5MlC_ODdD_.H,I8-0ED_#LI0H8E*-U[[+H2ERIC5MRF_k0CdM_.RR='24'R#CDCZR''R;
RRRRRRRRRRRRRCRRMo8RCsMCNR0CNH##o
M;RRRRRRRRRRRRCRM8oCCMsCN0RUz.;S
SCRM8oCCMsCN0REzO	C_D6S;
SEzO	0_o6RR:H5VRI0H8E=R>RNURMI8RHE80R8lFR>UR=2R6RMoCC0sNCR
RRRRRRRRRRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqz)vRd.:NRDLRCDH"#R1"1aRH&RMo0CCHs'lCNo58IH0RE2&7R""RR&HCM0o'CsHolNCk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*2ncR"&RW&"RR0HMCsoC'NHloIC5HE80RD-R#IL_HE802RR&"R "&MRH0CCosl'HN5oCo_C0C_M880CbEk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*Rnc+.Rd,CR8b20E2RR&"RX"&MRH0CCosl'HN5oCI0H8ERR-D_#LI0H8ERR+U
2;RRRRRRRRRRRRRRRRRRRRLHCoMS
SRRRRzv)qd:.RRqX)vXd.US1
SRSRRFRbsl0RN5bR7>R=R8bN5H#_MC_soH5I8-0E4FR8IFM0R8IH0DE-#IL_HE802U,R,#RDLH_I8-0E4R2,q=jR>FRDI8_N8js52S,
SSSSSqRR4>R=RIDF_8N8s254,.RqRR=>D_FINs885,.2RRqd=D>RFNI_858sdR2,q=cR>FRDI8_N8cs52W,R >R=R0Is__CMdR.,WiBpRR=>B,pi
SSSSRSSR=mR>lR0b__Ud#.5_8IH0NE_s$sN5-d24;22
SSSS#N#HRoM:FRVs[RHRRHMI0H8ER-48MFI0IFRHE80-LD#_8IH0oERCsMCN
0CSSSSRkRF0k_L#._d5lMk_DOCD._d,2H[RR<=0_lbU._d5I#_HE80_sNsNd$522-45-H[I0H8E#+DLH_I820E;R
RRRRRRRRRRRRRRRRR#k_F0C_so[5H2=R<R0Fk_#Lk_5d.M_klODCD_,d.HR[2IMECRk5F0M_C_Rd.=4R''C2RDR#C';Z'
SSSS8CMRMoCC0sNC#RN#MHo;R
RRRRRRRRRR.RzURR:VRFs[MRHRI#_HE80_sNsNd$52R-.8MFI0jFRRMoCC0sNCR
RRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FzVR)dqv.RR:DCNLD#RHR1"1a&"RR0HMCsoC'NHloIC5HE802RR&"R7"&MRH0CCosl'HN5oCM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*c&2RR""WRH&RMo0CCHs'lCNo5U[*2RR&"R "&MRH0CCosl'HN5oCo_C0C_M880CbEk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*Rnc+.Rd,CR8b20E2RR&"RX"&MRH0CCosl'HN5oC54[+22*U;R
RRRRRRRRRRRRRLHCoMR
RRRRRRRRRRRRRzv)qd:.RRqX)vXd.U
1RRRRRRRRRRRRRRRRRb0FsRblNRR57=#>R__HMs5CoU+*[(FR8IFM0R[U*2q,Rj>R=RIDF_8N8s25j,4RqRR=>D_FINs885,42RRq.=D>RFNI_858s.
2,RRRRRRRRRRRRRRRRRRRRRRRRRdRqRR=>D_FINs885,d2RRqc=D>RFNI_858scR2,W= R>sRI0M_C_,d.RpWBi>R=RiBp,RRm=0>RlUb__5d.[;22
SSSS#N#HRoM:FRVs[RHRRHM(FR8IFM0RojRCsMCN
0CSSSSRkRF0k_L#._d5lMk_DOCD._d,[U*+2H[RR<=0_lbU._d55[2H;[2
RRRRRRRRRRRRRRRR#RR_0Fk_osC5[U*+2H[RR<=F_k0L_k#dM.5kOl_C_DDdU.,*H[+[I2RERCM50Fk__CMd=.RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRCRM8oCCMsCN0R#N#H;oM
RRRRRRRRRRRR8CMRMoCC0sNC.RzUS;
S8CMRMoCC0sNCORzEo	_0
6;SOSzEM	_RH:RVIR5HE80RU<R2CRoMNCs0RC
RRRRRRRRRRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)Rzq.vdRD:RNDLCRRH#"a11"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloMC5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*n2RR&"RW"&MRH0CCosl'HN5oCj&2RR"" RH&RMo0CCHs'lCNo50oC_8CM_b8C0ME5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*nRd+R.8,RCEb02&2RR""XRH&RMo0CCHs'lCNo5;U2
RRRRRRRRRRRRRRRRRRRRoLCHSM
SRRRRqz)vRd.:)RXq.vdX
U1SRSSRbRRFRs0lRNb5=7R>NRb8_5#HsM_CIo5HE80-84RF0IMFHRI8-0ED_#LI0H8ER2,UD,R#IL_HE80-,42RRqj=D>RFNI_858sj
2,SSSSSRSRq=4R>FRDI8_N84s52q,R.>R=RIDF_8N8s25.,dRqRR=>D_FINs885,d2RRqc=D>RFNI_858scR2,W= R>sRI0M_C_,d.RpWBi>R=RiBp,S
SSSSSRRRm=0>RlUb__5d.j;22
SSSS#N#HRoM:FRVs[RHRRHMI0H8ER-48MFI0jFRRMoCC0sNCS
SSRSRF_k0L_k#dM.5kOl_C_DDdH.,[<2R=lR0b__Udj.52[5H2R;
RRRRRRRRRRRRRRRRRF#_ks0_CHo5[<2R=kRF0k_L#._d5lMk_DOCD._d,2H[RCIEMFR5kC0_M._dR'=R4R'2CCD#R''Z;S
SSMSC8CRoMNCs0NCR#o#HMS;
S8CMRMoCC0sNCORzEM	_;S
SCRM8oCCMsCN0REzO	;_U
zSSO_E	cRR:H5VR#H_I8_0ENNss$25.Rj>R2CRoMNCs0RC
RRRRRzRR.cc_RH:RVIR5HE80RR>=co2RCsMCN
0CRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FzVR)dqv.RR:DCNLD#RHR1"1a&"RR0HMCsoC'NHloIC5HE802RR&"R7"&MRH0CCosl'HN5oCM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*c&2RR""WRH&RMo0CCHs'lCNo5Rj2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50EM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*cRR+dR.,80CbER22&XR""RR&HCM0o'CsHolNC25c;R
RRRRRRRRRRCRLo
HMRRRRRRRRRRRRzv)qd:.RRqX)vXd.c
1RRRRRRRRRRRRRRRRRb0FsRblNRd57RR=>#M_H_osC5,d2RR7.=#>R__HMs5Co.R2,7=4R>_R#HsM_C4o527,Rj>R=RH#_MC_so25j,S
SSRRRRRRRRRRRRqRRj>R=RIDF_8N8s25j,4RqRR=>D_FINs885,42RRq.=D>RFNI_858s.
2,RRRRRRRRRRRRRRRRRRRRRRRRRdRqRR=>D_FINs885,d2RRqc=D>RFNI_858scR2,W= R>sRI0M_C_,d.RpWBi>R=RiBp,SR
SSSSSmRRd>R=R0Fk_#Lk_5d.M_klODCD_,d.dR2,m=.R>kRF0k_L#._d5lMk_DOCD._d,,.2
SSSSRSSRRm4=F>RkL0_kd#_.k5MlC_ODdD_.2,4,jRmRR=>F_k0L_k#dM.5kOl_C_DDdj.,2
2;RRRRRRRRRRRRRRRR#k_F0C_so25dRR<=F_k0L_k#dM.5kOl_C_DDdd.,2ERIC5MRF_k0CdM_.RR='24'R#CDCZR''R;
RRRRRRRRRRRRR#RR_0Fk_osC5R.2<F=RkL0_kd#_.k5MlC_ODdD_.2,.RCIEMFR5kC0_M._dR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRR_R#F_k0s5Co4<2R=kRF0k_L#._d5lMk_DOCD._d,R42IMECRk5F0M_C_Rd.=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRF#_ks0_Cjo52=R<R0Fk_#Lk_5d.M_klODCD_,d.jI2RERCM50Fk__CMd=.RR''42DRC#'CRZ
';RRRRRRRRCRM8oCCMsCN0Rcz._
c;RRRRRRRRz_.cdRR:H5VRI0H8ERR=do2RCsMCN
0CRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FzVR)dqv.RR:DCNLD#RHR1"1a&"RR0HMCsoC'NHloIC5HE802RR&"R7"&MRH0CCosl'HN5oCM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*c&2RR""WRH&RMo0CCHs'lCNo5Rj2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50EM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*cRR+dR.,80CbER22&XR""RR&HCM0o'CsHolNC25c;R
RRRRRRRRRRCRLo
HMRRRRRRRRRRRRzv)qd:.RRqX)vXd.c
1RRRRRRRRRRRRRRRRRb0FsRblNRd57RR=>',j'RR7.=#>R__HMs5Co.R2,7=4R>_R#HsM_C4o527,Rj>R=RH#_MC_so25j,S
SSRRRRRRRRRRRRqRRj>R=RIDF_8N8s25j,4RqRR=>D_FINs885,42RRq.=D>RFNI_858s.
2,RRRRRRRRRRRRRRRRRRRRRRRRRdRqRR=>D_FINs885,d2RRqc=D>RFNI_858scR2,W= R>sRI0M_C_,d.RpWBi>R=RiBp,SR
SSSSSmRRd>R=RCFbMm,R.>R=R0Fk_#Lk_5d.M_klODCD_,d..
2,SSSSSRSRm=4R>kRF0k_L#._d5lMk_DOCD._d,,42RRmj=F>RkL0_kd#_.k5MlC_ODdD_.2,j2R;
RRRRRRRRRRRRR#RR_0Fk_osC5R.2<F=RkL0_kd#_.k5MlC_ODdD_.2,.RCIEMFR5kC0_M._dR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRR_R#F_k0s5Co4<2R=kRF0k_L#._d5lMk_DOCD._d,R42IMECRk5F0M_C_Rd.=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRF#_ks0_Cjo52=R<R0Fk_#Lk_5d.M_klODCD_,d.jI2RERCM50Fk__CMd=.RR''42DRC#'CRZ
';RRRRRRRRCRM8oCCMsCN0Rcz._
d;SMSC8CRoMNCs0zCRO_E	cS;
SEzO	R_.:VRHR_5#I0H8Es_Ns5N$4>2RRRj2oCCMsCN0
RRRRRRRRcz.RV:RF[sRRRHM5I#_HE80_sNsN4$52RR-482RF0IMFRRjoCCMsCN0
RRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVzv)qd:.RRLDNCHDR#1R"1Ra"&MRH0CCosl'HN5oCI0H8E&2RR""7RH&RMo0CCHs'lCNo5lMk_DOCD._4U.*4URR+M_klODCD_*ncnRc2&WR""RR&HCM0o'CsHolNCH5I8-0EU_*#I0H8Es_Ns5N$d.2-*.[-2RR&"R "&MRH0CCosl'HN5oCo_C0C_M880CbEk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*Rnc+.Rd,CR8b20E2RR&"RX"&MRH0CCosl'HN5oCI0H8E*-U#H_I8_0ENNss$25d-[.*2R;
RRRRRRRRRLRRCMoH
RRRRRRRRRRRRqz)vRd.:qR)vXd..
1RRRRRRRRRRRRRRRRRb0FsRblNRj57RR=>#M_H_osC58IH0UE-*I#_HE80_sNsNd$52*-.[2-.,4R7RR=>#M_H_osC58IH0UE-*I#_HE80_sNsNd$52*-.[2-4,jRqRR=>D_FINs885,j2RRq4=D>RFNI_858s4R2,q=.R>FRDI8_N8.s52R,
RRRRRRRRRRRRRRRRRRRRRRRRRRqd=D>RFNI_858sdR2,q=cR>FRDI8_N8cs52W,R >R=R0Is__CMdR.,WiBpRR=>B,piRRmj=F>RkL0_kd#_.k5MlC_ODdD_.H,I8-0EU_*#I0H8Es_Ns5N$d.2-*.[-2S,
SSSSSmRR4>R=R0Fk_#Lk_5d.M_klODCD_,d.I0H8E*-U#H_I8_0ENNss$25d-[.*-242;R
RRRRRRRRRRRRRR_R#F_k0s5CoI0H8E*-U#H_I8_0ENNss$25d-[.*-R42<F=RkL0_kd#_.k5MlC_ODdD_.H,I8-0EU_*#I0H8Es_Ns5N$d.2-*4[-2ERIC5MRF_k0CdM_.RR='24'R#CDCZR''R;
RRRRRRRRRRRRR#RR_0Fk_osC58IH0UE-*I#_HE80_sNsNd$52*-.[2-.RR<=F_k0L_k#dM.5kOl_C_DDdI.,HE80-#U*_8IH0NE_s$sN5-d2.-*[.I2RERCM50Fk__CMd=.RR''42DRC#'CRZ
';RRRRRRRRCRM8oCCMsCN0Rcz.;S
SCRM8oCCMsCN0REzO	;_.
zSSO_E	4RR:H5VR#H_I8_0ENNss$25jRj>R2CRoMNCs0RC
RRRRRzRR.:cRRRHV58IH0lERFU8RR4=R2CRoMNCs0RC
RRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)Rzq.vdRD:RNDLCRRH#"a11"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloMC5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*n2RR&"RW"&MRH0CCosl'HN5oCj&2RR"" RH&RMo0CCHs'lCNo50oC_8CM_b8C0ME5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*nRd+R.8,RCEb02&2RR""XRH&RMo0CCHs'lCNo5;42
RRRRRRRRRRRRoLCHRM
RRRRRRRRRzRR)dqv.RR:)dqv.1X4RR
RRRRRRRRRRRRRRFRbsl0RN5bR7>R=RH#_MC_so25j,jRqRR=>D_FINs885,j2RRq4=D>RFNI_858s4R2,q=.R>FRDI8_N8.s52R,
RRRRRRRRRRRRRRRRRRRRRRRRRRqd=D>RFNI_858sdR2,q=cR>FRDI8_N8cs52W,R >R=R0Is__CMdR.,WiBpRR=>B,piR=mR>kRF0k_L#._d5lMk_DOCD._d,2j2;R
RRRRRRRRRRRRRR_R#F_k0s5Coj<2R=kRF0k_L#._d5lMk_DOCD._d,Rj2IMECRk5F0M_C_Rd.=4R''C2RDR#C';Z'
RRRRRRRR8CMRMoCC0sNC.RzcS;
S8CMRMoCC0sNCORzE4	_;R
RRMRC8CRoMNCs0zCR.R4;RRRRRRRRRR

R-RR-CRtMNCs0NCRRR4nI8FsRC8CbqR)vCRODHDRVbRNbbsFs0HNCRRRRRRRRRRRRRRR
RRRR6z.RH:RVMR5kOl_C_DD4=nRRR42oCCMsCN0
RRRRR--Q5VRNs88I0H8ERR>6M2RCRC80OFRs0CNCsRIHR0CCLMNDNCRMF8Rkk0b0MRCNCLDRD#CCRO0DHFoOR
RRRRRR.Rzn:NRRRHV58N8s8IH0>ERRN(RMM8RkOl_C_DDn=cRRN4RMM8RkOl_C_DDd=.RRR42oCCMsCN0
RRRRRRRRRRRRRRRR0Fk__CM4<nR=4R''ERIC5MR5N#_8C_so85N8HsI8-0E4FR8IFM0RR(2=kRMlC_OD4D_.RU2NRM85N#_8C_so25nR'=R4R'2NRM85N#_8C_so256R'=R4R'2NRM85N#_8C_so25cR'=Rj2'2R#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_Mn_4RR<=WI RERCM5_5#Ns8_CNo58I8sHE80-84RF0IMF2R(RM=RkOl_C_DD42.UR8NMR_5#Ns8_Cno52RR='24'R8NMR_5#Ns8_C6o52RR='24'R8NMR_5#Ns8_Cco52RR='2j'2DRC#'CRj
';RRRRRRRRCRM8oCCMsCN0Rnz.NR;
RRRRRzRR.RnL:VRHR85N8HsI8R0E>RR(NRM8M_klODCD_Rnc=RR4NRM8M_klODCD_Rd.=2RjRMoCC0sNCR
RRRRRRRRRRRRRRkRF0M_C_R4n<'=R4I'RERCM5_5#Ns8_CNo58I8sHE80-84RF0IMF2R(RM=RkOl_C_DD42.UR8NMR_5#Ns8_Cno52RR='24'R8NMR_5#Ns8_C6o52RR='2j'R8NMR_5#Ns8_Cco52RR='2j'2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0C4M_n=R<RRW IMECR#55__N8s5CoNs88I0H8ER-48MFI0(FR2RR=M_klODCD_U4.2MRN8#R5__N8s5Con=2RR''42MRN8#R5__N8s5Co6=2RR''j2MRN8#R5__N8s5Coc=2RR''j2C2RDR#C';j'
RRRRRRRR8CMRMoCC0sNC.Rzn
L;RRRRRRRRzO.nRH:RVNR58I8sHE80R(>RR8NMRlMk_DOCDc_nRj=RR8NMRlMk_DOCD._dR4=R2CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_Mn_4RR<='R4'IMECR#55__N8s5CoNs88I0H8ER-48MFI0(FR2RR=M_klODCD_U4.2MRN8#R5__N8s5Con=2RR''j2MRN8#R5__N8s5Co6=2RR''42MRN8#R5__N8s5Coc=2RR''j2C2RDR#C';j'
RRRRRRRRRRRRRRRR0Is__CM4<nR= RWRCIEM5R5#8_N_osC58N8s8IH04E-RI8FMR0F(=2RRlMk_DOCD._4UN2RM58R#8_N_osC5Rn2=jR''N2RM58R#8_N_osC5R62=4R''N2RM58R#8_N_osC5Rc2=jR''R22CCD#R''j;R
RRRRRRMRC8CRoMNCs0zCR.;nO
RRRRRRRRnz.8RR:H5VRNs88I0H8ERR>(MRN8kRMlC_ODnD_cRR=jMRN8kRMlC_ODdD_.RR=jo2RCsMCN
0CRRRRRRRRRRRRRRRRF_k0C4M_n=R<R''4RCIEM5R5#8_N_osC58N8s8IH04E-RI8FMR0F(=2RRlMk_DOCD._4UN2RM58R#8_N_osC5Rn2=jR''N2RM58R#8_N_osC5R62=jR''N2RM58R#8_N_osC5Rc2=jR''R22CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C_R4n<W=R ERIC5MR5N#_8C_so85N8HsI8-0E4FR8IFM0RR(2=kRMlC_OD4D_.RU2NRM85N#_8C_so25nR'=RjR'2NRM85N#_8C_so256R'=RjR'2NRM85N#_8C_so25cR'=Rj2'2R#CDCjR''R;
RRRRRCRRMo8RCsMCNR0Cz8.n;R
RRRRRR.Rzn:CRRRHV58N8s8IH0=ERRN(RMM8RkOl_C_DDn=cRRN4RMM8RkOl_C_DDd=.RRR42oCCMsCN0
RRRRRRRRRRRRRRRR0Fk__CM4<nR=4R''ERIC5MR5N#_8C_so25nR'=R4R'2NRM85N#_8C_so256R'=R4R'2NRM85N#_8C_so25cR'=Rj2'2R#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_Mn_4RR<=WI RERCM5_5#Ns8_Cno52RR='24'R8NMR_5#Ns8_C6o52RR='24'R8NMR#R5__N8s5Coc=2RR''j2C2RDR#C';j'
RRRRRRRR8CMRMoCC0sNC.Rzn
C;RRRRRRRRzV.nRH:RVNR58I8sHE80R(=RR8NMRlMk_DOCDc_nR4=RR8NMRlMk_DOCD._dRj=R2CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_Mn_4RR<='R4'IMECR#55__N8s5Con=2RR''42MRN8#R5__N8s5Co6=2RR''j2MRN8#R5__N8s5Coc=2RR''j2C2RDR#C';j'
RRRRRRRRRRRRRRRR0Is__CM4<nR= RWRCIEM5R5#8_N_osC5Rn2=4R''N2RM58R#8_N_osC5R62=jR''N2RM58R#8_N_osC5Rc2=jR''R22CCD#R''j;R
RRRRRRMRC8CRoMNCs0zCR.;nV
RRRRRRRRnz.oRR:H5VRNs88I0H8ERR=nMRN8kRMlC_ODnD_cRR=jMRN8kRMlC_ODdD_.RR=4o2RCsMCN
0CRRRRRRRRRRRRRRRRF_k0C4M_n=R<R''4RCIEM5R5#8_N_osC5R62=4R''N2RM58R#8_N_osC5Rc2=jR''R22CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C_R4n<W=R ERIC5MR5N#_8C_so256R'=R4R'2NRM85N#_8C_so25cR'=Rj2'2R#CDCjR''R;
RRRRRCRRMo8RCsMCNR0Czo.n;R
RRRRRR.Rzn:ERRRHV58N8s8IH0=ERRN6RMM8RkOl_C_DDd/.R=2R4RMoCC0sNCR
RRRRRRRRRRRRRRkRF0M_C_R4n<'=R4I'RERCM5_5#Ns8_CNo58I8sHE80-84RF0IMF2RcRM=RkOl_C_DDd2.2R#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_Mn_4RR<=WI RERCM5_5#Ns8_CNo58I8sHE80-84RF0IMF2RcRM=RkOl_C_DDd2.2R#CDCjR''R;
RRRRRCRRMo8RCsMCNR0CzE.n;R
RR-R-RRQV58N8s8IH0<ER=2R6RRMFI0sHCMRCNCLDRRFsFbk0kC0RMDNLCCR#D0CORoDFHMORCCC88R
RRRRRR.Rz(RR:H5VRNs88I0H8E=R<RRc2oCCMsCN0
RRRRRRRRRRRRRRRR0Fk__CM4<nR=4R''R;
RRRRRRRRRRRRRIRRsC0_Mn_4RR<=W
 ;RRRRRRRRCRM8oCCMsCN0R(z.;R
RR-R-RMtCC0sNCER0CqR)vCRODNDRM08Rs#H-0CN0
RSRRORzEU	_RH:RV#R5_8IH0NE_s$sN5Rd2>2RjRMoCC0sNCS
Sz	OE_6DCRH:RVIR5HE80RR>=U_*#I0H8Es_Ns5N$dN2RMI8RHE80RR>=Uo2RCsMCN
0CRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FzVR)4qvnRR:DCNLD#RHR1"1a&"RR0HMCsoC'NHloIC5HE802RR&"R7"&MRH0CCosl'HN5oCM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*cRR+M_klODCD_*d.dR.2&WR""RR&HCM0o'CsHolNCH5I8R0E-#RDLH_I820ER"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05lMk_DOCD._4U.*4URR+M_klODCD_*ncn+cRRlMk_DOCD._d*Rd.+nR4,CR8b20E2RR&"RX"&MRH0CCosl'HN5oCI0H8ERR-D_#LI0H8ERR+U
2;RRRRRRRRRRRRLHCoMS
SRRRRzv)q4:nRRqX)vX4nUS1
SRSRRFRbsl0RN5bR7>R=R8bN5H#_MC_soH5I8-0E4FR8IFM0R8IH0DE-#IL_HE802U,R,#RDLH_I8-0E4R2,q=jR>FRDI8_N8js52S,
SSSSSqRR4>R=RIDF_8N8s254,.RqRR=>D_FINs885,.2RRqd=D>RFNI_858sdR2,W= R>sRI0M_C_,4nRpWBi>R=RiBp,S
SSSSSRRRm=0>RlUb__54nj;22
SSSS#N#HRoM:FRVs[RHRRHMI0H8ER-48MFI0IFRHE80-LD#_8IH0oERCsMCN
0CSSSSRkRF0k_L#n_45lMk_DOCDn_4,2H[RR<=0_lbUn_455j2HI[-HE80+LD#_8IH0;E2
RRRRRRRRRRRRRRRR#RR_0Fk_osC52H[RR<=F_k0L_k#4Mn5kOl_C_DD4Hn,[I2RERCM50Fk__CM4=nRR''42DRC#'CRZ
';SSSSCRM8oCCMsCN0R#N#H;oM
RRRRRRRRRRRRUz.RV:RF[sRRRHM#H_I8_0ENNss$25d-84RF0IMFRR4oCCMsCN0
RRRRRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)Rzqnv4RD:RNDLCRRH#"a11"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloMC5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*nRM+RkOl_C_DDdd.*.&2RR""WRH&RMo0CCHs'lCNo58IH0-ERRLD#_8IH0-ERRU[*2RR&"R "&MRH0CCosl'HN5oCo_C0C_M880CbEk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*Rnc+kRMlC_ODdD_..*dR4+Rn8,RCEb02&2RR""XRH&RMo0CCHs'lCNo58IH0-ERRLD#_8IH0-ERR-5[4U2*2R;
RRRRRRRRRRRRRoLCHRM
RRRRRRRRRRRRRqz)vR4n:)RXqnv4XRU1
RRRRRRRRRRRRRRRRsbF0NRlb7R5RR=>#M_H_osC58IH0DE-#IL_HE80-[U*+8(RF0IMFHRI8-0ED_#LI0H8E*-U[R2,q=jR>FRDI8_N8js52q,R4>R=RIDF_8N8s254,.RqRR=>D_FINs885,.2
RRRRRRRRRRRRRRRRRRRRRRRRqRRd>R=RIDF_8N8s25d, RWRR=>I_s0C4M_nW,RBRpi=B>RpRi,m>R=Rb0l_4U_n25[2S;
SRSRR#RN#MHoRV:RFHsR[MRHR8(RF0IMFRRjoCCMsCN0
SSSSFRRkL0_k4#_nk5MlC_OD4D_nH,I8-0ED_#LI0H8E*-U[[+H2=R<Rb0l_4U_n25[52H[;R
RRRRRRRRRRRRRRRRR#k_F0C_soH5I8-0ED_#LI0H8E*-U[[+H2=R<R0Fk_#Lk_54nM_klODCD_,4nI0H8E#-DLH_I8-0EU+*[HR[2IMECRk5F0M_C_R4n=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR8CMRMoCC0sNC#RN#MHo;R
RRRRRRRRRRMRC8CRoMNCs0zCR.
U;SMSC8CRoMNCs0zCRO_E	D;C6
zSSO_E	oR06:VRHRH5I8R0E>U=RR8NMR8IH0lERFU8RRR>=6o2RCsMCN
0CRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FzVR)4qvnRR:DCNLD#RHR1"1a&"RR0HMCsoC'NHloIC5HE802RR&"R7"&MRH0CCosl'HN5oCM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*cRR+M_klODCD_*d.dR.2&WR""RR&HCM0o'CsHolNCH5I8R0E-#RDLH_I820ER"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05lMk_DOCD._4U.*4URR+M_klODCD_*ncn+cRRlMk_DOCD._d*Rd.+nR4,CR8b20E2RR&"RX"&MRH0CCosl'HN5oCI0H8ERR-D_#LI0H8ERR+U
2;RRRRRRRRRRRRLHCoMS
SRRRRzv)q4:nRRqX)vX4nUS1
SRSRRFRbsl0RN5bR7>R=R8bN5H#_MC_soH5I8-0E4FR8IFM0R8IH0DE-#IL_HE802U,R,#RDLH_I8-0E4R2,q=jR>FRDI8_N8js52S,
SSSSSqRR4>R=RIDF_8N8s254,.RqRR=>D_FINs885,.2RRqd=D>RFNI_858sdR2,W= R>sRI0M_C_,4nRpWBi>R=RiBp,S
SSSSSRRRm=0>RlUb__54n#H_I8_0ENNss$25d-242;S
SS#SN#MHoRV:RFHsR[MRHR8IH04E-RI8FMR0FI0H8E#-DLH_I8R0EoCCMsCN0
SSSSFRRkL0_k4#_nk5MlC_OD4D_n[,H2=R<Rb0l_4U_n_5#I0H8Es_Ns5N$d42-2[5H-8IH0DE+#IL_HE802R;
RRRRRRRRRRRRRRRRRF#_ks0_CHo5[<2R=kRF0k_L#n_45lMk_DOCDn_4,2H[RCIEMFR5kC0_Mn_4R'=R4R'2CCD#R''Z;S
SSMSC8CRoMNCs0NCR#o#HMR;
RRRRRRRRRzRR.:URRsVFRH[RM_R#I0H8Es_Ns5N$d.2-RI8FMR0FjCRoMNCs0RC
RRRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVzv)q4:nRRLDNCHDR#1R"1Ra"&MRH0CCosl'HN5oCI0H8E&2RR""7RH&RMo0CCHs'lCNo5lMk_DOCD._4U.*4URR+M_klODCD_*ncn+cRRlMk_DOCD._d*2d.R"&RW&"RR0HMCsoC'NHlo[C5*RU2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50EM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*cRR+M_klODCD_*d.d+.RR,4nRb8C02E2R"&RX&"RR0HMCsoC'NHlo5C5[2+4*;U2
RRRRRRRRRRRRLRRCMoH
RRRRRRRRRRRRzRR)4qvnRR:Xv)q4UnX1RR
RRRRRRRRRRRRRbRRFRs0lRNb5=7R>_R#HsM_CUo5*([+RI8FMR0FU2*[,jRqRR=>D_FINs885,j2RRq4=D>RFNI_858s4R2,q=.R>FRDI8_N8.s52R,
RRRRRRRRRRRRRRRRRRRRRRRRRRqd=D>RFNI_858sdR2,W= R>sRI0M_C_,4nRpWBi>R=RiBp,RRm=0>RlUb__54n[;22
SSSS#N#HRoM:FRVs[RHRRHM(FR8IFM0RojRCsMCN
0CSSSSRkRF0k_L#n_45lMk_DOCDn_4,[U*+2H[RR<=0_lbUn_455[2H;[2
RRRRRRRRRRRRRRRR#RR_0Fk_osC5[U*+2H[RR<=F_k0L_k#4Mn5kOl_C_DD4Un,*H[+[I2RERCM50Fk__CM4=nRR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRCRM8oCCMsCN0R#N#H;oM
RRRRRRRRRRRR8CMRMoCC0sNC.RzUS;
S8CMRMoCC0sNCORzEo	_0
6;SOSzEM	_RH:RVIR5HE80RU<R2CRoMNCs0RC
RRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)Rzqnv4RD:RNDLCRRH#"a11"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloMC5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*nRM+RkOl_C_DDdd.*.&2RR""WRH&RMo0CCHs'lCNo5Rj2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50EM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*cRR+M_klODCD_*d.d+.RR,4nRb8C02E2R"&RX&"RR0HMCsoC'NHloUC52R;
RRRRRRRRRLRRCMoH
RSSRzRR)4qvnRR:Xv)q4UnX1S
SSRRRRsbF0NRlb7R5RR=>b5N8#M_H_osC58IH04E-RI8FMR0FI0H8E#-DLH_I820E,,RURLD#_8IH04E-2q,Rj>R=RIDF_8N8s25j,S
SSSSSR4RqRR=>D_FINs885,42RRq.=D>RFNI_858s.R2,q=dR>FRDI8_N8ds52W,R >R=R0Is__CM4Rn,WiBpRR=>B,pi
SSSSRSSR=mR>lR0b__U4jn52
2;SSSSNH##o:MRRsVFRRH[HIMRHE80-84RF0IMFRRjoCCMsCN0
SSSSFRRkL0_k4#_nk5MlC_OD4D_n[,H2=R<Rb0l_4U_n25j52H[;R
RRRRRRRRRRRRRRRRR#k_F0C_so[5H2=R<R0Fk_#Lk_54nM_klODCD_,4nHR[2IMECRk5F0M_C_R4n=4R''C2RDR#C';Z'
SSSS8CMRMoCC0sNC#RN#MHo;S
SCRM8oCCMsCN0REzO	;_M
CSSMo8RCsMCNR0Cz	OE_
U;SOSzEc	_RH:RV#R5_8IH0NE_s$sN5R.2>2RjRMoCC0sNCR
RRRRRR.RzgR_c:VRHRH5I8R0E>c=R2CRoMNCs0RC
RRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)Rzqnv4RD:RNDLCRRH#"a11"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloMC5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*nRM+RkOl_C_DDdd.*.&2RR""WRH&RMo0CCHs'lCNo5Rj2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50EM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*cRR+M_klODCD_*d.d+.RR,4nRb8C02E2R"&RX&"RR0HMCsoC'NHlocC52R;
RRRRRRRRRLRRCMoH
RRRRRRRRRRRRqz)vR4n:qR)vX4nc
1RRRRRRRRRRRRRRRRRb0FsRblNRd57RR=>#M_H_osC5,d2RR7.=#>R__HMs5Co.R2,7=4R>_R#HsM_C4o527,Rj>R=RH#_MC_so25j,S
SSRRRRRRRRRRRRqRRj>R=RIDF_8N8s25j,4RqRR=>D_FINs885,42RRq.=D>RFNI_858s.
2,RRRRRRRRRRRRRRRRRRRRRRRRRdRqRR=>D_FINs885,d2RRW =I>RsC0_Mn_4,BRWp=iR>pRBi
,RSSSSSRSRm=dR>kRF0k_L#n_45lMk_DOCDn_4,,d2RRm.=F>RkL0_k4#_nk5MlC_OD4D_n2,.,S
SSSSSR4RmRR=>F_k0L_k#4Mn5kOl_C_DD44n,2m,Rj>R=R0Fk_#Lk_54nM_klODCD_,4nj;22
RRRRRRRRRRRRRRRRF#_ks0_Cdo52=R<R0Fk_#Lk_54nM_klODCD_,4ndI2RERCM50Fk__CM4=nRR''42DRC#'CRZ
';RRRRRRRRRRRRRRRR#k_F0C_so25.RR<=F_k0L_k#4Mn5kOl_C_DD4.n,2ERIC5MRF_k0C4M_nRR='24'R#CDCZR''R;
RRRRRRRRRRRRR#RR_0Fk_osC5R42<F=RkL0_k4#_nk5MlC_OD4D_n2,4RCIEMFR5kC0_Mn_4R'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRR_R#F_k0s5Coj<2R=kRF0k_L#n_45lMk_DOCDn_4,Rj2IMECRk5F0M_C_R4n=4R''C2RDR#C';Z'
RRRRRRRR8CMRMoCC0sNC.Rzg;_c
RRRRRRRRgz._:dRRRHV58IH0=ERRRd2oCCMsCN0
RRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVzv)q4:nRRLDNCHDR#1R"1Ra"&MRH0CCosl'HN5oCI0H8E&2RR""7RH&RMo0CCHs'lCNo5lMk_DOCD._4U.*4URR+M_klODCD_*ncn+cRRlMk_DOCD._d*2d.R"&RW&"RR0HMCsoC'NHlojC52RR&"R "&MRH0CCosl'HN5oCo_C0C_M880CbEk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*Rnc+kRMlC_ODdD_..*dR4+Rn8,RCEb02&2RR""XRH&RMo0CCHs'lCNo5;c2
RRRRRRRRRRRRoLCHRM
RRRRRRRRRzRR)4qvnRR:)4qvn1XcRR
RRRRRRRRRRRRRRFRbsl0RN5bR7=dR>jR''7,R.>R=RH#_MC_so25.,4R7RR=>#M_H_osC5,42RR7j=#>R__HMs5Coj
2,SRSSRRRRRRRRRRRRRRqj=D>RFNI_858sjR2,q=4R>FRDI8_N84s52q,R.>R=RIDF_8N8s25.,R
RRRRRRRRRRRRRRRRRRRRRRRRRq=dR>FRDI8_N8ds52W,R >R=R0Is__CM4Rn,WiBpRR=>B,piRS
SSSSSRdRmRR=>FMbC,.RmRR=>F_k0L_k#4Mn5kOl_C_DD4.n,2S,
SSSSSmRR4>R=R0Fk_#Lk_54nM_klODCD_,4n4R2,m=jR>kRF0k_L#n_45lMk_DOCDn_4,2j2;R
RRRRRRRRRRRRRR_R#F_k0s5Co.<2R=kRF0k_L#n_45lMk_DOCDn_4,R.2IMECRk5F0M_C_R4n=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRF#_ks0_C4o52=R<R0Fk_#Lk_54nM_klODCD_,4n4I2RERCM50Fk__CM4=nRR''42DRC#'CRZ
';RRRRRRRRRRRRRRRR#k_F0C_so25jRR<=F_k0L_k#4Mn5kOl_C_DD4jn,2ERIC5MRF_k0C4M_nRR='24'R#CDCZR''R;
RRRRRCRRMo8RCsMCNR0Cz_.gdS;
S8CMRMoCC0sNCORzEc	_;S
Sz	OE_:.RRRHV5I#_HE80_sNsN4$52RR>jo2RCsMCN
0CRRRRRRRRzRdj:FRVsRR[H5MR#H_I8_0ENNss$254R4-R2FR8IFM0RojRCsMCN
0CRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FzVR)4qvnRR:DCNLD#RHR1"1a&"RR0HMCsoC'NHloIC5HE802RR&"R7"&MRH0CCosl'HN5oCM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*cRR+M_klODCD_*d.dR.2&WR""RR&HCM0o'CsHolNCH5I8-0EU_*#I0H8Es_Ns5N$d.2-*.[-2RR&"R "&MRH0CCosl'HN5oCo_C0C_M880CbEk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*Rnc+kRMlC_ODdD_..*dR4+Rn8,RCEb02&2RR""XRH&RMo0CCHs'lCNo58IH0UE-*I#_HE80_sNsNd$52*-.[
2;RRRRRRRRRRRRLHCoMR
RRRRRRRRRR)Rzqnv4R):Rqnv4XR.1
RRRRRRRRRRRRRRRRsbF0NRlb7R5j>R=RH#_MC_soH5I8-0EU_*#I0H8Es_Ns5N$d.2-*.[-27,R4>R=RH#_MC_soH5I8-0EU_*#I0H8Es_Ns5N$d.2-*4[-2q,Rj>R=RIDF_8N8s25j,4RqRR=>D_FINs885,42RRq.=D>RFNI_858s.
2,RRRRRRRRRRRRRRRRRRRRRRRRRdRqRR=>D_FINs885,d2RRW =I>RsC0_Mn_4,BRWp=iR>pRBim,Rj>R=R0Fk_#Lk_54nM_klODCD_,4nI0H8E*-U#H_I8_0ENNss$25d-[.*-,.2
SSSSRSSRRm4=F>RkL0_k4#_nk5MlC_OD4D_nH,I8-0EU_*#I0H8Es_Ns5N$d.2-*4[-2
2;RRRRRRRRRRRRRRRR#k_F0C_soH5I8-0EU_*#I0H8Es_Ns5N$d.2-*4[-2=R<R0Fk_#Lk_54nM_klODCD_,4nI0H8E*-U#H_I8_0ENNss$25d-[.*-R42IMECRk5F0M_C_R4n=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRF#_ks0_CIo5HE80-#U*_8IH0NE_s$sN5-d2.-*[.<2R=kRF0k_L#n_45lMk_DOCDn_4,8IH0UE-*I#_HE80_sNsNd$52*-.[2-.RCIEMFR5kC0_Mn_4R'=R4R'2CCD#R''Z;R
RRRRRRMRC8CRoMNCs0zCRd
j;SMSC8CRoMNCs0zCRO_E	.S;
SEzO	R_4:VRHR_5#I0H8Es_Ns5N$j>2RRRj2oCCMsCN0
RRRRRRRR4zdRH:RVIR5HE80R8lFR=URRR42oCCMsCN0
RRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVzv)q4:nRRLDNCHDR#1R"1Ra"&MRH0CCosl'HN5oCI0H8E&2RR""7RH&RMo0CCHs'lCNo5lMk_DOCD._4U.*4URR+M_klODCD_*ncn+cRRlMk_DOCD._d*2d.R"&RW&"RR0HMCsoC'NHlojC52RR&"R "&MRH0CCosl'HN5oCo_C0C_M880CbEk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*Rnc+kRMlC_ODdD_..*dR4+Rn8,RCEb02&2RR""XRH&RMo0CCHs'lCNo5;42
RRRRRRRRRRRRoLCHRM
RRRRRRRRRzRR)4qvnRR:)4qvn1X4RR
RRRRRRRRRRRRRRFRbsl0RN5bR7>R=RH#_MC_so25j,jRqRR=>D_FINs885,j2RRq4=D>RFNI_858s4R2,q=.R>FRDI8_N8.s52R,
RRRRRRRRRRRRRRRRRRRRRRRRRRqd=D>RFNI_858sdR2,W= R>sRI0M_C_,4nRpWBi>R=RiBp,RRm=F>RkL0_k4#_nk5MlC_OD4D_n2,j2R;
RRRRRRRRRRRRR#RR_0Fk_osC5Rj2<F=RkL0_k4#_nk5MlC_OD4D_n2,jRCIEMFR5kC0_Mn_4R'=R4R'2CCD#R''Z;R
RRRRRRMRC8CRoMNCs0zCRd
4;SMSC8CRoMNCs0zCRO_E	4R;
RRRRCRM8oCCMsCN0R6z.;RRRRRRRR
RRRCRRMo8RCsMCNR0Cz;cc
8CMRONsECH0Os0kCFRM__sIOOEC	
;
---
--
--p-RNR#0HDlbCMlC0HN0FHMR#CR8VDNk0-
-
ONsECH0Os0kCCR#D0CO_lsNRRFV)_qv)HWR#F
OlMbFCRM0Xv)q4X.U4R1
b0FsRR5
RRRm:kRF00R#8F_Do;HO
RRRq:jRRRHM#_08DHFoOR;
R4RqRH:RM0R#8F_Do;HO
RRRq:.RRRHM#_08DHFoOR;
RdRqRH:RM0R#8F_Do;HO
RRRq:cRRRHM#_08DHFoOR;
R6RqRH:RM0R#8F_Do;HO
RRRq:nRRRHM#_08DHFoOR;
RRR7:MRHR8#0_oDFH
O;RWRRBRpi:MRHR8#0_oDFH
O;RWRR RR:H#MR0D8_FOoH
;R2
8CMRlOFbCFMM
0;
F
OlMbFCRM0Xv)qn.cX1b
RFRs05R
RRRmj:kRF00R#8F_Do;HO
RRRm:4RR0FkR8#0_oDFH
O;RqRRjRR:H#MR0D8_FOoH;R
RRRq4:MRHR8#0_oDFH
O;RqRR.RR:H#MR0D8_FOoH;R
RRRqd:MRHR8#0_oDFH
O;RqRRcRR:H#MR0D8_FOoH;R
RRRq6:MRHR8#0_oDFH
O;R7RRjRR:H#MR0D8_FOoH;R
RRR74:MRHR8#0_oDFH
O;RWRRBRpi:MRHR8#0_oDFH
O;RWRR RR:H#MR0D8_FOoH
;R2
8CMRlOFbCFMM
0;
lOFbCFMMX0R)dqv.1Xc
FRbs50R
RRRm:jRR0FkR8#0_oDFH
O;RmRR4RR:FRk0#_08DHFoOR;
R.RmRF:Rk#0R0D8_FOoH;R
RRRmd:kRF00R#8F_Do;HO
RRRq:jRRRHM#_08DHFoOR;
R4RqRH:RM0R#8F_Do;HO
RRRq:.RRRHM#_08DHFoOR;
RdRqRH:RM0R#8F_Do;HO
RRRq:cRRRHM#_08DHFoOR;
RjR7RH:RM0R#8F_Do;HO
RRR7:4RRRHM#_08DHFoOR;
R.R7RH:RM0R#8F_Do;HO
RRR7:dRRRHM#_08DHFoOR;
RBRWp:iRRRHM#_08DHFoOR;
R RWRH:RM0R#8F_Do
HOR
2;CRM8ObFlFMMC0O;
FFlbM0CMRqX)vXd.U
1
RsbF0
R5RmRRRF:Rk#0R0D8_FOoH_OPC05Fs(FR8IFM0R;j2
RRRq:jRRRHM#_08DHFoOR;
R4RqRH:RM0R#8F_Do;HO
RRRq:.RRRHM#_08DHFoOR;
RdRqRH:RM0R#8F_Do;HO
RRRq:cRRRHM#_08DHFoOR;
RRR7:MRHR8#0_oDFHPO_CFO0sR5(8MFI0jFR2R;
RBRWp:iRRRHM#_08DHFoOR;
R RWRH:RM0R#8F_Do
HOR
2;CRM8ObFlFMMC0
;
ObFlFMMC0)RXqnv4X
U1RsbF0
R5RmRRRF:Rk#0R0D8_FOoH_OPC05Fs(FR8IFM0R;j2
RRRq:jRRRHM#_08DHFoOR;
R4RqRH:RM0R#8F_Do;HO
RRRq:.RRRHM#_08DHFoOR;
RdRqRH:RM0R#8F_Do;HO
RRR7RR:H#MR0D8_FOoH_OPC05Fs(FR8IFM0R;j2
RRRWiBpRH:RM0R#8F_Do;HO
RRRW: RRRHM#_08DHFoO2
R;M
C8FROlMbFC;M0
$
0bDCRCFV0P_Cs0#RHRsNsN5$RjFR0RRd2FHVRMo0CC
s;0C$bRVDC0CFPs__0.#RHRsNsN5$RjFR0RR42FHVRMo0CC
s;VOkM0MHFR8bN5:HRR8#0_oDFHPO_CFO0sI;R4I,R.RR:HCM0o2CsR0sCkRsM#_08DHFoOC_POs0FR
H#PHNsNCLDRsPNR#:R0D8_FOoH_OPC05FsI44-RI8FMR0Fj
2;LHCoMR
RVRFs[MRHRsPN'MsNoDCRF
FbRRRRH5VR[=R<R2I.RC0EMSR
RNRPs25[RR:=H'5HD+FI[
2;S#CDCR
SRsPN5R[2:'=Rj
';S8CMR;HV
CRRMD8RF;Fb
sRRCs0kMNRPsC;
Mb8RN
8;VOkM0MHFR0oC_8IH0UE_58IH0RE:HCM0o2CsR0sCkRsMHCM0oRCsHP#
NNsHLRDCPRND:MRH0CCos=R:R
j;LHCoMR
RPRND:I=RHE80/
U;RVRHRI55HE80R8lFRRU2>2RcRC0EMR
RRNRPD=R:RDPNR4+R;R
RCRM8H
V;RCRs0MksRDPN;M
C8CRo0H_I8_0EUV;
k0MOHRFMo_C0I0H8E5_.I0H8EH:RMo0CCRs2skC0sHMRMo0CCHsR#N
PsLHNDPCRN:DRR0HMCsoCRR:=jL;
CMoH
PRRN:DR=HRI8/0E.R;
R0sCkRsMP;ND
8CMR0oC_8IH0.E_;k
VMHO0FoMRCI0_HE8058IH0:ERR0HMCsoC2CRs0MksRVDC0CFPs__0.#RH
sPNHDNLCNRPDRR:D0CVFsPC_.0_;C
Lo
HMRNRPD254RR:=o_C0I0H8E5_.I0H8E
2;RVRHRH5I8R0ElRF8.RR=j02RE
CMRRRRP5NDj:2R=;Rj
CRRD
#CRRRRP5NDj:2R=;R4
CRRMH8RVR;
R0sCkRsMP;ND
8CMR0oC_8IH0
E;VOkM0MHFR0oC_8IH0IE5HE80RH:RMo0CCRs2skC0sDMRCFV0P_Cs0#RH
sPNHDNLCNRPDRR:D0CVFsPC_:0R=jR5,,RjRRj,j
2;LHCoMR
RP5NDd:2R=CRo0H_I8_0EUH5I820E;R
ROCN#RH5I8R0ElRF8UH2R#R
RIMECR|cRR=dR>NRPD25.RR:=4R;
RCIEMRR.=P>RN4D52=R:R
4;RERIC4MRRR=>P5NDj:2R=;R4
IRRERCMFC0Es=#R>kRMD
D;RMRC8NRO#
C;RCRs0MksRDPN;M
C8CRo0H_I8;0E
MOF#M0N0HRI8_0ENNss$RR:D0CVFsPC_:0R=CRo0H_I850EI0H8E
2;O#FM00NMR8IH0NE_s$sN_Rnc:CRDVP0FC0s__:.R=CRo0H_I850EI0H8E
2;VOkM0MHFR0oC_lMk_U4.5b8C0RE:HCM0o2CsR0sCkRsMHCM0oRCsHP#
NNsHLRDCPRND:MRH0CCos=R:R
j;LHCoMR
RPRND:8=RCEb0/U4.;R
RH5VR5b8C0lERF48R.RU2>4R4.02RE
CMRRRRPRND:P=RN+DRR
4;RMRC8VRH;R
RskC0sPMRN
D;CRM8o_C0M_kl4;.U
MVkOF0HMCRo0C_DVP0FCns_cC58bR0E:MRH0CCoss2RCs0kMMRH0CCos#RH
oLCHRM
R0sCk5sM80CbEFRl8.R4U
2;CRM8o_C0D0CVFsPC_;nc
MVkOF0HMCRo0k_Mlc_n5b8C0:ERR0HMCsoC2CRs0MksR0HMCsoCR
H#PHNsNCLDRDPNRH:RMo0CC:sR=;Rj
oLCHRM
RRHV5b8C0<ER=4R4.MRN8CR8bR0E>URc2ER0CRM
RRRRPRND:4=R;R
RCRM8H
V;RCRs0MksRDPN;M
C8CRo0k_Mlc_n;k
VMHO0FoMRCD0_CFV0P5Cs80CbERR:HCM0o;CsRGlNRH:RMo0CCRs2skC0sHMRMo0CCHsR#N
PsLHNDPCRN:DRR0HMCsoCRR:=jL;
CMoH
HRRV8R5CEb0Rl-RN>GR=2RjRC0EMR
RRNRPD=R:Rb8C0-ERRGlN;R
RCCD#
RRRRDPNRR:=80CbER;
R8CMR;HV
sRRCs0kMN5PD
2;CRM8o_C0D0CVFsPC;k
VMHO0FoMRCM0_kdl_.C58bR0E:MRH0CCoss2RCs0kMMRH0CCos#RH
sPNHDNLCNRPDRR:HCM0oRCs:j=R;C
Lo
HMRVRHRC58bR0E<c=RUMRN8CR8bR0E>nR42ER0CRM
RRRRPRND:4=R;R
RCRM8H
V;RCRs0MksRDPN;M
C8CRo0k_Ml._d;k
VMHO0FoMRCM0_k4l_nC58bR0E:MRH0CCoss2RCs0kMMRH0CCos#RH
sPNHDNLCNRPDRR:HCM0oRCs:j=R;C
Lo
HMRVRHRC58bR0E<4=RnMRN8CR8bR0E>2RjRC0EMR
RRPRRN:DR=;R4
CRRMH8RVR;
R0sCkRsMP;ND
8CMR0oC_lMk_;4n
MVkOF0HMCRo0M_C8C_8b50E#CHxRH:RMo0CC;sRRb8C0:ERR0HMCsoC2CRs0MksR0HMCsoCR
H#PHNsNCLDRMlH_x#HCRR:HCM0oRCs:j=R;C
Lo
HMRHRlMH_#x:CR=CR8b;0E
HRRV#R5HRxC<CR8b20ERC0EMR
RRHRlMH_#x:CR=HR#x
C;RMRC8VRH;R
RskC0slMRH#M_H;xC
8CMR0oC_8CM_b8C0
E;-F-OMN#0MM0RkOl_C#DDRH:RMo0CC:sR=5R55b8C0-ERRR42/.Rd2RR+5855CEb0R4-R2FRl8.Rd2RR/42n2;RRR-y-RRRFV)dqv.1X4RDOCDM#RCCC88OR
F0M#NRM0M_klODCD_U4.RH:RMo0CC:sR=CRo0k_Ml._4UC58b20E;F
OMN#0MD0RCFV0P_Csn:cRR0HMCsoCRR:=o_C0D0CVFsPC_5nc80CbE
2;O#FM00NMRlMk_DOCDc_nRH:RMo0CC:sR=CRo0k_Mlc_n5VDC0CFPsc_n2O;
F0M#NRM0D0CVFsPC_Rd.:MRH0CCos=R:R0oC_VDC0CFPsC5DVP0FCns_cn,Rc
2;O#FM00NMRlMk_DOCD._dRH:RMo0CC:sR=CRo0k_Ml._d5VDC0CFPs._d2O;
F0M#NRM0D0CVFsPC_R4n:MRH0CCos=R:R0oC_VDC0CFPsC5DVP0FCds_.d,R.
2;O#FM00NMRlMk_DOCDn_4RH:RMo0CC:sR=CRo0k_Mln_45VDC0CFPsn_42
;
0C$bR0Fk_#Lk_b0$C._4U#RHRsNsN5$RM_klODCD_U4.RI8FMR0FjI,RHE80-84RF0IMF2RjRRFV#_08DHFoO0;
$RbCF_k0L_k#0C$b_RncHN#Rs$sNRk5MlC_ODnD_cFR8IFM0RRj,I0H8ER-48MFI0jFR2VRFR8#0_oDFH
O;0C$bR0Fk_#Lk_b0$C._dRRH#NNss$MR5kOl_C_DDd8.RF0IMF,RjR8IH04E-RI8FMR0FjF2RV0R#8F_Do;HO
b0$CkRF0k_L#$_0b4C_n#RHRsNsN5$RM_klODCD_R4n8MFI0jFR,HRI8-0E4FR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNR0Fk_#Lk_U4.RF:RkL0_k0#_$_bC4;.URRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$F8VRFRk05bHMk00RFsR0H0-#N#0C2H
#oDMNR0Fk_#Lk_Rnc:kRF0k_L#$_0bnC_cR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFRk8F0HR5M0bkRR0F0-sH#00NC
#2#MHoNFDRkL0_kd#_.RR:F_k0L_k#0C$b_;d.RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$F8VRFRk05bHMk00RFsR0H0-#N#0C2H
#oDMNR0Fk_#Lk_R4n:kRF0k_L#$_0b4C_nR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFRk8F0HR5M0bkRR0F0-sH#00NC
#2#MHoNFDRkC0_MRR:#_08DHFoOC_POs0F5lMk_DOCD._4UFR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--CLMNDRC#VRFs0-sH#00NC##
HNoMDkRF0M_C_Rnc:0R#8F_Do;HO
o#HMRNDF_k0CdM_.RR:#_08DHFoO#;
HNoMDkRF0M_C_R4n:0R#8F_Do;HO
o#HMRNDI_s0C:MRR8#0_oDFHPO_CFO0sk5MlC_OD4D_.8URF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RHIs0CCRMDNLCV#RFCsRNROEsRFIF)VRqOvRC#DD
o#HMRNDI_s0CnM_cRR:#_08DHFoO#;
HNoMDsRI0M_C_Rd.:0R#8F_Do;HO
o#HMRNDI_s0C4M_nRR:#_08DHFoO#;
HNoMDMRH_osCR#:R0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--k8#CRR0FsHCo#s0CRh7QRH
#oDMNR0Fk_osCR#:R0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-k-R#RC80sFRC#oH0RCs7amz
o#HMRNDNs8_C:oRR8#0_oDFHPO_CFO0s85N8HsI8-0E4FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-#RkC08RFCRso0H#CqsR7
7)#MHoNDDRFNI_8R8s:0R#8F_Do_HOP0COFns5RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-R8N8sHRL0H#RM0bkRR0F)RqvODCD#cR5R0LH#CRsJskHC
82O#FM00NMRLD#_8IH0:ERR0HMCsoCRR:=I0H8E*-U58IH0NE_s$sN5-d24c2-*8IH0NE_s$sN5-.2.H*I8_0ENNss$254-8IH0NE_s$sN5;j2
b0$ClR0bs_NsUN$RRH#NNss$IR5HE80_sNsNd$52R-48MFI0jFR2VRFR8#0_oDFHPO_CFO0sR5(8MFI0jFR2#;
HNoMDlR0b__UdR.,0_lbUn_4R0:RlNb_s$sNUN;
0H0sLCk0Rs\3NFl_VCV#0:\RRs#0H;Mo
oLCH
M
RRRR-Q-RV8RN8HsI8R0E<RR(NH##o'MRj0'RFMRkk8#CR0LH#R
RRjRzRRR:H5VRNs88I0H8ERR=4o2RCsMCN
0CRRRRRRRRD_FINs88RR<="jjjj"jjRN&R8C_so25j;R
RRMRC8CRoMNCs0zCRjR;
RzRR4:RRRRHV58N8s8IH0=ERRR.2oCCMsCN0
RRRRRRRRIDF_8N8s=R<Rj"jj"jjRN&R8C_soR548MFI0jFR2R;
RCRRMo8RCsMCNR0Cz
4;RRRRzR.R:VRHR85N8HsI8R0E=2RdRMoCC0sNCR
RRRRRRFRDI8_N8<sR=jR"j"jjRN&R8C_soR5.8MFI0jFR2R;
RCRRMo8RCsMCNR0Cz
.;RRRRzRdR:VRHR85N8HsI8R0E=2RcRMoCC0sNCR
RRRRRRFRDI8_N8<sR=jR"jRj"&8RN_osC58dRF0IMF2Rj;R
RRMRC8CRoMNCs0zCRdS;
z:cSRRHV58N8s8IH0=ERRR62oCCMsCN0
DSSFNI_8R8s<"=RjRj"&8RN_osC58cRF0IMF2Rj;C
SMo8RCsMCNR0Cz
c;SSz6:VRHR85N8HsI8R0E=2RnRMoCC0sNCS
SD_FINs88RR<='Rj'&8RN_osC586RF0IMF2Rj;R
RRMRC8CRoMNCs0zCR6R;
RzRRn:RRRRHV58N8s8IH0>ERRRn2oCCMsCN0
RRRRRRRRIDF_8N8s=R<R_N8s5ConFR8IFM0R;j2
RRRR8CMRMoCC0sNCnRz;R

R-RR-VRQRH58MC_sos2RC#oH0RCs7RQhkM#HopRBiR
RR(RzRRR:H5VR8_HMs2CoRMoCC0sNCR
RRRRRRsRbF#OC#BR5pRi,72QhRoLCHRM
RRRRRRRRRHRRVBR5p=iRR''4R8NMRiBp'CCPMR020MEC
RRRRRRRRRRRRRRRR_HMsRCo<7=RQ
h;RRRRRRRRRRRRCRM8H
V;RRRRRRRRCRM8bOsFC;##
RRRR8CMRMoCC0sNC(Rz;R
RRURzRRR:H5VRMRF08_HMs2CoRMoCC0sNCR
RRRRRRRRRRMRH_osCRR<=7;Qh
RRRR8CMRMoCC0sNCURz;R

R-RR-VRQRF58ks0_CRo2sHCo#s0CRz7ma#RkHRMomiBp
RRRRRzgRH:RV8R5F_k0s2CoRMoCC0sNCR
RRRRRRsRbF#OC#mR5B,piR0Fk_osC2CRLo
HMRRRRRRRRRRRRH5VRmiBpR'=R4N'RMm8RB'piCMPC002RE
CMRRRRRRRRRRRRRRRR7amzRR<=F_k0s;Co
RRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMRFbsO#C#;R
RRMRC8CRoMNCs0zCRgR;
RzRR4RjR:VRHRF5M0FR8ks0_CRo2oCCMsCN0
RRRRRRRRRRRRz7ma=R<R0Fk_osC;R
RRMRC8CRoMNCs0zCR4
j;
RRRRR--Q5VRNs88_osC2CRso0H#CqsR7R7)kM#HopRBiR
RR4Rz4:RRRRHV58N8sC_soo2RCsMCN
0CRRRRRRRRbOsFCR##5iBp,7Rq7R)2LHCoMR
RRRRRRRRRRVRHRp5BiRR='R4'NRM8B'piCMPC002RE
CMRRRRRRRRRRRRRRRRNs8_C<oR=7Rq7N)58I8sHE80-84RF0IMF2Rj;R
RRRRRRRRRRMRC8VRH;R
RRRRRRMRC8sRbF#OC#R;
RCRRMo8RCsMCNR0Cz;44
RRRR.z4RH:RVMR5FN0R8_8ss2CoRMoCC0sNCR
RRRRRRRRRR8RN_osCRR<=q)77;R
RRMRC8CRoMNCs0zCR4
.;RRRRRRRR
RRRRR--tCCMsCN0RC0ERv)qRDOCDN#RM#8RCODC0FRDo
HORRRRzR4d:FRVsRRHH5MRM_klODCD_U4.R4-R2FR8IFM0RojRCsMCN
0CRRRR-Q-RVNR58I8sHE80R6>R2CRMC08RFsROCCN0RHIs0CCRMDNLCMRN8kRF00bkRNCMLRDC#CCDOD0RFOoH
RRRRRRRRcz4RH:RVNR58I8sHE80R(>R2CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_M25HRR<='R4'IMECR85N_osC58N8s8IH04E-RI8FMR0F(=2RRRH2CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R ERIC5MRNs8_CNo58I8sHE80-84RF0IMF2R(RH=R2DRC#'CRj
';RRRRRRRRCRM8oCCMsCN0Rcz4;R
RR-R-RRQV58N8s8IH0<ER=2R6RRMFI0sHCMRCNCLDRRFsFbk0kC0RMDNLCCR#D0CORoDFHMORCCC88R
RRRRRR4Rz6RR:H5VRNs88I0H8E=R<RR(2oCCMsCN0
RRRRRRRRRRRRRRRR0Fk_5CMH<2R=4R''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=W
 ;RRRRRRRRCRM8oCCMsCN0R6z4;R
RR-R-RMtCC0sNCER0CqR)vCRODRD#NRM80-sH#00NCR#
RRRRRzRR4:nRRsVFRH[RMIR5HE80R4-R2FR8IFM0RojRCsMCN
0CRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FzVR)4qv.:URRLDNCHDR#1R"1Ra"&MRH0CCosl'HN5oCI0H8E&2RR""7RH&RMo0CCHs'lCNo54H*.RU2&WR""RR&HCM0o'CsHolNC25[R"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05+5H442*.RU,80CbER22&XR""RR&HCM0o'CsHolNC+5[4
2;RRRRRRRRRRRRLHCoMR
RRRRRRRRRR)Rzq.v4URR:Xv)q4X.U4
1RRRRRRRRRRRRRRRRRb0FsRblNRR57=H>RMC_so25[,jRqRR=>D_FINs885,j2RRq4=D>RFNI_858s4R2,q=.R>FRDI8_N8.s52R,
RRRRRRRRRRRRRRRRRRRRRRRRRRqd=D>RFNI_858sdR2,q=cR>FRDI8_N8cs52q,R6>R=RIDF_8N8s256,nRqRR=>D_FINs885,n2
SSSSRSSRRW =I>RsC0_M25H,BRWp=iR>pRBim,RRR=>F_k0L_k#45.UH2,[2R;
RRRRRRRRRRRRRFRRks0_C[o52=R<R0Fk_#Lk_U4.5[H,2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRCRRMo8RCsMCNR0Cz;4n
RRRRMRC8CRoMNCs0zCR4Rd;RRRRRRRRR
RRRRRRRRR
R-RR-CRtMNCs0NCRRR4nI8FsRC8CbqR)vCRODHDRVbRNbbsFs0HNCRRRRRRRRRRRRRRR
RRRR(z4RH:RVMR5kOl_C_DDn=cRRR42oCCMsCN0
RRRRR--Q5VRNs88I0H8ERR>(M2RCRC80OFRs0CNCsRIHR0CCLMNDNCRMF8Rkk0b0MRCNCLDRD#CCRO0DHFoOR
RRRRRR4RzU:NRRRHV58N8s8IH0>ERRR(2oCCMsCN0
RRRRRRRRRRRRRRRR0Fk__CMn<cR=4R''ERIC5MR5_N8s5CoNs88I0H8ER-48MFI0(FR2RR=M_klODCD_U4.2MRN8NR58C_so25nR'=Rj2'2R#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_Mc_nRR<=WI RERCM585N_osC58N8s8IH04E-RI8FMR0F(=2RRlMk_DOCD._4UN2RM58RNs8_Cno52RR='2j'2DRC#'CRj
';RRRRRRRRCRM8oCCMsCN0RUz4NR;
RRRRRzRR4RUL:VRHR85N8HsI8R0E=RR(NRM8M_klODCD_U4.Rj=R2CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_Mc_nRR<='R4'IMECRN558C_so25nR'=Rj2'2R#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_Mc_nRR<=WI RERCM585N_osC5Rn2=jR''R22CCD#R''j;R
RRRRRRMRC8CRoMNCs0zCR4;UL
RRRRR--Q5VRNs88I0H8E=R<RR62MIFRsCH0RNCMLRDCFFsRkk0b0MRCNCLDRD#CCRO0DHFoOCRMC88C
RRRRRRRRgz4RH:RVNR58I8sHE80RR<=no2RCsMCN
0CRRRRRRRRRRRRRRRRF_k0CnM_c=R<R''4;R
RRRRRRRRRRRRRRsRI0M_C_Rnc<W=R R;
RRRRRCRRMo8RCsMCNR0Cz;4g
RRRRR--tCCMsCN0RC0ERv)qRDOCDMRN8sR0H0-#N
0CSRRRREzO	R_.:VRHRH5I8_0ENNss$c_n5R42>2RjRMoCC0sNCR
RRRRRR.RzjRR:VRFs[MRHRH5I8_0ENNss$c_n5R42-2R4RI8FMR0FjCRoMNCs0RC
RRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)RzqcvnRD:RNDLCRRH#"a11"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloMC5kOl_C_DD4*.U42.UR"&RW&"RR0HMCsoC'NHloIC5HE80R.-R*-[RRR.2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50EM_klODCD_U4.*U4.Rn+Rc8,RCEb02&2RR""XRH&RMo0CCHs'lCNo58IH0-ERR[.*2R;
RRRRRRRRRLRRCMoH
RRRRRRRRRRRRqz)vRnc:)RXqcvnXR.1
RRRRRRRRRRRRRRRRsbF0NRlb7R54>R=R_HMs5CoI0H8E*-.[2-4,jR7RR=>HsM_CIo5HE80-[.*-,.2RRqj=D>RFNI_858sjR2,q=4R>FRDI8_N84s52q,R.>R=RIDF_8N8s25.,R
RRRRRRRRRRRRRRRRRRRRRRRRRq=dR>FRDI8_N8ds52q,Rc>R=RIDF_8N8s25c,6RqRR=>D_FINs885,62
SSSSRSSRRW =I>RsC0_Mc_n,BRWp=iR>pRBim,R4>R=R0Fk_#Lk_5ncM_klODCD_,ncI0H8E*-.[2-4,jRmRR=>F_k0L_k#nMc5kOl_C_DDnIc,HE80-[.*-2.2;R
RRRRRRRRRRRRRRkRF0C_soH5I8-0E.-*[4<2R=kRF0k_L#c_n5lMk_DOCDc_n,8IH0.E-*4[-2ERIC5MRF_k0CnM_cRR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_CIo5HE80-[.*-R.2<F=RkL0_kn#_ck5MlC_ODnD_cH,I8-0E.-*[.I2RERCM50Fk__CMn=cRR''42DRC#'CRZ
';RRRRRRRRR8CMRMoCC0sNC.RzjS;
SMRC8CRoMNCs0zCRO_E	.S;
SORzE4	_RH:RVIR5HE80_sNsNn$_c25jRj>R2CRoMNCs0RC
RRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)RzqcvnRD:RNDLCRRH#"a11"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloMC5kOl_C_DD4*.U42.UR"&RW&"RR0HMCsoC'NHloIC5HE80R.-R*8IH0NE_s$sN_5nc4-2RRR42& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50EM_klODCD_U4.*U4.Rn+Rc8,RCEb02&2RR""XRH&RMo0CCHs'lCNo58IH0-ERRI.*HE80_sNsNn$_c2542R;
RRRRRRRRRLRRCMoH
RRRRRRRRRRRRqz)vRnc:qR)vXnc4
1RRRRRRRRRRRRRRRRRb0FsRblNRR57=H>RMC_soH5I8-0E.H*I8_0ENNss$c_n5-424R2,q=jR>FRDI8_N8js52q,R4>R=RIDF_8N8s254,.RqRR=>D_FINs885,.2
RRRRRRRRRRRRRRRRRRRRRRRRqRRd>R=RIDF_8N8s25d,cRqRR=>D_FINs885,c2RRq6=D>RFNI_858s6
2,SSSSSRSRW= R>sRI0M_C_,ncRpWBi>R=RiBp,RRm=F>RkL0_kn#_ck5MlC_ODnD_cH,I8-0E.H*I8_0ENNss$c_n5-424;22
RRRRRRRRRRRRRRRR0Fk_osC58IH0.E-*8IH0NE_s$sN_5nc442-2=R<R0Fk_#Lk_5ncM_klODCD_,ncI0H8E*-.I0H8Es_Ns_N$n4c522-4RCIEMFR5kC0_Mc_nR'=R4R'2CCD#R''Z;R
RRRRRRCRRMo8RCsMCNR0Cz	OE_
4;RRRRRCSRMo8RCsMCNR0Cz;4(RRRRRRRRR
R
RRRR-t-RCsMCNR0CNnR4RsIF8CR8C)bRqOvRCRDDHNVRbFbsbNsH0RCRRRRRRRRRRRRRRR
RR.Rz4RR:H5VRM_klODCD_Rd.=2R4RMoCC0sNCR
RR-R-RRQV58N8s8IH0>ERRR62M8CCRR0FONsC0ICRsCH0RNCMLRDCNRM8Fbk0kC0RMDNLCCR#D0CORoDFHRO
RRRRRzRR.R.N:VRHR85N8HsI8R0E>RR(NRM8M_klODCD_Rnc=2R4RMoCC0sNCR
RRRRRRRRRRRRRRkRF0M_C_Rd.<'=R4I'RERCM585N_osC58N8s8IH04E-RI8FMR0F(=2RRlMk_DOCD._4UN2RM58RNs8_Cno52RR='24'R8NMR85N_osC5R62=jR''R22CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C_Rd.<W=R ERIC5MR5_N8s5CoNs88I0H8ER-48MFI0(FR2RR=M_klODCD_U4.2MRN8NR58C_so25nR'=R4R'2NRM85_N8s5Co6=2RR''j2C2RDR#C';j'
RRRRRRRR8CMRMoCC0sNC.Rz.
N;RRRRRRRRzL..RH:RVNR58I8sHE80R(>RR8NMRlMk_DOCDc_nRR/=4o2RCsMCN
0CRRRRRRRRRRRRRRRRF_k0CdM_.=R<R''4RCIEM5R5Ns8_CNo58I8sHE80-84RF0IMF2R(RM=RkOl_C_DD42.UR8NMR85N_osC5Rn2=jR''N2RM58RNs8_C6o52RR='2j'2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0CdM_.=R<RRW IMECRN558C_so85N8HsI8-0E4FR8IFM0RR(2=kRMlC_OD4D_.RU2NRM85_N8s5Con=2RR''j2MRN8NR58C_so256R'=Rj2'2R#CDCjR''R;
RRRRRCRRMo8RCsMCNR0CzL..;R
RRRRRR.Rz.:ORRRHV58N8s8IH0=ERRN(RMM8RkOl_C_DDn=cRRR42oCCMsCN0
RRRRRRRRRRRRRRRR0Fk__CMd<.R=4R''ERIC5MR5_N8s5Con=2RR''42MRN8NR58C_so256R'=Rj2'2R#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_M._dRR<=WI RERCM585N_osC5Rn2=4R''N2RM58RNs8_C6o52RR='2j'2DRC#'CRj
';RRRRRRRRCRM8oCCMsCN0R.z.OR;
RRRRRzRR.R.8:VRHR85N8HsI8R0E=RRnNRM8M_klODCD_Rnc/4=R2CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_M._dRR<='R4'IMECRN558C_so85N8HsI8-0E4FR8IFM0RR62=kRMlC_ODnD_cR22CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C_Rd.<W=R ERIC5MR5_N8s5CoNs88I0H8ER-48MFI06FR2RR=M_klODCD_2nc2DRC#'CRj
';RRRRRRRRCRM8oCCMsCN0R.z.8R;
R-RR-VRQR85N8HsI8R0E<6=R2FRMRHIs0CCRMDNLCsRFR0FkbRk0CLMND#CRCODC0FRDoRHOM8CCCR8
RRRRRzRR.:dRRRHV58N8s8IH0<ER=2R6RMoCC0sNCR
RRRRRRRRRRRRRRkRF0M_C_Rd.<'=R4
';RRRRRRRRRRRRRRRRI_s0CdM_.=R<R;W 
RRRRRRRR8CMRMoCC0sNC.RzdR;
R-RR-CRtMNCs00CRE)CRqOvRCRDDNRM80-sH#00NCR
SRzRRO_E	URR:H5VRI0H8Es_Ns5N$d>2RRRj2oCCMsCN0
zSSO_E	DRC6:VRHRH5I8R0E>U=R*8IH0NE_s$sN5Rd2NRM8I0H8E=R>RRU2oCCMsCN0
RRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVzv)qd:.RRLDNCHDR#1R"1Ra"&MRH0CCosl'HN5oCI0H8E&2RR""7RH&RMo0CCHs'lCNo5lMk_DOCD._4U.*4URR+M_klODCD_*ncnRc2&WR""RR&HCM0o'CsHolNCH5I8R0E-#RDLH_I820ER"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05lMk_DOCD._4U.*4URR+M_klODCD_*ncn+cRR,d.Rb8C02E2R"&RX&"RR0HMCsoC'NHloIC5HE80RD-R#IL_HE80RU+R2R;
RRRRRRRRRLRRCMoH
RSSRzRR)dqv.RR:Xv)qdU.X1S
SSRRRRsbF0NRlb7R5RR=>b5N8HsM_CIo5HE80-84RF0IMFHRI8-0ED_#LI0H8ER2,UD,R#IL_HE80-,42RRqj=D>RFNI_858sj
2,SSSSSRSRq=4R>FRDI8_N84s52q,R.>R=RIDF_8N8s25.,dRqRR=>D_FINs885,d2RRqc=D>RFNI_858scR2,W= R>sRI0M_C_,d.RpWBi>R=RiBp,S
SSSSSRRRm=0>RlUb__5d.j;22
SSSS#N#HRoM:FRVs[RHRRHMI0H8ER-48MFI0IFRHE80-LD#_8IH0oERCsMCN
0CSSSSRkRF0k_L#._d5lMk_DOCD._d,2H[RR<=0_lbU._d55j2HI[-HE80+LD#_8IH0;E2
RRRRRRRRRRRRRRRRFRRks0_CHo5[<2R=kRF0k_L#._d5lMk_DOCD._d,2H[RCIEMFR5kC0_M._dR'=R4R'2CCD#R''Z;S
SSMSC8CRoMNCs0NCR#o#HMR;
RRRRRRRRRzRR.:URRsVFRH[RMHRI8_0ENNss$25d-84RF0IMFRR4oCCMsCN0
RRRRRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)Rzq.vdRD:RNDLCRRH#"a11"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloMC5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*n2RR&"RW"&MRH0CCosl'HN5oCI0H8ERR-D_#LI0H8ERR-[2*UR"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05lMk_DOCD._4U.*4URR+M_klODCD_*ncn+cRR,d.Rb8C02E2R"&RX&"RR0HMCsoC'NHloIC5HE80RD-R#IL_HE80R5-R[2-4*;U2
RRRRRRRRRRRRLRRCMoH
RRRRRRRRRRRRzRR)dqv.RR:Xv)qdU.X1RR
RRRRRRRRRRRRRbRRFRs0lRNb5=7R>MRH_osC58IH0DE-#IL_HE80-[U*+8(RF0IMFHRI8-0ED_#LI0H8E*-U[R2,q=jR>FRDI8_N8js52q,R4>R=RIDF_8N8s254,.RqRR=>D_FINs885,.2
RRRRRRRRRRRRRRRRRRRRRRRRqRRd>R=RIDF_8N8s25d,cRqRR=>D_FINs885,c2RRW =I>RsC0_M._d,BRWp=iR>pRBim,RRR=>0_lbU._d52[2;S
SSRRRR#N#HRoM:FRVs[RHRRHM(FR8IFM0RojRCsMCN
0CSSSSRkRF0k_L#._d5lMk_DOCD._d,8IH0DE-#IL_HE80-[U*+2H[RR<=0_lbU._d55[2H;[2
RRRRRRRRRRRRRRRRFRRks0_CIo5HE80-LD#_8IH0UE-*H[+[<2R=kRF0k_L#._d5lMk_DOCD._d,8IH0DE-#IL_HE80-[U*+2H[RCIEMFR5kC0_M._dR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRMRC8CRoMNCs0NCR#o#HMR;
RRRRRRRRRCRRMo8RCsMCNR0Cz;.U
CSSMo8RCsMCNR0Cz	OE_6DC;S
Sz	OE_6o0RH:RVIR5HE80RR>=UMRN8HRI8R0ElRF8U=R>RR62oCCMsCN0
RRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVzv)qd:.RRLDNCHDR#1R"1Ra"&MRH0CCosl'HN5oCI0H8E&2RR""7RH&RMo0CCHs'lCNo5lMk_DOCD._4U.*4URR+M_klODCD_*ncnRc2&WR""RR&HCM0o'CsHolNCH5I8R0E-#RDLH_I820ER"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05lMk_DOCD._4U.*4URR+M_klODCD_*ncn+cRR,d.Rb8C02E2R"&RX&"RR0HMCsoC'NHloIC5HE80RD-R#IL_HE80RU+R2R;
RRRRRRRRRLRRCMoH
RSSRzRR)dqv.RR:Xv)qdU.X1S
SSRRRRsbF0NRlb7R5RR=>b5N8HsM_CIo5HE80-84RF0IMFHRI8-0ED_#LI0H8ER2,UD,R#IL_HE80-,42RRqj=D>RFNI_858sj
2,SSSSSRSRq=4R>FRDI8_N84s52q,R.>R=RIDF_8N8s25.,dRqRR=>D_FINs885,d2RRqc=D>RFNI_858scR2,W= R>sRI0M_C_,d.RpWBi>R=RiBp,S
SSSSSRRRm=0>RlUb__5d.I0H8Es_Ns5N$d42-2
2;SSSSNH##o:MRRsVFRRH[HIMRHE80-84RF0IMFHRI8-0ED_#LI0H8ECRoMNCs0SC
SRSSR0Fk_#Lk_5d.M_klODCD_,d.HR[2<0=RlUb__5d.I0H8Es_Ns5N$d42-2[5H-8IH0DE+#IL_HE802R;
RRRRRRRRRRRRRRRRR0Fk_osC52H[RR<=F_k0L_k#dM.5kOl_C_DDdH.,[I2RERCM50Fk__CMd=.RR''42DRC#'CRZ
';SSSSCRM8oCCMsCN0R#N#H;oM
RRRRRRRRRRRRUz.RV:RF[sRRRHMI0H8Es_Ns5N$d.2-RI8FMR0FjCRoMNCs0RC
RRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)Rzq.vdRD:RNDLCRRH#"a11"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloMC5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*n2RR&"RW"&MRH0CCosl'HN5oC[2*UR"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05lMk_DOCD._4U.*4URR+M_klODCD_*ncn+cRR,d.Rb8C02E2R"&RX&"RR0HMCsoC'NHlo5C5[2+4*;U2
RRRRRRRRRRRRLRRCMoH
RRRRRRRRRRRRzRR)dqv.RR:Xv)qdU.X1RR
RRRRRRRRRRRRRbRRFRs0lRNb5=7R>MRH_osC5[U*+8(RF0IMF*RU[R2,q=jR>FRDI8_N8js52q,R4>R=RIDF_8N8s254,.RqRR=>D_FINs885,.2
RRRRRRRRRRRRRRRRRRRRRRRRqRRd>R=RIDF_8N8s25d,cRqRR=>D_FINs885,c2RRW =I>RsC0_M._d,BRWp=iR>pRBim,RRR=>0_lbU._d52[2;S
SS#SN#MHoRV:RFHsR[MRHR8(RF0IMFRRjoCCMsCN0
SSSSFRRkL0_kd#_.k5MlC_ODdD_.*,U[[+H2=R<Rb0l_dU_.25[52H[;R
RRRRRRRRRRRRRRRRRF_k0s5CoU+*[HR[2<F=RkL0_kd#_.k5MlC_ODdD_.*,U[[+H2ERIC5MRF_k0CdM_.RR='24'R#CDCZR''R;
RRRRRRRRRRRRRCRRMo8RCsMCNR0CNH##o
M;RRRRRRRRRRRRCRM8oCCMsCN0RUz.;S
SCRM8oCCMsCN0REzO	0_o6S;
SEzO	R_M:VRHRH5I8R0E<2RURMoCC0sNCR
RRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqz)vRd.:NRDLRCDH"#R1"1aRH&RMo0CCHs'lCNo58IH0RE2&7R""RR&HCM0o'CsHolNCk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*2ncR"&RW&"RR0HMCsoC'NHlojC52RR&"R "&MRH0CCosl'HN5oCo_C0C_M880CbEk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*Rnc+.Rd,CR8b20E2RR&"RX"&MRH0CCosl'HN5oCU
2;RRRRRRRRRRRRLHCoMS
SRRRRzv)qd:.RRqX)vXd.US1
SRSRRFRbsl0RN5bR7>R=R8bN5_HMs5CoI0H8ER-48MFI0IFRHE80-LD#_8IH0,E2RRU,D_#LI0H8E2-4,jRqRR=>D_FINs885,j2
SSSSRSSRRq4=D>RFNI_858s4R2,q=.R>FRDI8_N8.s52q,Rd>R=RIDF_8N8s25d,cRqRR=>D_FINs885,c2RRW =I>RsC0_M._d,BRWp=iR>pRBiS,
SSSSSmRRRR=>0_lbU._d52j2;S
SS#SN#MHoRV:RFHsR[MRHR8IH04E-RI8FMR0FjCRoMNCs0SC
SRSSR0Fk_#Lk_5d.M_klODCD_,d.HR[2<0=RlUb__5d.jH25[
2;RRRRRRRRRRRRRRRRRkRF0C_so[5H2=R<R0Fk_#Lk_5d.M_klODCD_,d.HR[2IMECRk5F0M_C_Rd.=4R''C2RDR#C';Z'
SSSS8CMRMoCC0sNC#RN#MHo;S
SCRM8oCCMsCN0REzO	;_M
CSSMo8RCsMCNR0Cz	OE_
U;SOSzEc	_RH:RVIR5HE80_sNsN.$52RR>jo2RCsMCN
0CRRRRRRRRz_.ccRR:H5VRI0H8E=R>RRc2oCCMsCN0
RRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVzv)qd:.RRLDNCHDR#1R"1Ra"&MRH0CCosl'HN5oCI0H8E&2RR""7RH&RMo0CCHs'lCNo5lMk_DOCD._4U.*4URR+M_klODCD_*ncnRc2&WR""RR&HCM0o'CsHolNC25jR"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05lMk_DOCD._4U.*4URR+M_klODCD_*ncn+cRR,d.Rb8C02E2R"&RX&"RR0HMCsoC'NHlocC52R;
RRRRRRRRRLRRCMoH
RRRRRRRRRRRRqz)vRd.:)RXq.vdXRc1
RRRRRRRRRRRRRRRRsbF0NRlb7R5d>R=R_HMs5CodR2,7=.R>MRH_osC5,.2RR74=H>RMC_so254,jR7RR=>HsM_Cjo52S,
SRSRRRRRRRRRRRRRq=jR>FRDI8_N8js52q,R4>R=RIDF_8N8s254,.RqRR=>D_FINs885,.2
RRRRRRRRRRRRRRRRRRRRRRRRqRRd>R=RIDF_8N8s25d,cRqRR=>D_FINs885,c2RRW =I>RsC0_M._d,BRWp=iR>pRBi
,RSSSSSRSRm=dR>kRF0k_L#._d5lMk_DOCD._d,,d2RRm.=F>RkL0_kd#_.k5MlC_ODdD_.2,.,S
SSSSSR4RmRR=>F_k0L_k#dM.5kOl_C_DDd4.,2m,Rj>R=R0Fk_#Lk_5d.M_klODCD_,d.j;22
RRRRRRRRRRRRRRRR0Fk_osC5Rd2<F=RkL0_kd#_.k5MlC_ODdD_.2,dRCIEMFR5kC0_M._dR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so25.RR<=F_k0L_k#dM.5kOl_C_DDd..,2ERIC5MRF_k0CdM_.RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o52=R<R0Fk_#Lk_5d.M_klODCD_,d.4I2RERCM50Fk__CMd=.RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Coj<2R=kRF0k_L#._d5lMk_DOCD._d,Rj2IMECRk5F0M_C_Rd.=4R''C2RDR#C';Z'
RRRRRRRR8CMRMoCC0sNC.Rzc;_c
RRRRRRRRcz._:dRRRHV58IH0=ERRRd2oCCMsCN0
RRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVzv)qd:.RRLDNCHDR#1R"1Ra"&MRH0CCosl'HN5oCI0H8E&2RR""7RH&RMo0CCHs'lCNo5lMk_DOCD._4U.*4URR+M_klODCD_*ncnRc2&WR""RR&HCM0o'CsHolNC25jR"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05lMk_DOCD._4U.*4URR+M_klODCD_*ncn+cRR,d.Rb8C02E2R"&RX&"RR0HMCsoC'NHlocC52R;
RRRRRRRRRLRRCMoH
RRRRRRRRRRRRqz)vRd.:)RXq.vdXRc1
RRRRRRRRRRRRRRRRsbF0NRlb7R5d>R=R''j,.R7RR=>HsM_C.o527,R4>R=R_HMs5Co4R2,7=jR>MRH_osC5,j2
SSSRRRRRRRRRRRRRjRqRR=>D_FINs885,j2RRq4=D>RFNI_858s4R2,q=.R>FRDI8_N8.s52R,
RRRRRRRRRRRRRRRRRRRRRRRRRRqd=D>RFNI_858sdR2,q=cR>FRDI8_N8cs52W,R >R=R0Is__CMdR.,WiBpRR=>B,piRS
SSSSSRdRmRR=>FMbC,.RmRR=>F_k0L_k#dM.5kOl_C_DDd..,2S,
SSSSSmRR4>R=R0Fk_#Lk_5d.M_klODCD_,d.4R2,m=jR>kRF0k_L#._d5lMk_DOCD._d,2j2;R
RRRRRRRRRRRRRRkRF0C_so25.RR<=F_k0L_k#dM.5kOl_C_DDd..,2ERIC5MRF_k0CdM_.RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o52=R<R0Fk_#Lk_5d.M_klODCD_,d.4I2RERCM50Fk__CMd=.RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Coj<2R=kRF0k_L#._d5lMk_DOCD._d,Rj2IMECRk5F0M_C_Rd.=4R''C2RDR#C';Z'
RRRRRRRR8CMRMoCC0sNC.Rzc;_d
CSSMo8RCsMCNR0Cz	OE_
c;SOSzE.	_RH:RVIR5HE80_sNsN4$52RR>jo2RCsMCN
0CRRRRRRRRzR.c:FRVsRR[H5MRI0H8Es_Ns5N$4-2RRR428MFI0jFRRMoCC0sNCR
RRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqz)vRd.:NRDLRCDH"#R1"1aRH&RMo0CCHs'lCNo58IH0RE2&7R""RR&HCM0o'CsHolNCk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*2ncR"&RW&"RR0HMCsoC'NHloIC5HE80-IU*HE80_sNsNd$52*-.[2-.R"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05lMk_DOCD._4U.*4URR+M_klODCD_*ncn+cRR,d.Rb8C02E2R"&RX&"RR0HMCsoC'NHloIC5HE80-IU*HE80_sNsNd$52*-.[
2;RRRRRRRRRRRRLHCoMR
RRRRRRRRRR)Rzq.vdR):Rq.vdXR.1
RRRRRRRRRRRRRRRRsbF0NRlb7R5j>R=R_HMs5CoI0H8E*-UI0H8Es_Ns5N$d.2-*.[-27,R4>R=R_HMs5CoI0H8E*-UI0H8Es_Ns5N$d.2-*4[-2q,Rj>R=RIDF_8N8s25j,4RqRR=>D_FINs885,42RRq.=D>RFNI_858s.
2,RRRRRRRRRRRRRRRRRRRRRRRRRdRqRR=>D_FINs885,d2RRqc=D>RFNI_858scR2,W= R>sRI0M_C_,d.RpWBi>R=RiBp,jRmRR=>F_k0L_k#dM.5kOl_C_DDdI.,HE80-IU*HE80_sNsNd$52*-.[2-.,S
SSSSSR4RmRR=>F_k0L_k#dM.5kOl_C_DDdI.,HE80-IU*HE80_sNsNd$52*-.[2-42R;
RRRRRRRRRRRRRFRRks0_CIo5HE80-IU*HE80_sNsNd$52*-.[2-4RR<=F_k0L_k#dM.5kOl_C_DDdI.,HE80-IU*HE80_sNsNd$52*-.[2-4RCIEMFR5kC0_M._dR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soH5I8-0EUH*I8_0ENNss$25d-[.*-R.2<F=RkL0_kd#_.k5MlC_ODdD_.H,I8-0EUH*I8_0ENNss$25d-[.*-R.2IMECRk5F0M_C_Rd.=4R''C2RDR#C';Z'
RRRRRRRR8CMRMoCC0sNC.RzcS;
S8CMRMoCC0sNCORzE.	_;S
Sz	OE_:4RRRHV58IH0NE_s$sN5Rj2>2RjRMoCC0sNCR
RRRRRR.RzcRR:H5VRI0H8EFRl8RRU=2R4RMoCC0sNCR
RRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqz)vRd.:NRDLRCDH"#R1"1aRH&RMo0CCHs'lCNo58IH0RE2&7R""RR&HCM0o'CsHolNCk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*2ncR"&RW&"RR0HMCsoC'NHlojC52RR&"R "&MRH0CCosl'HN5oCo_C0C_M880CbEk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*Rnc+.Rd,CR8b20E2RR&"RX"&MRH0CCosl'HN5oC4
2;RRRRRRRRRRRRLHCoMR
RRRRRRRRRR)Rzq.vdR):Rq.vdXR41
RRRRRRRRRRRRRRRRsbF0NRlb7R5RR=>HsM_Cjo52q,Rj>R=RIDF_8N8s25j,4RqRR=>D_FINs885,42RRq.=D>RFNI_858s.
2,RRRRRRRRRRRRRRRRRRRRRRRRRdRqRR=>D_FINs885,d2RRqc=D>RFNI_858scR2,W= R>sRI0M_C_,d.RpWBi>R=RiBp,RRm=F>RkL0_kd#_.k5MlC_ODdD_.2,j2R;
RRRRRRRRRRRRRFRRks0_Cjo52=R<R0Fk_#Lk_5d.M_klODCD_,d.jI2RERCM50Fk__CMd=.RR''42DRC#'CRZ
';RRRRRRRRCRM8oCCMsCN0Rcz.;S
SCRM8oCCMsCN0REzO	;_4
RRRR8CMRMoCC0sNC.Rz4R;RRRRRRRRR
R
RR-R-RMtCC0sNCRRN4InRFRs88bCCRv)qRDOCDVRHRbNbssFbHCN0RRRRRRRRRRRRR
RRRRRRzR.6:VRHRk5MlC_OD4D_nRR=4o2RCsMCN
0CRRRR-Q-RVNR58I8sHE80R6>R2CRMC08RFsROCCN0RHIs0CCRMDNLCMRN8kRF00bkRNCMLRDC#CCDOD0RFOoH
RRRRRRRRnz.NRR:H5VRNs88I0H8ERR>(MRN8kRMlC_ODnD_cRR=4MRN8kRMlC_ODdD_.RR=4o2RCsMCN
0CRRRRRRRRRRRRRRRRF_k0C4M_n=R<R''4RCIEM5R5Ns8_CNo58I8sHE80-84RF0IMF2R(RM=RkOl_C_DD42.UR8NMR85N_osC5Rn2=4R''N2RM58RNs8_C6o52RR='24'R8NMR85N_osC5Rc2=jR''R22CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C_R4n<W=R ERIC5MR5_N8s5CoNs88I0H8ER-48MFI0(FR2RR=M_klODCD_U4.2MRN8NR58C_so25nR'=R4R'2NRM85_N8s5Co6=2RR''42MRN8NR58C_so25cR'=Rj2'2R#CDCjR''R;
RRRRRCRRMo8RCsMCNR0CzN.n;R
RRRRRR.Rzn:LRRRHV58N8s8IH0>ERRN(RMM8RkOl_C_DDn=cRRN4RMM8RkOl_C_DDd=.RRRj2oCCMsCN0
RRRRRRRRRRRRRRRR0Fk__CM4<nR=4R''ERIC5MR5_N8s5CoNs88I0H8ER-48MFI0(FR2RR=M_klODCD_U4.2MRN8NR58C_so25nR'=R4R'2NRM85_N8s5Co6=2RR''j2MRN8NR58C_so25cR'=Rj2'2R#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_Mn_4RR<=WI RERCM585N_osC58N8s8IH04E-RI8FMR0F(=2RRlMk_DOCD._4UN2RM58RNs8_Cno52RR='24'R8NMR85N_osC5R62=jR''N2RM58RNs8_Cco52RR='2j'2DRC#'CRj
';RRRRRRRRCRM8oCCMsCN0Rnz.LR;
RRRRRzRR.RnO:VRHR85N8HsI8R0E>RR(NRM8M_klODCD_Rnc=RRjNRM8M_klODCD_Rd.=2R4RMoCC0sNCR
RRRRRRRRRRRRRRkRF0M_C_R4n<'=R4I'RERCM585N_osC58N8s8IH04E-RI8FMR0F(=2RRlMk_DOCD._4UN2RM58RNs8_Cno52RR='2j'R8NMR85N_osC5R62=4R''N2RM58RNs8_Cco52RR='2j'2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0C4M_n=R<RRW IMECRN558C_so85N8HsI8-0E4FR8IFM0RR(2=kRMlC_OD4D_.RU2NRM85_N8s5Con=2RR''j2MRN8NR58C_so256R'=R4R'2NRM85_N8s5Coc=2RR''j2C2RDR#C';j'
RRRRRRRR8CMRMoCC0sNC.Rzn
O;RRRRRRRRz8.nRH:RVNR58I8sHE80R(>RR8NMRlMk_DOCDc_nRj=RR8NMRlMk_DOCD._dRj=R2CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_Mn_4RR<='R4'IMECRN558C_so85N8HsI8-0E4FR8IFM0RR(2=kRMlC_OD4D_.RU2NRM85_N8s5Con=2RR''j2MRN8NR58C_so256R'=RjR'2NRM85_N8s5Coc=2RR''j2C2RDR#C';j'
RRRRRRRRRRRRRRRR0Is__CM4<nR= RWRCIEM5R5Ns8_CNo58I8sHE80-84RF0IMF2R(RM=RkOl_C_DD42.UR8NMR85N_osC5Rn2=jR''N2RM58RNs8_C6o52RR='2j'R8NMR85N_osC5Rc2=jR''R22CCD#R''j;R
RRRRRRMRC8CRoMNCs0zCR.;n8
RRRRRRRRnz.CRR:H5VRNs88I0H8ERR=(MRN8kRMlC_ODnD_cRR=4MRN8kRMlC_ODdD_.RR=4o2RCsMCN
0CRRRRRRRRRRRRRRRRF_k0C4M_n=R<R''4RCIEM5R5Ns8_Cno52RR='24'R8NMR85N_osC5R62=4R''N2RM58RNs8_Cco52RR='2j'2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0C4M_n=R<RRW IMECRN558C_so25nR'=R4R'2NRM85_N8s5Co6=2RR''42MRN85RRNs8_Cco52RR='2j'2DRC#'CRj
';RRRRRRRRCRM8oCCMsCN0Rnz.CR;
RRRRRzRR.RnV:VRHR85N8HsI8R0E=RR(NRM8M_klODCD_Rnc=RR4NRM8M_klODCD_Rd.=2RjRMoCC0sNCR
RRRRRRRRRRRRRRkRF0M_C_R4n<'=R4I'RERCM585N_osC5Rn2=4R''N2RM58RNs8_C6o52RR='2j'R8NMR85N_osC5Rc2=jR''R22CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C_R4n<W=R ERIC5MR5_N8s5Con=2RR''42MRN8NR58C_so256R'=RjR'2NRM85_N8s5Coc=2RR''j2C2RDR#C';j'
RRRRRRRR8CMRMoCC0sNC.Rzn
V;RRRRRRRRzo.nRH:RVNR58I8sHE80Rn=RR8NMRlMk_DOCDc_nRj=RR8NMRlMk_DOCD._dR4=R2CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_Mn_4RR<='R4'IMECRN558C_so256R'=R4R'2NRM85_N8s5Coc=2RR''j2C2RDR#C';j'
RRRRRRRRRRRRRRRR0Is__CM4<nR= RWRCIEM5R5Ns8_C6o52RR='24'R8NMR85N_osC5Rc2=jR''R22CCD#R''j;R
RRRRRRMRC8CRoMNCs0zCR.;no
RRRRRRRRnz.ERR:H5VRNs88I0H8ERR=6MRN8kRMlC_ODdD_.=R/RR42oCCMsCN0
RRRRRRRRRRRRRRRR0Fk__CM4<nR=4R''ERIC5MR5_N8s5CoNs88I0H8ER-48MFI0cFR2RR=M_klODCD_2d.2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0C4M_n=R<RRW IMECRN558C_so85N8HsI8-0E4FR8IFM0RRc2=kRMlC_ODdD_.R22CCD#R''j;R
RRRRRRMRC8CRoMNCs0zCR.;nE
RRRRR--Q5VRNs88I0H8E=R<RR62MIFRsCH0RNCMLRDCFFsRkk0b0MRCNCLDRD#CCRO0DHFoOCRMC88C
RRRRRRRR(z.RH:RVNR58I8sHE80RR<=co2RCsMCN
0CRRRRRRRRRRRRRRRRF_k0C4M_n=R<R''4;R
RRRRRRRRRRRRRRsRI0M_C_R4n<W=R R;
RRRRRCRRMo8RCsMCNR0Cz;.(
RRRRR--tCCMsCN0RC0ERv)qRDOCDMRN8sR0H0-#N
0CSRRRREzO	R_U:VRHRH5I8_0ENNss$25dRj>R2CRoMNCs0SC
SEzO	C_D6RR:H5VRI0H8E=R>RIU*HE80_sNsNd$52MRN8HRI8R0E>U=R2CRoMNCs0RC
RRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)Rzqnv4RD:RNDLCRRH#"a11"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloMC5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*nRM+RkOl_C_DDdd.*.&2RR""WRH&RMo0CCHs'lCNo58IH0-ERRLD#_8IH0RE2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50EM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*cRR+M_klODCD_*d.d+.RR,4nRb8C02E2R"&RX&"RR0HMCsoC'NHloIC5HE80RD-R#IL_HE80RU+R2R;
RRRRRRRRRLRRCMoH
RSSRzRR)4qvnRR:Xv)q4UnX1S
SSRRRRsbF0NRlb7R5RR=>b5N8HsM_CIo5HE80-84RF0IMFHRI8-0ED_#LI0H8ER2,UD,R#IL_HE80-,42RRqj=D>RFNI_858sj
2,SSSSSRSRq=4R>FRDI8_N84s52q,R.>R=RIDF_8N8s25.,dRqRR=>D_FINs885,d2RRW =I>RsC0_Mn_4,BRWp=iR>pRBiS,
SSSSSmRRRR=>0_lbUn_452j2;S
SS#SN#MHoRV:RFHsR[MRHR8IH04E-RI8FMR0FI0H8E#-DLH_I8R0EoCCMsCN0
SSSSFRRkL0_k4#_nk5MlC_OD4D_n[,H2=R<Rb0l_4U_n25j5-H[I0H8E#+DLH_I820E;R
RRRRRRRRRRRRRRRRRF_k0s5CoHR[2<F=RkL0_k4#_nk5MlC_OD4D_n[,H2ERIC5MRF_k0C4M_nRR='24'R#CDCZR''S;
SCSSMo8RCsMCNR0CNH##o
M;RRRRRRRRRRRRzR.U:FRVsRR[HIMRHE80_sNsNd$52R-48MFI04FRRMoCC0sNCR
RRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FzVR)4qvnRR:DCNLD#RHR1"1a&"RR0HMCsoC'NHloIC5HE802RR&"R7"&MRH0CCosl'HN5oCM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*cRR+M_klODCD_*d.dR.2&WR""RR&HCM0o'CsHolNCH5I8R0E-#RDLH_I8R0E-*R[U&2RR"" RH&RMo0CCHs'lCNo50oC_8CM_b8C0ME5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*nRM+RkOl_C_DDdd.*.RR+4Rn,80CbER22&XR""RR&HCM0o'CsHolNCH5I8R0E-#RDLH_I8R0E-[R5-*42U
2;RRRRRRRRRRRRRCRLo
HMRRRRRRRRRRRRR)Rzqnv4RX:R)4qvn1XURR
RRRRRRRRRRRRRRFRbsl0RN5bR7>R=R_HMs5CoI0H8E#-DLH_I8-0EU+*[(FR8IFM0R8IH0DE-#IL_HE80-[U*2q,Rj>R=RIDF_8N8s25j,4RqRR=>D_FINs885,42RRq.=D>RFNI_858s.
2,RRRRRRRRRRRRRRRRRRRRRRRRRdRqRR=>D_FINs885,d2RRW =I>RsC0_Mn_4,BRWp=iR>pRBim,RRR=>0_lbUn_452[2;S
SSRRRR#N#HRoM:FRVs[RHRRHM(FR8IFM0RojRCsMCN
0CSSSSRkRF0k_L#n_45lMk_DOCDn_4,8IH0DE-#IL_HE80-[U*+2H[RR<=0_lbUn_455[2H;[2
RRRRRRRRRRRRRRRRFRRks0_CIo5HE80-LD#_8IH0UE-*H[+[<2R=kRF0k_L#n_45lMk_DOCDn_4,8IH0DE-#IL_HE80-[U*+2H[RCIEMFR5kC0_Mn_4R'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRMRC8CRoMNCs0NCR#o#HMR;
RRRRRRRRRCRRMo8RCsMCNR0Cz;.U
CSSMo8RCsMCNR0Cz	OE_6DC;S
Sz	OE_6o0RH:RVIR5HE80RR>=UMRN8HRI8R0ElRF8U=R>RR62oCCMsCN0
RRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVzv)q4:nRRLDNCHDR#1R"1Ra"&MRH0CCosl'HN5oCI0H8E&2RR""7RH&RMo0CCHs'lCNo5lMk_DOCD._4U.*4URR+M_klODCD_*ncn+cRRlMk_DOCD._d*2d.R"&RW&"RR0HMCsoC'NHloIC5HE80RD-R#IL_HE802RR&"R "&MRH0CCosl'HN5oCo_C0C_M880CbEk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*Rnc+kRMlC_ODdD_..*dR4+Rn8,RCEb02&2RR""XRH&RMo0CCHs'lCNo58IH0-ERRLD#_8IH0+ERR;U2
RRRRRRRRRRRRoLCHSM
SRRRRqz)vR4n:)RXqnv4X
U1SRSSRbRRFRs0lRNb5=7R>NRb8M5H_osC58IH04E-RI8FMR0FI0H8E#-DLH_I820E,,RURLD#_8IH04E-2q,Rj>R=RIDF_8N8s25j,S
SSSSSR4RqRR=>D_FINs885,42RRq.=D>RFNI_858s.R2,q=dR>FRDI8_N8ds52W,R >R=R0Is__CM4Rn,WiBpRR=>B,pi
SSSSRSSR=mR>lR0b__U4In5HE80_sNsNd$522-42S;
SNSS#o#HMRR:VRFsHH[RMHRI8-0E4FR8IFM0R8IH0DE-#IL_HE80RMoCC0sNCS
SSRSRF_k0L_k#4Mn5kOl_C_DD4Hn,[<2R=lR0b__U4In5HE80_sNsNd$522-45-H[I0H8E#+DLH_I820E;R
RRRRRRRRRRRRRRRRRF_k0s5CoHR[2<F=RkL0_k4#_nk5MlC_OD4D_n[,H2ERIC5MRF_k0C4M_nRR='24'R#CDCZR''S;
SCSSMo8RCsMCNR0CNH##o
M;RRRRRRRRRRRRzR.U:FRVsRR[HIMRHE80_sNsNd$52R-.8MFI0jFRRMoCC0sNCR
RRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FzVR)4qvnRR:DCNLD#RHR1"1a&"RR0HMCsoC'NHloIC5HE802RR&"R7"&MRH0CCosl'HN5oCM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*cRR+M_klODCD_*d.dR.2&WR""RR&HCM0o'CsHolNC*5[U&2RR"" RH&RMo0CCHs'lCNo50oC_8CM_b8C0ME5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*nRM+RkOl_C_DDdd.*.RR+4Rn,80CbER22&XR""RR&HCM0o'CsHolNC[55+*42U
2;RRRRRRRRRRRRRCRLo
HMRRRRRRRRRRRRR)Rzqnv4RX:R)4qvn1XURR
RRRRRRRRRRRRRRFRbsl0RN5bR7>R=R_HMs5CoU+*[(FR8IFM0R[U*2q,Rj>R=RIDF_8N8s25j,4RqRR=>D_FINs885,42RRq.=D>RFNI_858s.
2,RRRRRRRRRRRRRRRRRRRRRRRRRdRqRR=>D_FINs885,d2RRW =I>RsC0_Mn_4,BRWp=iR>pRBim,RRR=>0_lbUn_452[2;S
SS#SN#MHoRV:RFHsR[MRHR8(RF0IMFRRjoCCMsCN0
SSSSFRRkL0_k4#_nk5MlC_OD4D_n*,U[[+H2=R<Rb0l_4U_n25[52H[;R
RRRRRRRRRRRRRRRRRF_k0s5CoU+*[HR[2<F=RkL0_k4#_nk5MlC_OD4D_n*,U[[+H2ERIC5MRF_k0C4M_nRR='24'R#CDCZR''R;
RRRRRRRRRRRRRCRRMo8RCsMCNR0CNH##o
M;RRRRRRRRRRRRCRM8oCCMsCN0RUz.;S
SCRM8oCCMsCN0REzO	0_o6S;
SEzO	R_M:VRHRH5I8R0E<2RURMoCC0sNCR
RRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqz)vR4n:NRDLRCDH"#R1"1aRH&RMo0CCHs'lCNo58IH0RE2&7R""RR&HCM0o'CsHolNCk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*Rnc+kRMlC_ODdD_..*d2RR&"RW"&MRH0CCosl'HN5oCj&2RR"" RH&RMo0CCHs'lCNo50oC_8CM_b8C0ME5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*nRM+RkOl_C_DDdd.*.RR+4Rn,80CbER22&XR""RR&HCM0o'CsHolNC25U;R
RRRRRRRRRRCRLo
HMSRSRR)Rzqnv4RX:R)4qvn1XU
SSSRRRRb0FsRblNRR57=b>RNH85MC_soH5I8-0E4FR8IFM0R8IH0DE-#IL_HE802U,R,#RDLH_I8-0E4R2,q=jR>FRDI8_N8js52S,
SSSSSqRR4>R=RIDF_8N8s254,.RqRR=>D_FINs885,.2RRqd=D>RFNI_858sdR2,W= R>sRI0M_C_,4nRpWBi>R=RiBp,S
SSSSSRRRm=0>RlUb__54nj;22
SSSS#N#HRoM:FRVs[RHRRHMI0H8ER-48MFI0jFRRMoCC0sNCS
SSRSRF_k0L_k#4Mn5kOl_C_DD4Hn,[<2R=lR0b__U4jn52[5H2R;
RRRRRRRRRRRRRRRRR0Fk_osC52H[RR<=F_k0L_k#4Mn5kOl_C_DD4Hn,[I2RERCM50Fk__CM4=nRR''42DRC#'CRZ
';SSSSCRM8oCCMsCN0R#N#H;oM
CSSMo8RCsMCNR0Cz	OE_
M;SMSC8CRoMNCs0zCRO_E	US;
SEzO	R_c:VRHRH5I8_0ENNss$25.Rj>R2CRoMNCs0RC
RRRRRzRR.cg_RH:RVIR5HE80RR>=co2RCsMCN
0CRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FzVR)4qvnRR:DCNLD#RHR1"1a&"RR0HMCsoC'NHloIC5HE802RR&"R7"&MRH0CCosl'HN5oCM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*cRR+M_klODCD_*d.dR.2&WR""RR&HCM0o'CsHolNC25jR"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05lMk_DOCD._4U.*4URR+M_klODCD_*ncn+cRRlMk_DOCD._d*Rd.+nR4,CR8b20E2RR&"RX"&MRH0CCosl'HN5oCc
2;RRRRRRRRRRRRLHCoMR
RRRRRRRRRR)Rzqnv4R):Rqnv4XRc1
RRRRRRRRRRRRRRRRsbF0NRlb7R5d>R=R_HMs5CodR2,7=.R>MRH_osC5,.2RR74=H>RMC_so254,jR7RR=>HsM_Cjo52S,
SRSRRRRRRRRRRRRRq=jR>FRDI8_N8js52q,R4>R=RIDF_8N8s254,.RqRR=>D_FINs885,.2
RRRRRRRRRRRRRRRRRRRRRRRRqRRd>R=RIDF_8N8s25d, RWRR=>I_s0C4M_nW,RBRpi=B>RpRi,
SSSSRSSRRmd=F>RkL0_k4#_nk5MlC_OD4D_n2,d,.RmRR=>F_k0L_k#4Mn5kOl_C_DD4.n,2S,
SSSSSmRR4>R=R0Fk_#Lk_54nM_klODCD_,4n4R2,m=jR>kRF0k_L#n_45lMk_DOCDn_4,2j2;R
RRRRRRRRRRRRRRkRF0C_so25dRR<=F_k0L_k#4Mn5kOl_C_DD4dn,2ERIC5MRF_k0C4M_nRR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C.o52=R<R0Fk_#Lk_54nM_klODCD_,4n.I2RERCM50Fk__CM4=nRR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4<2R=kRF0k_L#n_45lMk_DOCDn_4,R42IMECRk5F0M_C_R4n=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5Rj2<F=RkL0_k4#_nk5MlC_OD4D_n2,jRCIEMFR5kC0_Mn_4R'=R4R'2CCD#R''Z;R
RRRRRRMRC8CRoMNCs0zCR.cg_;R
RRRRRR.RzgR_d:VRHRH5I8R0E=2RdRMoCC0sNCR
RRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqz)vR4n:NRDLRCDH"#R1"1aRH&RMo0CCHs'lCNo58IH0RE2&7R""RR&HCM0o'CsHolNCk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*Rnc+kRMlC_ODdD_..*d2RR&"RW"&MRH0CCosl'HN5oCj&2RR"" RH&RMo0CCHs'lCNo50oC_8CM_b8C0ME5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*nRM+RkOl_C_DDdd.*.RR+4Rn,80CbER22&XR""RR&HCM0o'CsHolNC25c;R
RRRRRRRRRRCRLo
HMRRRRRRRRRRRRzv)q4:nRRv)q4cnX1RR
RRRRRRRRRRRRRbRRFRs0lRNb5R7d='>RjR',7=.R>MRH_osC5,.2RR74=H>RMC_so254,jR7RR=>HsM_Cjo52S,
SRSRRRRRRRRRRRRRq=jR>FRDI8_N8js52q,R4>R=RIDF_8N8s254,.RqRR=>D_FINs885,.2
RRRRRRRRRRRRRRRRRRRRRRRRqRRd>R=RIDF_8N8s25d, RWRR=>I_s0C4M_nW,RBRpi=B>RpRi,
SSSSRSSRRmd=F>Rb,CMRRm.=F>RkL0_k4#_nk5MlC_OD4D_n2,.,S
SSSSSR4RmRR=>F_k0L_k#4Mn5kOl_C_DD44n,2m,Rj>R=R0Fk_#Lk_54nM_klODCD_,4nj;22
RRRRRRRRRRRRRRRR0Fk_osC5R.2<F=RkL0_k4#_nk5MlC_OD4D_n2,.RCIEMFR5kC0_Mn_4R'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so254RR<=F_k0L_k#4Mn5kOl_C_DD44n,2ERIC5MRF_k0C4M_nRR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cjo52=R<R0Fk_#Lk_54nM_klODCD_,4njI2RERCM50Fk__CM4=nRR''42DRC#'CRZ
';RRRRRRRRCRM8oCCMsCN0Rgz._
d;SMSC8CRoMNCs0zCRO_E	cS;
SEzO	R_.:VRHRH5I8_0ENNss$254Rj>R2CRoMNCs0RC
RRRRRzRRd:jRRsVFRH[RMIR5HE80_sNsN4$52RR-482RF0IMFRRjoCCMsCN0
RRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVzv)q4:nRRLDNCHDR#1R"1Ra"&MRH0CCosl'HN5oCI0H8E&2RR""7RH&RMo0CCHs'lCNo5lMk_DOCD._4U.*4URR+M_klODCD_*ncn+cRRlMk_DOCD._d*2d.R"&RW&"RR0HMCsoC'NHloIC5HE80-IU*HE80_sNsNd$52*-.[2-.R"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05lMk_DOCD._4U.*4URR+M_klODCD_*ncn+cRRlMk_DOCD._d*Rd.+nR4,CR8b20E2RR&"RX"&MRH0CCosl'HN5oCI0H8E*-UI0H8Es_Ns5N$d.2-*;[2
RRRRRRRRRRRRoLCHRM
RRRRRRRRRzRR)4qvnRR:)4qvn1X.RR
RRRRRRRRRRRRRRFRbsl0RN5bR7=jR>MRH_osC58IH0UE-*8IH0NE_s$sN5-d2.-*[.R2,7=4R>MRH_osC58IH0UE-*8IH0NE_s$sN5-d2.-*[4R2,q=jR>FRDI8_N8js52q,R4>R=RIDF_8N8s254,.RqRR=>D_FINs885,.2
RRRRRRRRRRRRRRRRRRRRRRRRqRRd>R=RIDF_8N8s25d, RWRR=>I_s0C4M_nW,RBRpi=B>RpRi,m=jR>kRF0k_L#n_45lMk_DOCDn_4,8IH0UE-*8IH0NE_s$sN5-d2.-*[.
2,SSSSSRSRm=4R>kRF0k_L#n_45lMk_DOCDn_4,8IH0UE-*8IH0NE_s$sN5-d2.-*[4;22
RRRRRRRRRRRRRRRR0Fk_osC58IH0UE-*8IH0NE_s$sN5-d2.-*[4<2R=kRF0k_L#n_45lMk_DOCDn_4,8IH0UE-*8IH0NE_s$sN5-d2.-*[4I2RERCM50Fk__CM4=nRR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5CoI0H8E*-UI0H8Es_Ns5N$d.2-*.[-2=R<R0Fk_#Lk_54nM_klODCD_,4nI0H8E*-UI0H8Es_Ns5N$d.2-*.[-2ERIC5MRF_k0C4M_nRR='24'R#CDCZR''R;
RRRRRCRRMo8RCsMCNR0Cz;dj
CSSMo8RCsMCNR0Cz	OE_
.;SOSzE4	_RH:RVIR5HE80_sNsNj$52RR>jo2RCsMCN
0CRRRRRRRRzRd4:VRHRH5I8R0ElRF8URR=4o2RCsMCN
0CRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FzVR)4qvnRR:DCNLD#RHR1"1a&"RR0HMCsoC'NHloIC5HE802RR&"R7"&MRH0CCosl'HN5oCM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*cRR+M_klODCD_*d.dR.2&WR""RR&HCM0o'CsHolNC25jR"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05lMk_DOCD._4U.*4URR+M_klODCD_*ncn+cRRlMk_DOCD._d*Rd.+nR4,CR8b20E2RR&"RX"&MRH0CCosl'HN5oC4
2;RRRRRRRRRRRRLHCoMR
RRRRRRRRRR)Rzqnv4R):Rqnv4XR41
RRRRRRRRRRRRRRRRsbF0NRlb7R5RR=>HsM_Cjo52q,Rj>R=RIDF_8N8s25j,4RqRR=>D_FINs885,42RRq.=D>RFNI_858s.
2,RRRRRRRRRRRRRRRRRRRRRRRRRdRqRR=>D_FINs885,d2RRW =I>RsC0_Mn_4,BRWp=iR>pRBim,RRR=>F_k0L_k#4Mn5kOl_C_DD4jn,2
2;RRRRRRRRRRRRRRRRF_k0s5Coj<2R=kRF0k_L#n_45lMk_DOCDn_4,Rj2IMECRk5F0M_C_R4n=4R''C2RDR#C';Z'
RRRRRRRR8CMRMoCC0sNCdRz4S;
S8CMRMoCC0sNCORzE4	_;R
RRCRRMo8RCsMCNR0Cz;.6RRRRRRRRR
R
CRM8NEsOHO0C0CksRD#CC_O0s;Nl
