--*****************************************************
@Ea--HC0D:RRRR_#LH_OCObFlFMMC0D#_OE3P8-R
-#7CH:oMR#RRLO_HCF_OlMbFC#M0_3DOPRE8
q--kF0EsR:RRD[oF
Mo-k-wMHO0FRM:BbFlFMMC0F#RVER0CERb$O#HNpDRFOoHRDBCD-
-BbFlN:M$RHR1DFHOMkADCCRaOFEMDHFoCR#,Q3MO
Q--h:QaRRRRRLwCR,4URj.jU-
-*****************************************************D*
HNLssH$RCRCC;#
kCCRHC#C30D8_FOoH_n44cD3ND
;
b	NONRoC#HL_OOC_FFlbM0CM#O_DR
H#
lOFbCFMMt0RhR7
RRRRRRRRRsbF0
5RRRRRRRRRRRRRRRRRYRR:FRk0R8#0_oDFH
ORRRRRRRRRRRRRRRRR2C;
MO8RFFlbM0CM;O

FFlbM0CMRBeB
RRRRRRRRbRRF5s0RR
RRRRRRRRRRRRRRRRY:kRF0#RR0D8_FOoHRR
RRRRRRRRRRRRRR;R2
8CMRlOFbCFMM
0;
F
OlMbFCRM0DHFoOC_ODRD
RRRRRRRRRsbF0R5
RRRRRRRRRORRN$ss_0FkRF:Rk#0R0D8_FOoH;R
RRRRRRRRRRORD_0FkRRRR:kRF00R#8F_Do;HO
RRRRRRRRR
RRRRRRRRRRNROs_s$H:MRRMRHR8#0_oDFH
O;RRRRRRRRRRRRORD	RRRRRR:RH#MR0D8_FOoH;R
RRRRRRRRRRDRO	RLRR:RRRMRHR8#0_oDFH
O;RRRRRRRRRRRRHRMjRRRRRR:RH#MR0D8_FOoH;R
RRRRRRRRRRMRH4RRRR:RRRMRHR8#0_oDFH
O;RRRRRRRRRRRRHRM.RRRRRR:RH#MR0D8_FOoH;R
RRRRRRRRRRMRHdRRRR:RRRMRHR8#0_oDFH
O;RRRRRRRRRRRRbosFRRRRRR:RH#MR0D8_FOoH;R
RRRRRRRRRRkRbsR#0R:RRRMRHR8#0_oDFH
O;RRRRRRRRRRRR#R_sRRRRRR:RH#MR0D8_FOoH;R
RRRRRRRRRRLROHR0RR:RRRMRHR8#0_oDFHPO_CFO0sj5.RI8FMR0FjR2
RRRRRRRRR2RR;M
C8FROlMbFC;M0
F
OlMbFCRM0pHFoODBCDR
RRRRRRRRRoCCMsRHO5RR
RRRRRRRRRSSSS S1Tm_v7R R:HRL0C_POs0F58dRF0IMF2RjRR:="jjjj
";RRRRRRRRRRRRSSSSBh_mRRRRRRR:LRH0:'=RjR';
RRRRRRRRRRRRSSSSapz_QQha:RRR0LH_OPC05Fs486RF0IMF2RjRR:=Xj"jj
j"RRRRRRRRRRRRRRRRRRR2;R
RRRRRRRRRb0Fs5RR
RRRRRRRRRRRRRORRN$ss_0FkRF:RkR0R#_08DHFoO
R;RRRRRRRRRRRRRRRRDFO_kR0RRRR:FRk0R8#0_oDFH;OR
R
RRRRRRRRRRRRRRNROs_s$HRMR:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRDRO	RRRRRRR:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRDRO	RLRRRRR:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRMRHjRRRRRRR:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRMRH4RRRRRRR:MRHR0R#8F_DoRHO;RR
RRRRRRRRRRRRRHRRMR.RRRRRRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRRHRRMRdRRRRRRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRR#RR_RsRRRRRRH:RM#RR0D8_FOoHRR
RRRRRRRRRRRRRR;R2
8CMRlOFbCFMM
0;
lOFbCFMMQ0RhRe
RRRRRRRRRsbF0
5RRRRRRRRRRRRRRRRRQ:RRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRR:mRR0FkR0R#8F_DoRHO
RRRRRRRRRRRRRRRR
2;CRM8ObFlFMMC0
;
ObFlFMMC0MRHPP_E0R
RRRRRRRRRb0Fs5RR
RRRRRRRRRRRRRQRRRRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRRmRR:FRk0R8#0_oDFH
ORRRRRRRRRRRRRRRRR2C;
MO8RFFlbM0CM;O

FFlbM0CMRsOFCV8VsR
RRRRRRRRRb0Fs5R
RRRRRRRRRRRRJRRRRRRR:FRk0#_08DHFoOR;
RRRRR
RRRRRRRRRRRRRR8RRRRRRR:MRHR8#0_oDFH
O;RRRRRRRRRRRRb#ks0RRR:MRHR8#0_oDFH
O;RRRRRRRRRRRR1R_)RRRR:MRHR8#0_oDFH
O;RRRRRRRRRRRRORD	RRRR:MRHR8#0_oDFH
O;RRRRRRRRRRRROLD	RRRR:MRHR8#0_oDFH
O;RRRRRRRRRRRRO0LHRRRR:MRHR8#0_oDFHPO_CFO0sR548MFI0jFR2R
RRRRRRRRRR;R2
8CMRlOFbCFMM
0;
lOFbCFMMO0RDck0
RRRRRRRRbRRF5s0
RRRRRRRRRRRR0DkcRR:FRk0#_08DHFoOR;
RRRRR
RRRRRRRRRRRRRRHRMjRH:RM0R#8F_Do;HO
RRRRRRRRRRRR4HMRRR:H#MR0D8_FOoH;R
RRRRRRRRRRMRH.:RRRRHM#_08DHFoOR;
RRRRRRRRRHRRMRdR:MRHR8#0_oDFH
O;RRRRRRRRRRRRHLMjRH:RM0R#8F_Do;HO
RRRRRRRRRRRR4HMLRR:H#MR0D8_FOoH;R
RRRRRRRRRRMRH.:LRRRHM#_08DHFoOR;
RRRRRRRRRHRRMRdL:MRHR8#0_oDFH
O;RRRRRRRRRRRRO0LHRH:RM0R#8F_Do_HOP0COF4s56FR8IFM0R
j2RRRRRRRRRRRR2C;
MO8RFFlbM0CM;O

FFlbM0CMRsONsD$_FOoH
RRRRRRRRbRRF5s0
RRRRRRRRRRRRkOF0RR:FRk0#_08DHFoOR;
RRRRR
RRRRRRRRRRRRRROsNs$M_HRRR:H#MR0D8_FOoH;R
RRRRRRRRRRRRNRRRRRRRR:MRHR8#0_oDFH
O;RRRRRRRRRRRRNN_LsRRRRRR:H#MR0D8_FOoH;R
RRRRRRRRRRRRLRRRRRRRR:MRHR8#0_oDFH
O;RRRRRRRRRRRRLN_LsRRRRRR:H#MR0D8_FOoH;R
RRRRRRRRRRoRP_RCMRRRR:MRHR8#0_oDFHRO
RRRRRRRRR2RR;M
C8FROlMbFC;M0
F
OlMbFCRM0Fk_lGR
RRRRRRRRRb0Fs5R
RRRRRRRRRRRRmR:RRR0FkR8#0_oDFH
O;RRRRRRRR
RRRRRRRRRRRRjHMRRR:H#MR0D8_FOoH;R
RRRRRRRRRRMRH4:RRRRHM#_08DHFoOR;
RRRRRRRRRORRLRH0:MRHR8#0_oDFH
O;RRRRRRRRRRRRbosFRH:RM0R#8F_Do
HORRRRRRRRRRRR2C;
MO8RFFlbM0CM;O

FFlbM0CMR7qh.R
RRRRRRRRRb0Fs5RR
RRRRRRRRRRRRRqRRRRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRRA:RRRRHMR8#0_oDFH;OR
R
RRRRRRRRRRRRRRRRmRF:RkR0R#_08DHFoORR
RRRRRRRRRRRRR2RR;M
C8FROlMbFC;M0
F
OlMbFCRM0BvD	kRG
RRRRRRRRRsbF0
5RRRRRRRRRRRRRRRRRQ:RRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRRmR:kRF0#RR0D8_FOoHRR
RRRRRRRRRRRRRR;R2
8CMRlOFbCFMM
0;
lOFbCFMM10R)Gvk
RRRRRRRRbRRF5s0RR
RRRRRRRRRRRRRRRRQRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRRmRRRRR:FRk0R8#0_oDFH
ORRRRRRRRRRRRRRRRR2C;
MO8RFFlbM0CM;O

FFlbM0CMRLtD.OpFNkDvGR
RRRRRRRRRb0Fs5RR
RRRRRRRRRRRRRQRRRRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRRm:RRR0FkR0R#8F_DoRHO
RRRRRRRRRRRRRRRR
2;CRM8ObFlFMMC0
;
ObFlFMMC0 RBv
kGRRRRRRRRRFRbsR05
RRRRRRRRRRRRRRRRRQR:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRRRmRF:RkR0R#_08DHFoORR
RRRRRRRRRRRRR2RR;M
C8FROlMbFC;M0
F
OlMbFCRM01MbN4k.vGR
RRRRRRRRRb0Fs5RR
RRRRRRRRRRRRRQRRRRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRRm:RRR0FkR0R#8F_DoRHO
RRRRRRRRRRRRRRRR
2;CRM8ObFlFMMC0
;
ObFlFMMC0bR14F.0cR
RRRRRRRRRb0Fs5RR
RRRRRRRRRRRRRQRRRRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRRm:RRR0FkR0R#8F_DoRHO
RRRRRRRRRRRRRRRR
2;CRM8ObFlFMMC0
;
ObFlFMMC08Rms
PcRRRRRRRRRFRbsR05
RRRRRRRRRRRRRRRRRQR:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRRRmRF:RkR0R#_08DHFoORR
RRRRRRRRRRRRR2RR;M
C8FROlMbFC;M0
F
OlMbFCRM0mP8s4R.
RRRRRRRRRsbF0
5RRRRRRRRRRRRRRRRRQ:RRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRRmR:kRF0#RR0D8_FOoHRR
RRRRRRRRRRRRRR;R2
8CMRlOFbCFMM
0;
lOFbCFMMp0RFDONv
kGRRRRRRRRRFRbsR05
RRRRRRRRRRRRRRRRRQR:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRRRmRF:RkR0R#_08DHFoORR
RRRRRRRRRRRRR2RR;M
C8FROlMbFC;M0
F
OlMbFCRM01MbNcGvk
RRRRRRRRbRRF5s0RR
RRRRRRRRRRRRRRRRQRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRRmRRRRR:FRk0R8#0_oDFH
ORRRRRRRRRRRRRRRRR2C;
MO8RFFlbM0CM;O

FFlbM0CMRvQMkRG
RRRRRRRRRsbF0
5RRRRRRRRRRRRRRRRRQ:RRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRRmR:kRF0#RR0D8_FOoHRR
RRRRRRRRRRRRRR;R2
8CMRlOFbCFMM
0;
lOFbCFMMQ0RFvQMkRG
RRRRRRRRRsbF0
5RRRRRRRRRRRRRRRRRQ:RRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRRmR:kRF0#RR0D8_FOoHRR
RRRRRRRRRRRRRR;R2
8CMRlOFbCFMM
0;
lOFbCFMMo0RHBF.0AsDkRV
RRRRRRRRRsbF0
5RRRRRRRRRRRRRRRRRQ:RRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRRmR:kRF0#RR0D8_FOoHRR
RRRRRRRRRRRRRR;R2
8CMRlOFbCFMM
0;
lOFbCFMMt0RDNFLDGvkRR
RRRRRRRRRb0Fs5RR
RRRRRRRRRRRRRQRRRRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRRm:RRR0FkR0R#8F_DoRHO
RRRRRRRRRRRRRRRR
2;CRM8ObFlFMMC0
;
ObFlFMMC0FRQ1MbNcGvkRR
RRRRRRRRRb0Fs5RR
RRRRRRRRRRRRRQRRRRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRRm:RRR0FkR0R#8F_DoRHO
RRRRRRRRRRRRRRRR
2;CRM8ObFlFMMC0
;
ObFlFMMC0bR1NvMckPG_RR
RRRRRRRRRb0Fs5RR
RRRRRRRRRRRRRQRRRRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRRm:RRR0FkR0R#8F_DoRHO
RRRRRRRRRRRRRRRR
2;CRM8ObFlFMMC0
;
ObFlFMMC0bR1NvMck#G_jR_P
RRRRRRRRbRRF5s0RR
RRRRRRRRRRRRRRRRQRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRRmRRRRR:FRk0R8#0_oDFH
ORRRRRRRRRRRRRRRRR2C;
MO8RFFlbM0CM;O

FFlbM0CMRN1bMkcvG4_#_
PRRRRRRRRRRFRbsR05
RRRRRRRRRRRRRRRRRQR:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRRRmRF:RkR0R#_08DHFoORR
RRRRRRRRRRRRR2RR;M
C8FROlMbFC;M0
F
OlMbFCRM01MbNcGvk__#.PRR
RRRRRRRRRsbF0
5RRRRRRRRRRRRRRRRRQ:RRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRRmR:kRF0#RR0D8_FOoHRR
RRRRRRRRRRRRRR;R2
8CMRlOFbCFMM
0;
lOFbCFMM10RbcNMv_kG#Pd_RR
RRRRRRRRRb0Fs5RR
RRRRRRRRRRRRRQRRRRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRRm:RRR0FkR0R#8F_DoRHO
RRRRRRRRRRRRRRRR
2;CRM8ObFlFMMC0
;
ObFlFMMC0bR1NvMckEG_RR
RRRRRRRRRb0Fs5RR
RRRRRRRRRRRRRQRRRRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRRm:RRR0FkR0R#8F_DoRHO
RRRRRRRRRRRRRRRR
2;CRM8ObFlFMMC0
;
ObFlFMMC0bR1NvMck#G_jR_E
RRRRRRRRbRRF5s0RR
RRRRRRRRRRRRRRRRQRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRRmRRRRR:FRk0R8#0_oDFH
ORRRRRRRRRRRRRRRRR2C;
MO8RFFlbM0CM;O

FFlbM0CMRN1bMkcvG4_#_
ERRRRRRRRRRFRbsR05
RRRRRRRRRRRRRRRRRQR:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRRRmRF:RkR0R#_08DHFoORR
RRRRRRRRRRRRR2RR;M
C8FROlMbFC;M0
F
OlMbFCRM01MbNcGvk__#.ERR
RRRRRRRRRsbF0
5RRRRRRRRRRRRRRRRRQ:RRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRRmR:kRF0#RR0D8_FOoHRR
RRRRRRRRRRRRRR;R2
8CMRlOFbCFMM
0;
lOFbCFMM10RbcNMv_kG#Ed_RR
RRRRRRRRRb0Fs5RR
RRRRRRRRRRRRRQRRRRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRRm:RRR0FkR0R#8F_DoRHO
RRRRRRRRRRRRRRRR
2;CRM8ObFlFMMC0
;
ObFlFMMC0bR1N.M4v_kGERR
RRRRRRRRRsbF0
5RRRRRRRRRRRRRRRRRQ:RRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRRmR:kRF0#RR0D8_FOoHRR
RRRRRRRRRRRRRR;R2
8CMRlOFbCFMM
0;
lOFbCFMM10Rb4NM.Gvk__#jERR
RRRRRRRRRsbF0
5RRRRRRRRRRRRRRRRRQ:RRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRRmR:kRF0#RR0D8_FOoHRR
RRRRRRRRRRRRRR;R2
8CMRlOFbCFMM
0;
lOFbCFMM10Rb4NM.Gvk__#4ERR
RRRRRRRRRsbF0
5RRRRRRRRRRRRRRRRRQ:RRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRRmR:kRF0#RR0D8_FOoHRR
RRRRRRRRRRRRRR;R2
8CMRlOFbCFMM
0;
lOFbCFMM10Rb4NM.Gvk__#.ERR
RRRRRRRRRsbF0
5RRRRRRRRRRRRRRRRRQ:RRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRRmR:kRF0#RR0D8_FOoHRR
RRRRRRRRRRRRRR;R2
8CMRlOFbCFMM
0;
lOFbCFMM10Rb4NM.Gvk__#dERR
RRRRRRRRRsbF0
5RRRRRRRRRRRRRRRRRQ:RRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRRmR:kRF0#RR0D8_FOoHRR
RRRRRRRRRRRRRR;R2
8CMRlOFbCFMM
0;
lOFbCFMM10Rb4NM.Gvk__#cERR
RRRRRRRRRsbF0
5RRRRRRRRRRRRRRRRRQ:RRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRRmR:kRF0#RR0D8_FOoHRR
RRRRRRRRRRRRRR;R2
8CMRlOFbCFMM
0;
lOFbCFMM10Rb4NM.Gvk__#6ERR
RRRRRRRRRsbF0
5RRRRRRRRRRRRRRRRRQ:RRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRRmR:kRF0#RR0D8_FOoHRR
RRRRRRRRRRRRRR;R2
8CMRlOFbCFMM
0;
lOFbCFMM10Rb4NM.Gvk__#nERR
RRRRRRRRRsbF0
5RRRRRRRRRRRRRRRRRQ:RRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRRmR:kRF0#RR0D8_FOoHRR
RRRRRRRRRRRRRR;R2
8CMRlOFbCFMM
0;
lOFbCFMM10Rb4NM.Gvk__#(ERR
RRRRRRRRRsbF0
5RRRRRRRRRRRRRRRRRQ:RRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRRmR:kRF0#RR0D8_FOoHRR
RRRRRRRRRRRRRR;R2
8CMRlOFbCFMM
0;
lOFbCFMM10Rb4NM.Gvk__#UERR
RRRRRRRRRsbF0
5RRRRRRRRRRRRRRRRRQ:RRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRRmR:kRF0#RR0D8_FOoHRR
RRRRRRRRRRRRRR;R2
8CMRlOFbCFMM
0;
lOFbCFMM10Rb4NM.Gvk__#gERR
RRRRRRRRRsbF0
5RRRRRRRRRRRRRRRRRQ:RRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRRmR:kRF0#RR0D8_FOoHRR
RRRRRRRRRRRRRR;R2
8CMRlOFbCFMM
0;
lOFbCFMM10Rb4NM.Gvk_j#4_
ERRRRRRRRRRFRbsR05
RRRRRRRRRRRRRRRRRQR:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRRRmRF:RkR0R#_08DHFoORR
RRRRRRRRRRRRR2RR;M
C8FROlMbFC;M0
F
OlMbFCRM01MbN4k.vG4_#4R_E
RRRRRRRRbRRF5s0RR
RRRRRRRRRRRRRRRRQRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRRmRRRRR:FRk0R8#0_oDFH
ORRRRRRRRRRRRRRRRR2C;
MO8RFFlbM0CM;O

FFlbM0CMRN1bMv4.kPG_RR
RRRRRRRRRb0Fs5RR
RRRRRRRRRRRRRQRRRRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRRm:RRR0FkR0R#8F_DoRHO
RRRRRRRRRRRRRRRR
2;CRM8ObFlFMMC0
;
ObFlFMMC0bR1N.M4v_kG#Pj_RR
RRRRRRRRRb0Fs5RR
RRRRRRRRRRRRRQRRRRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRRm:RRR0FkR0R#8F_DoRHO
RRRRRRRRRRRRRRRR
2;CRM8ObFlFMMC0
;
ObFlFMMC0bR1N.M4v_kG#P4_RR
RRRRRRRRRb0Fs5RR
RRRRRRRRRRRRRQRRRRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRRm:RRR0FkR0R#8F_DoRHO
RRRRRRRRRRRRRRRR
2;CRM8ObFlFMMC0
;
ObFlFMMC0bR1N.M4v_kG#P._RR
RRRRRRRRRb0Fs5RR
RRRRRRRRRRRRRQRRRRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRRm:RRR0FkR0R#8F_DoRHO
RRRRRRRRRRRRRRRR
2;CRM8ObFlFMMC0
;
ObFlFMMC0bR1N.M4v_kG#Pd_RR
RRRRRRRRRb0Fs5RR
RRRRRRRRRRRRRQRRRRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRRm:RRR0FkR0R#8F_DoRHO
RRRRRRRRRRRRRRRR
2;CRM8ObFlFMMC0
;
ObFlFMMC0bR1N.M4v_kG#Pc_RR
RRRRRRRRRb0Fs5RR
RRRRRRRRRRRRRQRRRRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRRm:RRR0FkR0R#8F_DoRHO
RRRRRRRRRRRRRRRR
2;CRM8ObFlFMMC0
;
ObFlFMMC0bR1N.M4v_kG#P6_RR
RRRRRRRRRb0Fs5RR
RRRRRRRRRRRRRQRRRRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRRm:RRR0FkR0R#8F_DoRHO
RRRRRRRRRRRRRRRR
2;CRM8ObFlFMMC0
;
ObFlFMMC0bR1N.M4v_kG#Pn_RR
RRRRRRRRRb0Fs5RR
RRRRRRRRRRRRRQRRRRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRRm:RRR0FkR0R#8F_DoRHO
RRRRRRRRRRRRRRRR
2;CRM8ObFlFMMC0
;
ObFlFMMC0bR1N.M4v_kG#P(_RR
RRRRRRRRRb0Fs5RR
RRRRRRRRRRRRRQRRRRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRRm:RRR0FkR0R#8F_DoRHO
RRRRRRRRRRRRRRRR
2;CRM8ObFlFMMC0
;
ObFlFMMC0bR1N.M4v_kG#PU_RR
RRRRRRRRRb0Fs5RR
RRRRRRRRRRRRRQRRRRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRRm:RRR0FkR0R#8F_DoRHO
RRRRRRRRRRRRRRRR
2;CRM8ObFlFMMC0
;
ObFlFMMC0bR1N.M4v_kG#Pg_RR
RRRRRRRRRb0Fs5RR
RRRRRRRRRRRRRQRRRRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRRm:RRR0FkR0R#8F_DoRHO
RRRRRRRRRRRRRRRR
2;CRM8ObFlFMMC0
;
ObFlFMMC0bR1N.M4v_kG#_4jPRR
RRRRRRRRRsbF0
5RRRRRRRRRRRRRRRRRQ:RRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRRmR:kRF0#RR0D8_FOoHRR
RRRRRRRRRRRRRR;R2
8CMRlOFbCFMM
0;
lOFbCFMM10Rb4NM.Gvk_4#4_
PRRRRRRRRRRFRbsR05
RRRRRRRRRRRRRRRRRQR:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRRRmRF:RkR0R#_08DHFoORR
RRRRRRRRRRRRR2RR;M
C8FROlMbFC;M0
F
OlMbFCRM0#O$M_	OD_NCMLRDC
RRRRRRRRbRRF5s0RR
RRRRRRRRRRRRRRRR7RH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRRhRRBRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRRT:RRR0FkR0R#8F_DoRHO
RRRRRRRRRRRRRRRR
2;CRM8ObFlFMMC0
;
ObFlFMMC0AR1_at.ARkVHo#
CsMCH5ORRS
SXRR:QCM0oRCs;S
SYRR:QCM0oRCs
RSR2R;
RsbF0R5
RmRRRF:Rk#0R0D8_FOoH;R
RRRRQ:MRHR8#0_oDFHRO
R2RR;M
C8FROlMbFC;M0
M
C8
R;




