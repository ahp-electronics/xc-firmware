------------------------------------------------------------------------
@E
---a-RERH#VCHDR#ENRR0FL#CREbHbCC8RM$Osb80C!
!!-a-RERH#VCHDRF#EkRD8MCCPsCRLRH#Eb8bCRRHMs8CNNCLDRsVFl!!!

---a-RERH#P#CsHRFMF0VREvCRq_a])p qRObN	CNoR
H#-1-RbHCOVRHO01FR$DMbHRV$NRM8HM#RFk0R#DNLCFRVsHR#lNkD0MHF
R--B$FbsEHo0OR52gR4gRc,1b$MDHHO0R$,Q3MORDqDRosHER0#sCC#s8PC

---a-RE=CR>bRFC0sNFHsR##RkC08RFbR#CVOH$RRNLDkH0MRHRbHlDCClM00NHRFM
R--VRFsN$R0bFCRskRVMHO0F
M3---
-ERaCsRF8RCsFVVRk0MOH#FMR8NMRO8CDNNs0MHF##RHR0MFRCH8MO0HN0DRFER0C-
-RHFsoNHMDCRPsF#HMFRVsCR#OHks0s$RCFN#M
#3---
-]RfCCN8s/:R/M#$bODHH/0$ObFl.Uj4J4.b/lOFbCHDsP#/E/8DP/E8lEN0_NsCDE3P8Ry4f-
-
R--wRFsw0ksERCs8OC#s0HbHRFM8NC0H,D#RCbDNR#CD	FFRRN0OlFlC#M0RDLCF
I:------------------------------------------------------------------------

---B-RFsb$H0oERg4gn$RLR Q  q3RDsDRH0oE#CRs#PCsC
83---
-ERaH##RFOksCHRVDHCR#MRNR#C#CHM0NbDRNRs0FQVR R  1R084nj(34.-g,gnR Q  0R1NNM8s
8R-e-R]R7pvEN0C0lNHDONROuN	CNo#a3RERH##sFkOVCRHRDClRN$MRF0LOCRFCbH8#,RF,D8RRFs
R--HDMOk88CR0IHEFR#VN0Is0CRERN0H##RFRD8IEH0FRk0I0sH0RCMblCsHH##FVMRsRFl0RECQ   
R--1M0N88Ns#CR7b0Nsl0CM3ERaH##RFOksCHRVDlCRNL$RC#RkC08RFlRHblDCCRM00#EHRN#0Ms8N8-R
-MRN8NRl$CRLR#8H0LsHk80CRRHMObFlH8DCRsVFlMRHR$NMRMlNMRCs#DFRFRMoN0#RE
CR-O-RFHlbDRC8VlFsRC8F#FRM0DRNDRFI8CHsO80RClOFbNHD0MHFRRFV0RECFosHHDMNRk#FsROCVCHD3-
-RHaE#FR#kCsORDVHCNRl$CRLRbOFHRC8VRFsHHM8PkH8NkDR#LCRCC0ICDMRHMOC#RC8ks#C#
3R-a-RERH##sFkOVCRHRDCHb#RsHFP8RC8FNMRM1RqRRQ1LHN##a3REQCR R  8OH#DlNH#hRqY-R
-qRW)h)qa YRX u)1m1R)vRQu pQ7hRQB7pzQRhtqRhYW)q)qYhaRRmwvB )]aqhqpAQQRaY
R--qRh7whQa R11wRm)zR1 wRm)qqRu)BaQz)pqR)uzu m13ERaC#RkCFsRVER0CFR#kCsOR-
-RDVHCER#NRDDHCM8lVMH$MRN8FREDQ8R R  ElNsD#C#RFVslMRN$NR8lCNo#sRFRNDHLHHD0
$R-N-RsHH#MFoRkF0RVER0C#RkCER0CFsCV-3
--
-R0aHDRC:RRRRR0R1NNM8se8R]R7pvEN0C0lNHDONROuN	CNo#QR5 R  1R084nj(34.-g,gnR-
-RRRRRRRRRRRRRqRva)]_ 2qp

---p-RHNLssR$:RRRRa#EHRObN	CNoRN#EDLDRCFROlDbHCH8RMR0FNHRDLssN$-
-RRRRRRRRRRRRR$R#lDLFHDONDM$RN8lCR Q  -3
--
-RP7CCbDFC:s#R RQ 7 RqR1Bep]7R0vNENCl0NHODNRuOo	NCW#RFHs	MtoRsbFk

---u-RkFsb#RC:RRRRa#EHRObN	CNoRV8CH#MCR#NR08NMNRs8VRFs8HC#osMC#FR0RCk#R
HM-R-RRRRRRRRRRRRR8OC#sHHLMeoR]R7plCF8D0#RERN0lCN	RCk#RRFVOlFlF)MR RqpO#FM00NM#-
-RRRRRRRRRRRRRMRN8FROlMlFRq) pDRCCMlC0$NsR0lNENCl0NHODkRVMHO0F3M#

---p-RH0lHNF0HMR:RaRECPkNDCo#RCsMCN80CRRL$0RECVOkM0MHF#MRHRH0E#NRbOo	NCNRl$-
-RRRRRRRRRRRRRNRPsV$RsRFlb0DNVlFsRR0Fb0DNVlFs,MRN8ER0CsRbC#OHHRFMFsVRCD#k0-#
-RRRRRRRRRRRRHRR#MRFDo$RkNNsMC0C8FR0RRLC0REClHHMlRklskCJH8sCRRL$Q   R810R(4jn--
-RRRRRRRRRRRR4RRg3gd

---h-RF#0C:-
-RRRRRRRRRRRRRFRhRO8CDNNs0MHF#sRFRV8CH0MHH#FMRN#EDLDRCMRHO8DkCH8RMF,Rs-
-RRRRRRRRRRRRRGRCO8DkCV8Rs,FlRH0E#NRbOo	NC-3
-RRRRRRRRRRRRaRRE"CRb	NONRoC8DCON0sNH"FMRV8CH#MCRC0ERb0$CR#,#0kL$#bC,MRN8-
-RRRRRRRRRRRRRCR8OsDNNF0HMF#RVqRva)]_ 3qp
R--RRRRRRRRRRRRRCaERN#0Ms8N8NRl0lECNO0HN8DRCMVHHF0HMMRN8FROMMPC0MHFNlDRCHNMM-o
-RRRRRRRRRRRRFRRVER0CNRl0lECNO0HNVDRk0MOH#FMRN0E0sRNCNRbsF0RVER0H##R08NMN
s8-R-RRRRRRRRRRRRRssCbCM#C0ER0CFRVsDlNRl#CNHM0OF#RVER0ClRHblDCCNM00MHFRRFV0
EC-R-RRRRRRRRRRRRRv]qa_q) pNRbOo	NCCR8OsDNNF0HMR3RaRECbbksFR#CF0VREvCRq_a])p q
R--RRRRRRRRRRRRRObN	CNoR8LF$#RHRR0FbPsFHR8CNkRoHD8CHRMCVRFsHDlbCMlC0HN0FRM#0-F
-RRRRRRRRRRRRPRRCVsH$ER0CRHsHDlbCMlC0HN0FFMRVqRva)]_ 3qpRFRaF8DRCDPCFsbC#NRl$-
-RRRRRRRRRRRRREROFCF#RR0FHDlbCMlC0ER0CNRbOo	NCFRL8H$RMER0CFRl#C0RVOVHH0CM
R--RRRRRRRRRRRRRMlNMRCsNHPNDDNLCFR0RC0El-3
--
-R------------------------------------------------------------------------------
-CResF#HMRRRR4:R3-6
-NR70RCRRRRRR.:RckRKD4$Rg
gn---R----------------------------------------------------------------------------
-
-#0$MEHC##MRH0MCsNbD_NNO	obC
NNO	ovCRq_a])p qR
H#RRRRO#FM00NMRbBF$o)HEF0h0CHO:aR1)tQh
RRRR:RR=BR"Fsb$H0oERg4gn RQ R 3qRDDsEHo0s#RCs#CP3C8"
;
RRRR-R-
R-RR-FRBMN#0M70RCMVHHF0HMR#
R-RR-R
RRFROMN#0MR0Rv]qa_m4_e_ ) RR:)p qRR:=jn3d(_U(g4cc44_(c_c.dn.4jR;
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--ekNDCVRFRC4/
RRRRMOF#M0N0vRRq_a] RR:)p qRR:=.43(U_.U4UU.cg_6j_c6.dd6nR;
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--ekNDCVRFRRC
RORRF0M#NRM0Ravq]__.u:QRRq) p=R:R.n3UUd4_j6d((4_gn6U_nc(g
d;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RDeNkFCRV*R.bRH
RORRF0M#NRM0Ravq]Q_uR):R Rqp:d=R344c6.g_n66d_(Ugg.d_dnUc;R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-e-RNCDkRRFVbRH
RORRF0M#NRM0Ravq]Q_u_ me)R_.: R)q:pR=3R46((jgd_n._n(ggcUn4_ng;.d
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-NReDRkCFbVRH
/.RRRRO#FM00NMRqRva4]__ me)Q_uR):R Rqp:j=R3Ud4dgj_U4Un_(Udgnj_(c46;R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-e-RNCDkRRFV4H/b
RRRRMOF#M0N0vRRq_a]umQ_e_ )dRR:)p qRR:=4c3j(_4g(4664n_g6_g((4cn6R;
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--ekNDCVRFR/bHdR
RRFROMN#0MR0Rv]qa__uQm)e _:cRRq) p=R:R(j3Ug6d_nU4dgd_(Ucc_gdjn
.;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RDeNkFCRVHRb/Rc
RORRF0M#NRM0Ravq]__dumQ_e_ ).RR:)p qRR:=c43(._dUUjgUdc_Un_UgUn6(gR;
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--ekNDC*Rdb.H/
RRRRMOF#M0N0vRRq_a]p_mtm.w_R):R Rqp:j=R3dng4(c_46Uj_g6gcd6_j.gc;R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-h-RNs0kNDDRFFoRV
R.RRRRO#FM00NMRqRvap]_mmt_wj_4R):R Rqp:.=R3.dj66U_jgg._jgccn6_U.cj;R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-h-RNs0kNDDRFFoRVjR4
RRRRMOF#M0N0vRRq_a]p.mt__mw RR:)p qRR:=4c3c._ng6jjcUU_Ug_ndccj(;R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-p-RFLoRNR#C.VRFRRC
RORRF0M#NRM0Ravq]m_pt_4jm w_: R)q:pR=3Rjc.dcgc_cU_4gj6d.4._U(;n6
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-FRpoNRL#4CRjVRFRRC
RORRF0M#NRM0Ravq]__4m)e _)1Ta:_.Rq) p=R:R(j3jj(4_Un(4U4_n(6c_c6.c
j;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-Rk#JNRsCs0FFRRFV4
/.RRRRO#FM00NMRqRva1]_T_)a.):R Rqp:4=R3cc4.d4_6dn._j(dgj6_cjUU;R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-#-RJskNCFRsFF0RV
R.RRRRO#FM00NMRqRva7]_ at_mq_)7):R Rqp:j=R3(j4cd6_.6g._g4gc.d_g(6(;R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-FRBMsPC#MHFROVN0RFsVlsFRo8CsRCC0sFRNN8HMR
RRFROMN#0MR0Rv]qa_)1TaQ_u: R)q:pR=3R4(c(.6U_d6_jgj466n._j(;dj
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-JR#kCNsRFsF0VRFR
bHRRRRO#FM00NMRqRva)]_qa7_m _7t):R Rqp:6=R(g3.6_((gd64j._Ud_.jUU(njR;
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-B-RFCMPsF#HMNRVOs0FRFVslNRs8MHNRR0F8sCoC
C
RRRR-R-
R-RR-kRwMHO0F7MRCNODsHN0F
M#RRRR-R-
RVRRk0MOHRFMBp QRR5X:MRHRq) pRR2skC0s)MR ;qp
RRRRRRRRR--ubksF:#C
RRRRRRRRR--RRRRRRRR)kC0sRM##DlND0C#RaQh )t RDPNk5CRN)#R 2qpR0MFR#DC#ER0NXMR
RRRRRRRRR--1ObCHRNDPkNDC
#:RRRRRRRR-R-RRRRRRhRRF
MCRRRRRRRR-7-RFHlNMR:
RRRRR-RR-RRRRRRRRRRXH)MR 
qpRRRRRRRR- -RsssFRMOF8HH0F:M#
RRRRRRRRR--RRRRRRRRhCFM
RRRRRRRRR--)oNMCR:
RRRRR-RR-RRRRRRRR RBQXp52#RHR0lNENCl0NHODRD$kFMLkCM88R
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRRNRR2lRQblDCCNM00MHF#NREP0CRFkR#bsbF00RNRNDC#00RE8CRFHlNMR
RRRRRR-R-RRRRRRRRRRRRRRRRq5A1X<2RRq) ph5Qa  t)Q']t
]2
RRRRMVkOF0HMQR1t5hRXH:RM R)q2pRR0sCkRsM)p q;R
RRRRRR-R-RsukbCF#:R
RRRRRR-R-RRRRRRRRR0)Ck#sMRj43RRHVXRR>j;3jRjj3RRHVXRR=j;3jR3-4jVRHR<XRRjj3
RRRRRRRRR--1ObCHRNDPkNDC
#:RRRRRRRR-R-RRRRRRhRRF
MCRRRRRRRR-7-RFHlNMR:
RRRRR-RR-RRRRRRRRRRXH)MR 
qpRRRRRRRR- -RsssFRMOF8HH0F:M#
RRRRRRRRR--RRRRRRRRhCFM
RRRRRRRRR--)oNMCR:
RRRRR-RR-RRRRRRRRARq1Q51tXh52<2R=3R4jR
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRRhRRF
MC
RRRRMVkOF0HMmR)zRh75:XRRRHM)p qRs2RCs0kM R)q
p;RRRRRRRR-u-RkFsb#
C:RRRRRRRR-R-RRRRRR)RRF8kM#RRX00FREMCRCCNs#H0RMo0CCPsRNCDkR#5NRNsCDR23QXVRR
H#RRRRRRRR-R-RRRRRRERRNIDVNL$RCC0IC0MRIHFRMo0CC,s#RksFMM8Ho#RHRNNI$sRVFjlR3Rj
RRRRR-RR-bR1CNOHDNRPD#kC:R
RRRRRR-R-RRRRRRRRRz)mhj753Rj2=3RjjR
RRRRRR-R-Rl7FN:HM
RRRRRRRRR--RRRRRRRRXMRHRq) pR
RRRRRR-R-Rs sFOsRFHM80MHF#R:
RRRRR-RR-RRRRRRRRFRhMRC
RRRRR-RR-NR)M:oC
RRRRRRRRR--RRRRRRRR)hmz725XRRH#lEN0C0lNHDONDk$RMkLFM88C
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRR2RNRbQlDCClM00NH#FMRPENCFR0Rb#kb0FsRRN0D#CN0ER0CFR8lMNH
RRRRRRRRR--RRRRRRRRRRRRRqRRAX152RR<)p q5aQh )t 't]Q]
2
RRRRVOkM0MHFRq) phvQR,5XR:YRRRHM)p qRs2RCs0kM R)q
p;RRRRRRRR-u-RkFsb#
C:RRRRRRRR-R-RRRRRR)RRCs0kM0#RENCRDLoCsONHN$DDRN#lDsDCRRFVXMRN8
RYRRRRRRRR-1-RbHCONPDRNCDk#R:
RRRRR-RR-RRRRRRRR R)qQpvh,5XY=2RRIXRERCMXRR=YR
RRRRRR-R-Rl7FN:HM
RRRRRRRRR--RRRRRRRRXMRHRq) pY;RRRHM)p q
RRRRRRRRR-- FsssFROM08HH#FM:R
RRRRRR-R-RRRRRRRRRMhFCR
RRRRRR-R-RM)No
C:RRRRRRRR-R-RRRRRR)RR vqpQXh5,RY2Hl#RNC0ElHN0ODND$MRkLMFk8
C8RRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRRMhFCR

RVRRk0MOHRFMah)zBXR5RH:RM R)q2pRR0sCkRsM)p q;R
RRRRRR-R-RsukbCF#:R
RRRRRR-R-RRRRRRRRRkasM0ONCX#RRI0FN#s8Rjj3R8NMR0sCk#sMRk0sM0ONCP8RNCDk
RRRRRRRRR--1ObCHRNDPkNDC
#:RRRRRRRR-R-RRRRRRaRR)Bzh5jj32RR=j
3jRRRRRRRR-7-RFHlNMR:
RRRRR-RR-RRRRRRRRRRXH)MR 
qpRRRRRRRR- -RsssFRMOF8HH0F:M#
RRRRRRRRR--RRRRRRRRhCFM
RRRRRRRRR--)oNMCR:
RRRRR-RR-RRRRRRRR)Raz5hBXH2R#NRl0lECNO0HN$DDRLkMF8kMCR8
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRRRRNQ2RlCbDl0CMNF0HME#RNRPC0#FRkFbbsN0R0CRDNR#00REC8NFlHRM
RRRRR-RR-RRRRRRRRRRRRRRRR1qA5RX2< R)qQp5hta  ])'Q2t]
R
RRkRVMHO0FwMRp)mmRR5X:MRHRq) pRR2skC0s)MR ;qp
RRRRRRRRR--ubksF:#C
RRRRRRRRR--RRRRRRRR)kC0sRM#DoNsCR#0Q hatR )PkNDCNR5# R)qRp2MRF0oNsC0RCs0MENRRX
RRRRR-RR-bR1CNOHDNRPD#kC:R
RRRRRR-R-RRRRRRRRRmwpmj)53Rj2=3RjjR
RRRRRR-R-Rl7FN:HM
RRRRRRRRR--RRRRRRRRXMRHRq) pR
RRRRRR-R-Rs sFOsRFHM80MHF#R:
RRRRR-RR-RRRRRRRRFRhMRC
RRRRR-RR-NR)M:oC
RRRRRRRRR--RRRRRRRRwmpm)25XRRH#lEN0C0lNHDONDk$RMkLFM88C
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRR2RNRbQlDCClM00NH#FMRPENCFR0Rb#kb0FsRRN0D#CN0ER0CFR8lMNH
RRRRRRRRR--RRRRRRRRRRRRRqRRAX152RR<)p q5aQh )t 't]Q]
2
RRRRVOkM0MHFRm"v75"RXY,R:MRHRq) pRR2skC0s)MR ;qp
RRRRRRRRR--ubksF:#C
RRRRRRRRR--RRRRRRRR)kC0sRM#VNDF0oHMRHbFMl0RFD8kkF#RV/RXYI,RHR0E0REC#CNlRo#HM#RN
RRRRRRRRR--RRRRRRRRYN,RMN8RLD#FkR0CPkNDCCRD#0#RERNM0RECNFL#DCk0RDPNkFCRV,RYR8NM
RRRRRRRRR--RRRRRRRRVRFs#CFlRaQh )t RDPNkhCRRC0ER#sCkRD0#HN0#CVH#ER0CCRsDHN0FRM
RRRRR-RR-RRRRRRRRRRX=*RYhRR+v5m7X2,Y
RRRRRRRRR--1ObCHRNDPkNDC
#:RRRRRRRR-R-RRRRRRhRRF
MCRRRRRRRR-7-RFHlNMR:
RRRRR-RR-RRRRRRRRRRXH)MR ;qpRHYRM R)qNpRMY8RRR/=j
3jRRRRRRRR- -RsssFRMOF8HH0F:M#
RRRRRRRRR--RRRRRRRR FsssVRHR=YRRjj3
RRRRRRRRR--)oNMCR:
RRRRR-RR-RRRRRRRRARq1m5v7,5XYR22<ARq125Y
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRRFRhM
C
RRRRVOkM0MHFRq) pXvqR,5XR:YRRRHM)p qRs2RCs0kM R)q
p;RRRRRRRR-u-RkFsb#
C:RRRRRRRR-R-RRRRRR)RRCs0kM0#RENCRDLoCsONHN$DDRsDNoRCsFXVRR8NMRRY
RRRRR-RR-bR1CNOHDNRPD#kC:R
RRRRRR-R-RRRRRRRRRq) pXvq5YX,2RR=XERICXMRRY=R
RRRRRRRRR--7NFlH
M:RRRRRRRR-R-RRRRRRXRRRRHM)p q;RRYH)MR 
qpRRRRRRRR- -RsssFRMOF8HH0F:M#
RRRRRRRRR--RRRRRRRRhCFM
RRRRRRRRR--)oNMCR:
RRRRR-RR-RRRRRRRR R)qqpvX,5XYH2R#NRl0lECNO0HN$DDRLkMF8kMCR8
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRRRRhCFM
R
RRkRVMHO0F1MRTR)a5:XRRRHM)p qRs2RCs0kM R)q
p;RRRRRRRR-u-RkFsb#
C:RRRRRRRR-R-RRRRRR)RRCs0kM##RJskNCFRsFF0RV
RXRRRRRRRR-1-RbHCONPDRNCDk#R:
RRRRR-RR-RRRRRRRRTR1)ja53Rj2=3RjjR
RRRRRR-R-RRRRRRRRR)1Ta354j=2RRj43
RRRRRRRRR--7NFlH
M:RRRRRRRR-R-RRRRRRXRRRR>=j
3jRRRRRRRR- -RsssFRMOF8HH0F:M#
RRRRRRRRR--RRRRRRRR FsssVRHR<XRRjj3
RRRRRRRRR--)oNMCR:
RRRRR-RR-RRRRRRRRTR1)Xa52=R>Rjj3
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRR2RNRCaERbkbCLsRF8kMRRFV0RECsOCNEDNLCNRsMRoCF1VRTR)aHR#
RRRRR-RR-RRRRRRRRRRRRbNbsHFGlCN0Do$RHMPCR:L$
RRRRRRRRR--RRRRRRRRRRRRR1RRT5)aX<2R=TR1))a5 'qp]]Qt2R

RbRRsCFO8CksRQzhwvm)5sPNHDNLC R1 ,7417  .M:HFRk0uQm1a Qe;NRPsLHNDXCR:0FkRq) p
2;RRRRRRRR-u-RkFsb#
C:RRRRRRRR-R-RRRRRR)RRCs0kMR#,HXMR,RRNbk#C8sF-NFM8lkRMlsLCR0IHEMRkHsVFlR
RRRRRR-R-RRRRRRRRR#8H0LsHkF0HMMRHRC0ERCFbMMRH0PCsN5DRj,3jRj432R3
RRRRR-RR-bR1CNOHDNRPD#kC:R
RRRRRR-R-RRRRRRRRRMhFCR
RRRRRR-R-Rl7FN:HM
RRRRRRRRR--RRRRRRRR4=R<R 1 7<4R=4R.cU(cd.6n;RR4<1=R . 7RR<=.(4ccdUdgRU
RRRRR-RR-sR sRFsO8FMHF0HM
#:RRRRRRRR-R-RRRRRR RRsssFRRHV17  4sRFR 1 7F.RkH0#8FCRVNRPDRH88NFlHRM
RRRRR-RR-NR)M:oC
RRRRRRRRR--RRRRRRRRjR3j<RRX<3R4jR
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRRNRR2ERaCCR#l0NMHRO#VRFs0#EHRMVkOF0HMsRNCCR8#HOsLRC8L0$RERC
RRRRR-RR-RRRRRRRRRRRRoNDF0sHEblRkHLD#8ECRRL$usHCspCR'k O$RCsH"MRBlFlkOMHNF0HMR#
RRRRR-RR-RRRRRRRRRRRRRFV0RECq,Bv"FRPDd3R4M,RFn3R,kRKM4CRg,UUR3bbR.(c-c((3R
RRRRRR-R-RRRRRRRRRRRRaRECNFDosEH0l#RHR#LNCF8RMER0CFROlMLHNF0HMVRFRF0I
RRRRRRRRR--RRRRRRRRRlRRkHD0bODHNP0HCHRDMsCNRMOFoCskMN0HDCRoMNCs0#FsRsVFR-d.L
H0RRRRRRRR-R-RRRRRRRRRRDRbNF0Vs3l#
RRRRRRRR
--RRRRRRRR-R-RRRRRRLRR2CRAVCFsRC0ERsVH#O0RNRDD0zFRhmQw)Rv,0REC#8CCRDPNk
C#RRRRRRRR-R-RRRRRRRRRR1R5 4 7, R1 27.RPENCFR0RRLCH0MHHHNDxRC80PFRNCDk#MRHRC0ERMsNoRC
RRRRR-RR-RRRRRRRRRRRR,r4Rc.4(dcU69n.R8NMR,r4Rc.4(dcUd9gUR#sCb0COHDPC$R3Ra
ECRRRRRRRR-R-RRRRRRRRRRCR#CP8RNCDk#sRNCFRl8HHVCN8RVs0CROCNENROD0DRFhRzQ)wmvR3
RRRRR-RR-R
RRRRRR-R-RRRRRRRRRRO2a#EHRMsN8RFlMLklCosRCsMCNs0FRRH#b0FsNCLDRsVFR-d.L
H0RRRRRRRR-R-RRRRRRRRRRFROl0bkC,s#R8NMRRH0ERN#NCRbs8HFRRFV~d.3jc6U*j54*U*42FRVsNRCORE
RRRRR-RR-RRRRRRRRRRRR0#CRRFV#8CCRDPNk3C#
RRRRRRRR
--RRRRRRRR-R-RRRRRR8RR2FRwsMRHVlFsNF0HMMRFRC#bON0sDCR0#R0#VRFs0RECNFDosEH0ls,RCsVC
RRRRRRRRR--RRRRRRRRR0RRFER0C'Rp $OkCNsRsO0HD
C3
RRRRMVkOF0HMARB)5aRXRR:H)MR Rqp2CRs0MksRq) pR;
RRRRR-RR-kRus#bFCR:
RRRRR-RR-RRRRRRRRCR)0Mks#kROLsCRFRF0FXVR
RRRRRRRRR--1ObCHRNDPkNDC
#:RRRRRRRR-R-RRRRRRBRRA5)aj23jRj=R3Rj
RRRRR-RR-RRRRRRRRARB)4a53Rj2=3R4jR
RRRRRR-R-RRRRRRRRR)BAa45-3Rj2=4R-3Rj
RRRRR-RR-FR7lMNH:R
RRRRRR-R-RRRRRRRRRHXRM R)qRp
RRRRR-RR-sR sRFsO8FMHF0HM
#:RRRRRRRR-R-RRRRRRhRRF
MCRRRRRRRR-)-RNCMo:R
RRRRRR-R-RRRRRRRRR)BAa25XRRH#lEN0C0lNHDONDk$RMkLFM88C
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRR2RNRCaERNsCOLENDsCRNCMoRRFVBaA)RRH#NsbbFlGHND0C$HRoPRCML
$:RRRRRRRR-R-RRRRRRRRRRRRRRARq1A5B)Xa52<2R=ARB))a5 'qp]]Qt2R

RVRRk0MOHRFM""**RR5X:MRHRaQh )t ;RRY:MRHRq) ps2RCs0kM R)q
p;RRRRRRRR-u-RkFsb#
C:RRRRRRRR-R-RRRRRR)RRCs0kMY#RRIbFCFsRVRRX=R=>R*X*YR
RRRRRR-R-RC1bODHNRDPNk:C#
RRRRRRRRR--RRRRRRRRXj**3=jRRj43;RRX/j=R
RRRRRRRRR--RRRRRRRRjY**Rj=R3Rj;YRR>j
3jRRRRRRRR-R-RRRRRRXRR*3*4jRR=)p q5;X2R>XR=
RjRRRRRRRR-R-RRRRRR4RR*R*Y=3R4jR
RRRRRR-R-Rl7FN:HM
RRRRRRRRR--RRRRRRRRXRR>jR
RRRRRR-R-RRRRRRRRR=XRRVjRFYsRRj>R3Rj
RRRRR-RR-RRRRRRRRRRX<RRjVRFsYRR=j
3jRRRRRRRR- -RsssFRMOF8HH0F:M#
RRRRRRRRR--RRRRRRRR FsssVRHR<XRRNjRMY8RRR/=j
3jRRRRRRRR-R-RRRRRR RRsssFRRHVXRR=jMRN8RRY<j=R3Rj
RRRRR-RR-NR)M:oC
RRRRRRRRR--RRRRRRRRXY**RR>=j
3jRRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRRRN2aRECkCbbsFRLkRM8F0VREsCRCENONCLDRMsNoVCRF"sR*R*"HR#
RRRRR-RR-RRRRRRRRRRRRbNbsHFGlCN0Do$RHMPCR:L$
RRRRRRRRR--RRRRRRRRRRRRRXRR*R*Y<)=R 'qp]]Qt
R
RRkRVMHO0F"MR*R*"5:XRRRHM)p q;RRY:MRHRq) ps2RCs0kM R)q
p;RRRRRRRR-u-RkFsb#
C:RRRRRRRR-R-RRRRRR)RRCs0kMY#RRIbFCFsRVRRX=R=>R*X*YR
RRRRRR-R-RC1bODHNRDPNk:C#
RRRRRRRRR--RRRRRRRRXj**3=jRRj43;RRX/j=R3Rj
RRRRR-RR-RRRRRRRR3RjjY**Rj=R3Rj;YRR>j
3jRRRRRRRR-R-RRRRRRXRR*3*4jRR=XX;RRR>=j
3jRRRRRRRR-R-RRRRRR4RR3*j*YRR=4
3jRRRRRRRR-7-RFHlNMR:
RRRRR-RR-RRRRRRRRRRX>3RjjR
RRRRRR-R-RRRRRRRRR=XRRjj3RsVFR>YRRjj3
RRRRRRRRR--RRRRRRRRXRR<jR3jVRFsYRR=j
3jRRRRRRRR- -RsssFRMOF8HH0F:M#
RRRRRRRRR--RRRRRRRR FsssVRHR<XRRjj3R8NMR/YR=3RjjR
RRRRRR-R-RRRRRRRRRs sFHsRVRRX=3RjjMRN8RRY<j=R3Rj
RRRRR-RR-NR)M:oC
RRRRRRRRR--RRRRRRRRXY**RR>=j
3jRRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRRRN2aRECkCbbsFRLkRM8F0VREsCRCENONCLDRMsNoVCRF"sR*R*"HR#
RRRRR-RR-RRRRRRRRRRRRbNbsHFGlCN0Do$RHMPCR:L$
RRRRRRRRR--RRRRRRRRRRRRRXRR*R*Y<)=R 'qp]]Qt
R
RRkRVMHO0FpMRm5tRXRR:H)MR Rqp2CRs0MksRq) p>R=Rs"l_oDF"R;
RRRRR-RR-kRus#bFCR:
RRRRR-RR-RRRRRRRRCR)0Mks#NRM0NksDFRDoHNs0RElFXVR
RRRRRRRRR--1ObCHRNDPkNDC
#:RRRRRRRR-R-RRRRRRpRRm4t53Rj2=3RjjR
RRRRRR-R-RRRRRRRRRtpm5avq]2_ R4=R3Rj
RRRRR-RR-FR7lMNH:R
RRRRRR-R-RRRRRRRRR>XRRjj3
RRRRRRRRR-- FsssFROM08HH#FM:R
RRRRRR-R-RRRRRRRRRs sFHsRVRRX<j=R3Rj
RRRRR-RR-NR)M:oC
RRRRRRRRR--RRRRRRRRp5mtXH2R#NRl0lECNO0HN$DDRLkMF8kMCR8
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRRRRNa2REsCRCENONCLDRMsNoFCRVmRpt#RHRbNbsHFGlCN0Do$RHMPCR:L$
RRRRRRRRR--RRRRRRRRRRRRRpRRmjt5+<2R=mRpt25XRR<=p5mt)p q't]Q]
2
RRRRVOkM0MHFRu XRR5X:MRHRq) pRR2skC0s)MR Rqp=">RlCs_G;b"
RRRRRRRRR--ubksF:#C
RRRRRRRRR--RRRRRRRR)kC0sRM#CX**;ERICRsCCRR=v]qa_R 
RRRRR-RR-bR1CNOHDNRPD#kC:R
RRRRRR-R-RRRRRRRRRu X5jj32RR=4
3jRRRRRRRR-R-RRRRRR RRX4u53Rj2=qRva ]_
RRRRRRRRR--RRRRRRRR 5Xu-j432RR=v]qa_m4_e_ ) R
RRRRRR-R-RRRRRRRRRu X5RX2=3RjjFRVsRRX<-=Rp5mt)p q't]Q]R2
RRRRR-RR-FR7lMNH:R
RRRRRR-R-RRRRRRRRRHXRM R)q#pRkROE00ENRu X5RX2<)=R 'qp]]Qt
RRRRRRRRR-- FsssFROM08HH#FM:R
RRRRRR-R-RRRRRRRRRs sFHsRVRRX>mRpt 5)q]p'Q2t]
RRRRRRRRR--)oNMCR:
RRRRR-RR-RRRRRRRRXR u25XRR>=j
3jRRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRRRN2aRECkL#ND8CRFHlNMVRFRu XRRH#NsbbFlGHND0C$HRoPRCML
$:RRRRRRRR-R-RRRRRRRRRRRRRRRRX<p=Rm)t5 'qp]]Qt2R

RVRRk0MOHRFMp.mtRR5X:MRHRq) pRR2skC0s)MR ;qp
RRRRRRRRR--ubksF:#C
RRRRRRRRR--RRRRRRRR)kC0sRM#DNFosEH0lNRL#.CRRRFVXR
RRRRRR-R-RC1bODHNRDPNk:C#
RRRRRRRRR--RRRRRRRRp.mt5j432RR=j
3jRRRRRRRR-R-RRRRRRpRRm5t..23jR4=R3Rj
RRRRR-RR-FR7lMNH:R
RRRRRR-R-RRRRRRRRR>XRRjj3
RRRRRRRRR-- FsssFROM08HH#FM:R
RRRRRR-R-RRRRRRRRRs sFHsRVRRX<j=R3Rj
RRRRR-RR-NR)M:oC
RRRRRRRRR--RRRRRRRRp.mt5RX2Hl#RNC0ElHN0ODND$MRkLMFk8
C8RRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRRRN2aRECsOCNEDNLCNRsMRoCFpVRmRt.HN#RbFbsGNHl0$CDRPoHCLMR$R:
RRRRR-RR-RRRRRRRRRRRRRRRRtpm.+5j2=R<Rtpm.25XRR<=p.mt5q) pQ']t
]2
RRRRMVkOF0HMmRptXR5:MRHRq) pA;Rq:1 RRHM)p q2CRs0MksRq) pR;
RRRRR-RR-kRus#bFCR:
RRRRR-RR-RRRRRRRRCR)0Mks#FRDoHNs0RElLCN#R1Aq VRFRRX
RRRRR-RR-bR1CNOHDNRPD#kC:R
RRRRRR-R-RRRRRRRRRtpm5j43,qRA1R 2=3RjjR
RRRRRR-R-RRRRRRRRRtpm51Aq A,Rq21 R4=R3Rj
RRRRR-RR-FR7lMNH:R
RRRRRR-R-RRRRRRRRR>XRRjj3
RRRRRRRRR--RRRRRRRRA q1Rj>R3Rj
RRRRR-RR-RRRRRRRRqRA1/ R=3R4jR
RRRRRR-R-Rs sFOsRFHM80MHF#R:
RRRRR-RR-RRRRRRRRsR sRFsHXVRRR<=j
3jRRRRRRRR-R-RRRRRR RRsssFRRHVA q1RR<=j
3jRRRRRRRR-R-RRRRRR RRsssFRRHVA q1R4=R3Rj
RRRRR-RR-NR)M:oC
RRRRRRRRR--RRRRRRRRp5mtXA,Rq21 RRH#lEN0C0lNHDONDk$RMkLFM88C
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRR2RNRCWEMqRA1> RRj43,ER0CCRsNNOELRDCsoNMCVRFRtpmR
H#RRRRRRRR-R-RRRRRRRRRRbRNbGsFH0lNCRD$oCHPM$RL:R
RRRRRR-R-RRRRRRRRRRRRRRRRp5mtjR+,A q12=R<Rtpm5RX,A q12=R<Rtpm5q) pQ']tR],A q12R
RRRRRR-R-RRRRRRRRRRL2WMECRjj3RA<RqR1 <3R4j0,REsCRCENONCLDRMsNoFCRVmRpt#RH
RRRRRRRRR--RRRRRRRRRNRRbFbsGNHl0$CDRPoHCLMR$R:
RRRRR-RR-RRRRRRRRRRRRRRRRtpm5q) pQ']tR],A q12=R<Rtpm5RX,A q12=R<Rtpm5,j+R1Aq 
2
RRRRVOkM0MHFRtpm45jRXRR:H)MR Rqp2CRs0MksRq) pR;
RRRRR-RR-kRus#bFCR:
RRRRR-RR-RRRRRRRRCR)0Mks#FRDoHNs0RElLCN#RR4jFXVR
RRRRRRRRR--1ObCHRNDPkNDC
#:RRRRRRRR-R-RRRRRRpRRmjt45j432RR=j
3jRRRRRRRR-R-RRRRRRpRRmjt4534jj=2RRj43
RRRRRRRRR--7NFlH
M:RRRRRRRR-R-RRRRRRXRRRj>R3Rj
RRRRR-RR-sR sRFsO8FMHF0HM
#:RRRRRRRR-R-RRRRRR RRsssFRRHVX=R<Rjj3
RRRRRRRRR--)oNMCR:
RRRRR-RR-RRRRRRRRmRpt54jXH2R#NRl0lECNO0HN$DDRLkMF8kMCR8
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRRRRNa2REsCRCENONCLDRMsNoFCRVmRptR4jHN#RbFbsGNHl0$CDRPoHCLMR$R:
RRRRR-RR-RRRRRRRRRRRRRRRRtpm4jj5+<2R=mRpt54jX<2R=mRpt54j)p q't]Q]
2
RRRRVOkM0MHFRQR1hXR5RH:RM R)q2pRR0sCkRsM)p qRR=>"_ls#"HM;R
RRRRRR-R-RsukbCF#:R
RRRRRR-R-RRRRRRRRR0)Ck#sMRM#HCVRFRRX;XMRHR8sNH#NM
RRRRRRRRR--1ObCHRNDPkNDC
#:RRRRRRRR-R-RRRRRR1RRQXh52RR=jR3jVRFsXRR=	q*vau]_QI,RECCsRH	R#MRNRaQh )t 
RRRRRRRRR--RRRRRRRR15QhX=2RRj43RsVFR=XRR*5c	2+4*avq]Q_u_ me),_.RCIEs	CRRRH#NRM
RRRRR-RR-RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRQ hat
 )RRRRRRRR-R-RRRRRR1RRQXh52RR=-j43RsVFR=XRR*5c	2+d*avq]Q_u_ me),_.RCIEs	CRRRH#NRM
RRRRR-RR-RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRQ hat
 )RRRRRRRR-7-RFHlNMR:
RRRRR-RR-RRRRRRRRRRXH)MR 
qpRRRRRRRR- -RsssFRMOF8HH0F:M#
RRRRRRRRR--RRRRRRRRhCFM
RRRRRRRRR--)oNMCR:
RRRRR-RR-RRRRRRRRARq1Q51h25X2=R<Rj43
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRR2RNRswFRsDNoRCsPkNDCF#RVARq125X,CR8o8sNCN8ROsOkNRO$HN#RDIDFC
83
RRRRMVkOF0HMBRRm51RR:XRRRHM)p qRs2RCs0kM R)q=pR>lR"sF_O#
";RRRRRRRR-u-RkFsb#
C:RRRRRRRR-R-RRRRRR)RRCs0kMO#RFM#HCVRFRRX;XMRHR8sNH#NM
RRRRRRRRR--1ObCHRNDPkNDC
#:RRRRRRRR-R-RRRRRRBRRmX152RR=jR3jVRFsXRR=5	.*+*42v]qa__uQm)e _R.,IsECCRR	HN#RMR
RRRRRR-R-RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRQ hat
 )RRRRRRRR-R-RRRRRRBRRmX152RR=4R3jVRFsXRR=5	.*2q*vau]_QI,RECCsRH	R#MRNRaQh )t 
RRRRRRRRR--RRRRRRRRB5m1X=2RR3-4jFRVsRRX=.R5*4	+2q*vau]_QI,RECCsRH	R#MRNRaQh )t 
RRRRRRRRR--7NFlH
M:RRRRRRRR-R-RRRRRRXRRRRHM)p q
RRRRRRRRR-- FsssFROM08HH#FM:R
RRRRRR-R-RRRRRRRRRMhFCR
RRRRRR-R-RM)No
C:RRRRRRRR-R-RRRRRRqRRAB15mX152<2R=3R4jR
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRRNRR2FRwsNRDssoCRDPNkRC#FqVRAX1528,RCNos8RC8NkOOs$NORRH#NFDDI3C8
R
RRkRVMHO0FRMRaRqh5:XRRRHM)p qRs2RCs0kM R)q
p;RRRRRRRR-u-RkFsb#
C:RRRRRRRR-R-RRRRRR)RRCs0kM0#RNCMoMF0RV;RXRHXRMNRs8MHN#R
RRRRRR-R-RC1bODHNRDPNk:C#
RRRRRRRRR--RRRRRRRRa5qhX=2RRjj3RsVFR=XRRv	*q_a]uRQ,IsECCRR	HN#RMhRQa  t)R
RRRRRR-R-Rl7FN:HM
RRRRRRRRR--RRRRRRRRXMRHRq) pMRN8R
RRRRRR-R-RRRRRRRRR/XR=.R5*4	+2q*vau]_Qe_m .)_,ERICRsC	#RHRRNMQ hat
 )RRRRRRRR- -RsssFRMOF8HH0F:M#
RRRRRRRRR--RRRRRRRR FsssVRHR=XRR.55*4	+2RR*v]qa__uQm)e _,.2RCIEs	CRRRH#NRM
RRRRR-RR-RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRQ hat
 )RRRRRRRR-)-RNCMo:R
RRRRRR-R-RRRRRRRRRhaq5RX2Hl#RNC0ElHN0ODND$MRkLMFk8
C8RRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRRRN2wRFsDoNsCPsRNCDk#VRFR1qA5,X2Ro8CsCN88ORNONksOH$R#DRNDCFI8
3
RRRRVOkM0MHFR)RqBh1QRR5X:MRHRq) pRR2skC0s)MR ;qp
RRRRRRRRR--ubksF:#C
RRRRRRRRR--RRRRRRRR)kC0sRM#HCMPsR#C#CHMRRFVXR
RRRRRR-R-RC1bODHNRDPNk:C#
RRRRRRRRR--RRRRRRRRq1)BQjh53Rj2=3RjjR
RRRRRR-R-RRRRRRRRRBq)15Qh423jRv=Rq_a]umQ_e_ ).R
RRRRRR-R-RRRRRRRRRBq)15Qh-j432RR=-avq]Q_u_ me)
_.RRRRRRRR-7-RFHlNMR:
RRRRR-RR-RRRRRRRRARq125XRR<=4
3jRRRRRRRR- -RsssFRMOF8HH0F:M#
RRRRRRRRR--RRRRRRRR FsssVRHR1qA5RX2>3R4jR
RRRRRR-R-RM)No
C:RRRRRRRR-R-RRRRRRqRRAq15)QB1h25XRR<=v]qa__uQm)e _R.
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRRRRhCFM
R
RRkRVMHO0FRMRqB)Bm51RXRR:H)MR Rqp2CRs0MksRq) pR;
RRRRR-RR-kRus#bFCR:
RRRRR-RR-RRRRRRRRCR)0Mks#MRHP#CsCFRO#CHMRRFVXR
RRRRRR-R-RC1bODHNRDPNk:C#
RRRRRRRRR--RRRRRRRRqB)Bm4153Rj2=3RjjR
RRRRRR-R-RRRRRRRRRBq)B5m1j23jRv=Rq_a]umQ_e_ ).R
RRRRRR-R-RRRRRRRRRBq)B5m1-j432RR=v]qa_
uQRRRRRRRR-7-RFHlNMR:
RRRRR-RR-RRRRRRRRARq125XRR<=4
3jRRRRRRRR- -RsssFRMOF8HH0F:M#
RRRRRRRRR--RRRRRRRR FsssVRHR1qA5RX2>3R4jR
RRRRRR-R-RM)No
C:RRRRRRRR-R-RRRRRRjRR3<jR=)RqB1Bm5RX2<v=Rq_a]uRQ
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRRRRhCFM
R
RRkRVMHO0FRMRqa)Bq5hRYRR:H)MR 2qpR0sCkRsM)p q;R
RRRRRR-R-RsukbCF#:R
RRRRRR-R-RRRRRRRRR0)Ck#sMRC0ERDPNkFCRVER0CMRNoRDCHsMRNN8HMF#RVER0CFRbH
M0RRRRRRRR-R-RRRRRR4R53Rj,YR2,IOEHE#RHRRHMs0CONkMoDRNsOsFF8NHM0
C#RRRRRRRR-1-RbHCONPDRNCDk#R:
RRRRR-RR-RRRRRRRR)RqBhaq5jj32RR=j
3jRRRRRRRR-7-RFHlNMR:
RRRRR-RR-RRRRRRRRRRYH)MR 
qpRRRRRRRR- -RsssFRMOF8HH0F:M#
RRRRRRRRR--RRRRRRRRhCFM
RRRRRRRRR--)oNMCR:
RRRRR-RR-RRRRRRRRARq1)5qBhaq52Y2RR<=v]qa__uQm)e _R.
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRRRRhCFM
R
RRkRVMHO0FRMRqa)Bq5hRYRR:H)MR ;qpR:XRRRHM)p q2CRs0MksRq) pR;
RRRRR-RR-kRus#bFCR:
RRRRR-RR-RRRRRRRRCR)0Mks#ER0CsRbHHMObRNDPkNDCVRFRC0ERoNMDHCRMNRs8MHN#VRF
RRRRRRRRR--RRRRRRRR0RECbMFH0XR5,2RY,ERIHROEHH#RMCRsOM0NoNkDsFROFHs8MCN0#R
RRRRRR-R-RC1bODHNRDPNk:C#
RRRRRRRRR--RRRRRRRRqa)Bqjh53Rj,X=2RRjj3RRHVXRR>j
3jRRRRRRRR-R-RRRRRRqRR)qBah35jjX,R2RR=v]qa_RuQHXVRRj<R3Rj
RRRRR-RR-RRRRRRRR)RqBhaq5RY,j23jRv=Rq_a]umQ_e_ ).VRHR>YRRjj3
RRRRRRRRR--RRRRRRRRqa)BqYh5,3Rjj=2RRq-vau]_Qe_m .)_RRHVYRR<j
3jRRRRRRRR-7-RFHlNMR:
RRRRR-RR-RRRRRRRRRRYH)MR 
qpRRRRRRRR-R-RRRRRRXRRRRHM)p q,RRX/j=R3IjRERCMYRR=j
3jRRRRRRRR- -RsssFRMOF8HH0F:M#
RRRRRRRRR--RRRRRRRR FsssVRHR=XRRjj3R8NMR=YRRjj3
RRRRRRRRR--)oNMCR:
RRRRR-RR-RRRRRRRRvR-q_a]u<QRRBq)a5qhY2,XRR<=v]qa_
uQRRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRRMhFCR

RVRRk0MOHRFM1]QhRR5X:MRHRq) ps2RCs0kM R)q
p;RRRRRRRR-u-RkFsb#
C:RRRRRRRR-R-RRRRRR)RRCs0kME#R$sbCLHFDOHR#MFCRV
RXRRRRRRRR-1-RbHCONPDRNCDk#R:
RRRRR-RR-RRRRRRRRQR1hj]53Rj2=3RjjR
RRRRRR-R-Rl7FN:HM
RRRRRRRRR--RRRRRRRRXMRHRq) pR
RRRRRR-R-Rs sFOsRFHM80MHF#R:
RRRRR-RR-RRRRRRRRFRhMRC
RRRRR-RR-NR)M:oC
RRRRRRRRR--RRRRRRRR1]Qh5RX2Hl#RNC0ElHN0ODND$MRkLMFk8
C8RRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRRRN2aRECkL#ND8CRFHlNMVRFRh1Q]#RHRbNbsHFGlCN0Do$RHMPCR:L$
RRRRRRRRR--RRRRRRRRRRRRRqRRAX152=R<Rtpm5q) pQ']t
]2
R
RRkRVMHO0FBMRmR1]5:XRRRHM)p q2CRs0MksRq) pR;
RRRRR-RR-kRus#bFCR:
RRRRR-RR-RRRRRRRRCR)0Mks#$REbLCsFODHR#OFHRMCFXVR
RRRRRRRRR--1ObCHRNDPkNDC
#:RRRRRRRR-R-RRRRRRBRRm51]j23jR4=R3Rj
RRRRR-RR-FR7lMNH:R
RRRRRR-R-RRRRRRRRRHXRM R)qRp
RRRRR-RR-sR sRFsO8FMHF0HM
#:RRRRRRRR-R-RRRRRRhRRF
MCRRRRRRRR-)-RNCMo:R
RRRRRR-R-RRRRRRRRR1Bm]25XRR>=4
3jRRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRRRN2aRECkL#ND8CRFHlNMVRFR1Bm]#RHRbNbsHFGlCN0Do$RHMPCR:L$
RRRRRRRRR--RRRRRRRRRRRRRqRRAX152=R<Rtpm5q) pQ']t
]2
RRRRMVkOF0HMqRah5]RXRR:H)MR 2qpR0sCkRsM)p q;R
RRRRRR-R-RsukbCF#:R
RRRRRR-R-RRRRRRRRR0)Ck#sMRbE$CFsLDRHO0oNMCRM0FXVR
RRRRRRRRR--1ObCHRNDPkNDC
#:RRRRRRRR-R-RRRRRRaRRq5h]j23jRj=R3Rj
RRRRR-RR-FR7lMNH:R
RRRRRR-R-RRRRRRRRRHXRM R)qRp
RRRRR-RR-sR sRFsO8FMHF0HM
#:RRRRRRRR-R-RRRRRRhRRF
MCRRRRRRRR-)-RNCMo:R
RRRRRR-R-RRRRRRRRR1qA5haq]25X2=R<Rj43
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRRFRhM
C
RRRRVOkM0MHFRBq)1]QhRR5X:MRHRq) ps2RCs0kM R)q
p;RRRRRRRR-u-RkFsb#
C:RRRRRRRR-R-RRRRRR)RRCs0kMH#RMsPC#ECR$sbCLHFDOHR#MFCRV
RXRRRRRRRR-1-RbHCONPDRNCDk#R:
RRRRR-RR-RRRRRRRR)RqBh1Q]35jj=2RRjj3
RRRRRRRRR--7NFlH
M:RRRRRRRR-R-RRRRRRXRRRRHM)p q
RRRRRRRRR-- FsssFROM08HH#FM:R
RRRRRR-R-RRRRRRRRRMhFCR
RRRRRR-R-RM)No
C:RRRRRRRR-R-RRRRRRqRR)QB1hX]52#RHR0lNENCl0NHODRD$kFMLkCM88R
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRRNRR2ERaCCRsNNOELRDCsoNMCVRFRBq)1]QhRRH#NsbbFlGHND0C$HRoPRCML
$:RRRRRRRR-R-RRRRRRRRRRRRRRARq1)5qBh1Q]25X2=R<Rtpm5q) pQ']t
]2
RRRRMVkOF0HM)RqB1Bm]XR5RH:RM R)qRp2skC0s)MR ;qp
RRRRRRRRR--ubksF:#C
RRRRRRRRR--RRRRRRRR)kC0sRM#HCMPsR#CEC$bsDLFHOORFM#HCVRFRRX
RRRRR-RR-bR1CNOHDNRPD#kC:R
RRRRRR-R-RRRRRRRRRBq)B]m15j432RR=j
3jRRRRRRRR-7-RFHlNMR:
RRRRR-RR-RRRRRRRRRRX>4=R3Rj
RRRRR-RR-sR sRFsO8FMHF0HM
#:RRRRRRRR-R-RRRRRR RRsssFRRHVXRR<4
3jRRRRRRRR-)-RNCMo:R
RRRRRR-R-RRRRRRRRRBq)B]m15RX2>j=R3Rj
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRRRRNa2REkCRbsbCRkLFMF8RVER0CCRsNNOELRDCsoNMCVRFRBq)B]m1R
H#RRRRRRRR-R-RRRRRRRRRRbRNbGsFH0lNCRD$oCHPM$RL:RRRqB)Bm51]X<2R=mRpt 5)q]p'Q2t]
R
RRkRVMHO0FqMR)qBah5]RXRR:H)MR 2qpR0sCkRsM)p q;R
RRRRRR-R-RsukbCF#:R
RRRRRR-R-RRRRRRRRR0)Ck#sMRPHMCCs#RbE$CFsLDRHO0oNMCRM0FXVR
RRRRRRRRR--1ObCHRNDPkNDC
#:RRRRRRRR-R-RRRRRRqRR)qBahj]53Rj2=3RjjR
RRRRRR-R-Rl7FN:HM
RRRRRRRRR--RRRRRRRRq5A1X<2RRj43
RRRRRRRRR-- FsssFROM08HH#FM:R
RRRRRR-R-RRRRRRRRRs sFHsRVARq125XRR>=4
3jRRRRRRRR-)-RNCMo:R
RRRRRR-R-RRRRRRRRRBq)a]qh5RX2Hl#RNC0ElHN0ODND$MRkLMFk8
C8RRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRRRN2aRECsOCNEDNLCNRsMRoCFqVR)qBahH]R#bRNbGsFH0lNCRD$oCHPM$RL:R
RRRRRR-R-RRRRRRRRRRRRRRRRq5A1qa)Bq5h]XR22<mRpt 5)q]p'Q2t]
V
Sk0MOHRFMPF_OsO8H_8lFCF_s0HN0FXM5js:RC;NDRRYj:CRsNRD;Z:jRRNsCDS;
S:MRR0MNkDsN;CRs0RR:MkN0s2NDR0sCkRsM)p qRR=>"sOF8_HOlCF8_0sFNF0HM
";
8CMRqRva)]_ ;qp
N
bOo	NCFRL8v$Rq_a])p qR
H#
RRRR
--RRRR-p-RFDONRMBF#M0N0V#RFzsR#HCRMER0CNRuOo	NCFRA8m$RM
D$RRRR-R-
RORRF0M#NRM0Ravq]__ u:.RR R)q:pR=3R(djUg6j_ng_Ugd6jnjR;RRR--C.**
RRRRMOF#M0N0vRRqBX_mazh:hRQa  t)=R:Rj46;-R-RGvNHllkRkOFMV0RFMsRkClLsVRFRH0sCR#
RORRF0M#NRM0Ravq]Q_ t_]au:QRRq) p=R:R3.64(d.c._4._U(4cUd6j_g(_(j4;46RU--*
bHRRRRO#FM00NMRqRvXa_Q R):RaQh )t RR:=.R(;RR--vHNGlRklbOsCHF#HMNRVOs0FRsVFRsOF8
HORRRRO#FM00NMRqRva ]__ju4RR:R)p qRR:=...jnn3c6_(gcnUj((_4;-R-R*C*4Rj
RORRF0M#NRM0RRiB: R)q:pR=3Rnj6(..6gdjUjUU.4cC4-j;-R-RMBF#M0N0FRVsFROsO8H
RRRRMOF#M0N0ARRq_1  :u1Rq) p=R:Rjj3j4jj;-RR-NRwOs0FRsVFRMOFPoCsCCMORHOs0HCsNR

R-RR-R
RR-R-ROpFNaDR$RbC7DCON0sNH#FMRsVFRsBF8RHOmsbCNF0HMR#
R-RR-R
RR$R0bBCRmQ)7Bm_v7a _YRu H5#R)qmaahQm, ReB)amQ2ht;R
RR$R0b)CR _qpea BmH)R#sRNsRN$5ahqzp)qRMsNo<CR>F2RV R)q
p;RRRR0C$bRahqzp)q_Be aRm)HN#Rs$sNRq5haqz)pNRsMRoC<R>2FhVRq)azq
p;RRRR#0kL$RbC)p q_)q)_H.R# R)qep_ mBa)jR5RR0F4
2;RRRR#0kL$RbC)p q_)q)_HdR# R)qep_ mBa)jR5RR0F.
2;RRRR#0kL$RbC)p q_Be a_m)h#RHRq) p _eB)amRR5j0vFRqQX_a2 );R
RRkR#Lb0$CzRTqq7)hHaR#hRQa  t)NRsMRoCjFR0R
d;
RRRR
--RRRR-q-RkDGHH$NsRMwkOF0HMV#RFBsRFHs8ODRqoHFs0#El
RRRR
--RRRRVOkM0MHFRWum m)_w__.1Q ) 51R7RR:HhMRq)azqep_ mBa)Q;RhQQaqep_q pzRH:RM R)q
p;RRRRRRRRRRRRRRRRhAzv m)_wq_ep1z RH:RMqRhaqz)ps2RCs0kM R)qep_ mBa)#RH
RRRRRRRRR--7OC#s0HbH:FM
RRRRRRRRR--RRRRR)RRCs0kMb#RFsICRRFV0RIFVRFsNCRPOs0FRRFVPkNDCR#
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRhRRF
MCRRRRRRRR-R-
RRRRRPRRNNsHLRDCeRR:)p q_Be aRm)50jRFzRhv)A __mwezqp ;12
RRRRRRRRsPNHDNLC Rav:uRRq) p=R:RQQhapQq_peqz
 ;RRRRRRRRPHNsNCLDRqwptRR:Apmm Rqh:a=R);z 
RRRRoLCHRM
RRRRRRRRRRRRRsVFRHQRMRRj0hFRz vA)w_m_peqzR 1DbFF
RRRRRRRRRRRRRRRR5ReQ:2R= Rav
u;RRRRRRRRRRRRRRRRRsVFRHuRM'R7)tqh FRDFRb
RRRRRRRRRRRRRRRRRRRRRRRRRHRRVRRQ=5R7u02RE
CMRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRwtpqRR:=w1qp R;
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRCRRG;H0
RRRRRRRRRRRRRRRRRRRRRRRRRRRR8CMR;HV
RRRRRRRRRRRRRRRRMRC8FRDF
b;RRRRRRRRRRRRRRRRRRHVwtpqRC0EMR
RRRRRRRRRRRRRRRRRRRRRRRRRR Rav:uR= Rav.u/3
j;RRRRRRRRRRRRRRRRR8CMR;HV
RRRRRRRRRRRRRRRRpRwq:tR=)Raz
 ;RRRRRRRRRRRRRMRC8FRDF
b;RRRRRRRRRRRRRCRs0MksR
e;RRRRCRM8u mW)w_m_1._  )Q1
;

RRRRMOF#M0N0WRama_q_hvQz:1RRq) p _eB)amRR:=u mW)w_m_1._  )Q1R5
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRqRhaqz)p _eB)am'j54jg,Rj42,3
j,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRqRvXa_Q ;)2
R
RRFROMN#0M 0Rup1Qm:hRRq) p _eB)am_:hR=
R5RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR(63Ud4gUngdd(Ucc.-(Cj
4,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRcd3nnnc(jjgjjnUjj-nCj
4,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR.c3cgn(Un.d4ncUn4-dCj
4,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR4c3.dg6cgcc6n4(nc-cCj
4,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRnc3.4jUUg6gggd6(6-4Cj
.,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRd.34ddgUdjcd..nU(-(Cj
.,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR4n36..d(Ujn.cU(nd-jCj
.,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR(43U.4dcj4njj4444-nCj
d,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRdj3gnj.d4gd4n(ng4-(Cj
d,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR463gd.4.6c4n(4UUU-gCj
d,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRgn3(64n.U6g6ggd4d-(Cj
c,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRcU3U..U44g44cUUg.-gCj
c,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR.c3c4ncj.cj4g4dn(-6Cj
c,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR4.3.jd(j4g4Udjn(.-4Cj
c,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRnj34d664nc4(.(jUn-UCj
6,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRd63j4((6U6446j.ng-dCj
6,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR4.366UU(g4jnd(46n-jCj
6,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR(.3ngcdg64d4jn4gg-gCj
n,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRd43Uc(ng.nn6jgncn-jCj
n,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR4j3g(UdcnUd.4Uj4(-jCj
n,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRgd36nd(c4jnc6jgnU-jCj
(,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRcn3(U4d(6jU.dUjU(-nCj
(,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR.U3dc64U(jg44U66j-4Cj
(,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR4g34..jgU6g6jj(Un-(Cj
(,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR6n3gjccnc6((d6gj6-dCj
U,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR.U3gj..d.(dUndg6j-dCj
U,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR4g3cjn444d4gUnc(6-cCj
U,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR(63cjj6U6ggn..dUU-4CjRg
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR;R2
R
RRkRVMHO0FBMRmQ)7BRR5X:jRRRHM)p q;R
RRRRRRRRRRRRRRRRRRRRRY:jRRRHM)p q;R
RRRRRRRRRRRRRRRRRRRRRZ:jRRRHM)p q;R
RRRRRRRRRRRRRRRRRRRRRhRR:HhMRq)azqRp;RRRRRRRRRRRRRRRR-R-RuOsCHF#HMNRVOs0F
RRRRRRRRRRRR)Bm7_QBv m7RH:RMmRB)B7Q_7vm Y_auR RRRRRR-RR-)RRF00NHRFM5-ZR>2Rj
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-FRRsCRPOs0FHRMo5-YR>2Rj
RRRRRRRRRRRRRRRRRRRRs2RCs0kM R)qqp_)d)_R
H#RRRRRRRR-7-RCs#OHHb0F
M:RRRRRRRR-R-RRRRRRFRBl0bkCFROsO8HRDPNk
C#RRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRRMhFCR
RRRRRRRRRRPRRNNsHLRDCXRR:)p qRR:=X
j;RRRRRRRRRRRRRsPNHDNLCRRY: R)q:pR=jRY;R
RRRRRRRRRRPRRNNsHLRDCZRR:)p qRR:=Z
j;RRRRRRRRRRRRRsPNHDNLC_RXau vR):R ;qp
RRRRoLCHRM
RRRRRVRHR)Bm7_QBv m7R)=RmaaqQRmh0MEC
RRRRRRRRRRRVRFsiMRHR0jRFRRhDbFF
RRRRRRRRRRRRRRRRRRRRXRR_va u=R:R
X;RRRRRRRRRRRRRRRRRRRRRVRHRZ5RRR>=j23jRC0EMR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRR:XR=RRX-RRY*WRama_q_hvQzi152R;
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRY:Y=RRX+R_va uRR*a_Wmqva_Q1hz5;i2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRZ=R:R-ZRR1 uQhpm5;i2
RRRRRRRRRRRRRRRRRRRRCRRD
#CRRRRRRRRRRRRRRRRRRRRRRRRRRRRRXRRRR:=XRR+YRR*a_Wmqva_Q1hz5;i2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRY=R:R-YRRaX_ Rvu*WRama_q_hvQzi152R;
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRZ:Z=RR +Rup1Qmih52R;
RRRRRRRRRRRRRRRRRRRRR8CMR;HV
RRRRRRRRRRRR8CMRFDFbR;
RRRRRCRRD
#CRRRRRRRRRRRRVRFsiMRHR0jRFRRhDbFF
RRRRRRRRRRRRRRRRRRRRaX_ Rvu:X=R;R
RRRRRRRRRRRRRRRRRRVRHRY5RRj<R3Rj20MEC
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRX=R:R-XRR*YRRmaW__qavzQh125i;R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRR:YR=RRY+_RXau vRa*RWqm_aQ_vh5z1i
2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRZRRRR:=ZRR- Qu1p5mhi
2;RRRRRRRRRRRRRRRRRRRRCCD#
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRX=R:R+XRR*YRRmaW__qavzQh125i;R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRR:YR=RRY-_RXau vRa*RWqm_aQ_vh5z1i
2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRZRRRR:=ZRR+ Qu1p5mhi
2;RRRRRRRRRRRRRRRRRRRRCRM8H
V;RRRRRRRRRRRRCRM8DbFF;R
RRRRRRMRC8VRH;R
RRRRRRCRs0MksRq) p)_q)'_d5RX,YZ,R2R;
RCRRMB8RmQ)7B
;
RRRR-R-
R-RR-FRA8#HCRsVFRFtDLRNDvEN0C0lNHDONRMwkOF0HM1#R00NsRs]CCR
RR-R-
RRRRMVkOF0HMQR1t5hRXH:RM R)q2pRR0sCkRsM)p qR
H#RRRRRRRR-7-RCs#OHHb0F
M:RRRRRRRR-R-RRRRRRCR1CkRVMHO0F8MRCNODsHN0FHMRM RQ 1 R048Rj3(n.g-4gRn
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRhRRF
MCRRRRLHCoMR
RRRRRRRRRRRHVRX5RRj>R32jRRER0CRM
RRRRRRRRRRRRRsRRCs0kM3R4jR;
RRRRRRRRRDRC#RHV5RRX<3RjjRR2RC0EMR
RRRRRRRRRRRRRRCRs0MksR3-4jR;
RRRRRRRRRDRC#RC
RRRRRRRRRRRRRsRRCs0kM3RjjR;
RRRRRRRRRMRC8VRH;R
RRMRC8QR1t
h;
RRRRMVkOF0HM RBQ5pRXRR:H)MR Rqp2CRs0MksRq) p#RH
RRRRRRRRR--7OC#s0HbH:FM
RRRRRRRRR--RRRRR1RRCVCRk0MOHRFM8DCON0sNHRFMHQMR R  1R084nj(34.-g
gnRRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRNh2RFFROMsPC#MHFRR0FNQMRhta  0)R$RbCHC#RGObC0,C8RR#F0MskOCN0
RRRRRRRRR--RRRRRRRRRNROM0MFRCFPsFVDIFRVsNRDsRoCNksol0CM#R
RRRRRR-R-RRRRRRRRLa2RE8CRFHlNMkR#bsbF0RC8L0$RERH#VOkM0MHFRRH#X=R<R)pqtR 
RRRRR-RR-RRRRRRRRRO2)kC0sRM#XVRHR1qA5RX2>p=Rq )t
R
RRRRRRFROMN#0Mp0Rq )t: R)qRpR:)=R 5qpQ hat' )]]Qt2R;
RRRRRPRRNNsHLRDC)R7:)p q;R

RLRRCMoH
RRRRRRRRVRHR1qA5RX2>p=Rq )tRC0EMR
RRRRRRRRRRRRRR0sCkRsMXR;
RRRRRRRRCRM8H
V;
RRRRRRRR7R)RR:=)p qRQ5Rhta  X)52
2;RRRRRRRRRRHV)=7RR0XRE
CMRRRRRRRRRRRRskC0s)MR7R;
RRRRRRRRCRM8H
V;
RRRRRRRRRRRRRHVXRR>jR3j0MEC
RRRRRRRRRRRRRRRRRRRRRRRH)VR7=R>R0XRE
CMRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRCRs0MksR;)7
RRRRRRRRRRRRRRRRRRRRRRRCCD#
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRsRRCs0kM7R)R4+R3
j;RRRRRRRRRRRRRRRRRRRRRCRRMH8RVR;
RRRRRRRRRCRRDV#HRRRX=3Rjj0RRE
CMRRRRRRRRRRRRRRRRskC0sjMR3
j;RRRRRRRRRRRRCCD#
RRRRRRRRRRRRRRRRRRRRRRRH)VR7=R<R0XRE
CMRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRCRs0MksRR)7+3R4jR;
RRRRRRRRRRRRRRRRRRRRRDRC#RC
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR0sCkRsM)
7;RRRRRRRRRRRRRRRRRRRRRCRRMH8RVR;
RRRRRRRRRCRRMH8RVR;
RCRRMB8R ;Qp
R
RRkRVMHO0FwMRp)mmRR5X:MRHRq) pRR2skC0s)MR RqpHR#
RRRRR-RR-CR7#HOsbF0HMR:
RRRRR-RR-RRRRRRRRC1CRMVkOF0HMCR8OsDNNF0HMMRHR Q  0R18jR4(.n3-g4gnR
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRR2RNRRhFOPFMCHs#F0MRFMRNRaQh )t Rb0$C#RHRbCGCCO08#,RFsR0kNMO0RC
RRRRR-RR-RRRRRRRRRRROMNMFF0RPVCsDRFIVRFsDoNsCsRNoCklM
0#RRRRRRRR-R-RRRRRR2RLRCaERl8FNRHM#bkbFCs08$RLRH0E#kRVMHO0FHMR#ARq125XRR<=ptq) R
RRRRRR-R-RRRRRRRRO)2RCs0kMX#RRRHVq5A1X>2R=qRp)
t 
RRRRRRRRMOF#M0N0qRp):t Rq) p:RR= R)qQp5hta  ])'Q2t];R
RRRRRRNRPsLHND)CR7):R ;qp
R
RRCRLo
HMRRRRRRRRHqVRAR15XRR2>p=Rq )tRC0EMR
RRRRRRRRRRRRRRRRRRCRs0MksR
X;RRRRRRRRCRM8H
V;
RRRRRRRRR)7:)=R Rqp5hRQa  t)25X2R;
RRRRRHRRV7R)RX=RRC0EMR
RRRRRRRRRRRRRRCRs0MksR;)7
RRRRRRRR8CMR;HV
R
RRRRRRVRHR>XRRjj3RC0EMR
RRRRRRRRRRRRRRRRRRRRRH)VR7=R<R0XRE
CMRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRCRs0MksR;)7
RRRRRRRRRRRRRRRRRRRRRRRCCD#
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRsRRCs0kM7R)R4-R3
j;RRRRRRRRRRRRRRRRRRRRRCRRMH8RVR;
RRRRRCRRDV#HRRRX=3Rjj0RRE
CMRRRRRRRRRRRRRRRRskC0sjMR3
j;RRRRRRRRCCD#
RRRRRRRRRRRRRRRRRRRH)VR7=R>R0XRE
CMRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRCRs0MksRR)7-3R4jR;
RRRRRRRRRRRRRRRRRDRC#RC
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR0sCkRsM)
7;RRRRRRRRRRRRRRRRRCRRMH8RVR;
RRRRRCRRMH8RVR;
RCRRMw8Rp)mm;R

RVRRk0MOHRFM)hmz7XR5RH:RM R)q2pRR0sCkRsM)p qR
H#RRRRRRRR-7-RCs#OHHb0F
M:RRRRRRRR-R-RRRRRRCR1CkRVMHO0F8MRCNODsHN0FHMRM RQ 1 R048Rj3(n.g-4gRn
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRRRRN)2RCs0kMj#R3HjRVRRX=3RjjR
RRRRRR-R-RRRRRRRRRRL2)kC0sRM#wmpm)R5X+3Rj6H2RVRRX>
RjRRRRRRRR-R-RRRRRRORR2CR)0Mks# RBQXp5Rj-R3R62HXVRRj<R
R
RRCRLo
HMRRRRRRRRRHRRVXRRRj>R3RjR0MEC
RRRRRRRRRRRRRRRR0sCkRsMwmpm)R5X+3Rj6
2;RRRRRRRRRCRRDV#HRRRX<3Rjj0RRE
CMRRRRRRRRRRRRRRRRskC0sBMR 5QpR-XRR6j32R;
RRRRRRRRRDRC#RC
RRRRRRRRRRRRRsRRCs0kM3RjjR;
RRRRRRRRRMRC8VRH;R
RRMRC8mR)z;h7
R
RRkRVMHO0FaMR)BzhRR5X:MRHRq) pRR2skC0s)MR RqpHR#
RRRRR-RR-CR7#HOsbF0HMR:
RRRRR-RR-RRRRRRRRC1CRMVkOF0HMCR8OsDNNF0HMMRHR Q  0R18jR4(.n3-g4gnR
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRRNRR2CR)0Mks#3RjjVRHR=XRRjj3
RRRRRRRRR--RRRRRRRRL)2RCs0kMw#Rp)mm5RX2HXVRRj>R
RRRRRRRRR--RRRRRRRRO)2RCs0kMB#R 5QpXH2RVRRX<
Rj
RRRRoLCHRM
RRRRRRRRRVRHRRRX>3Rjj0RRE
CMRRRRRRRRRRRRRRRRskC0swMRp)mm5;X2
RRRRRRRRRRRCHD#VXRRRj<R3RjR0MEC
RRRRRRRRRRRRRRRR0sCkRsMBp Q52RX;R
RRRRRRRRRR#CDCR
RRRRRRRRRRRRRRCRs0MksRjj3;R
RRRRRRRRRR8CMR;HV
RRRR8CMRza)h
B;



RRRRVOkM0MHFRm"v75"RXY,R:MRHRq) pRR2skC0s)MR RqpHR#
RRRRR-RR-CR7#HOsbF0HMR:
RRRRR-RR-RRRRRRRRC1CRMVkOF0HMCR8OsDNNF0HMMRHR Q  0R18jR4(.n3-g4gnR
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRR2RNR0)Ck#sMRjj3RRFMCFsssR

RRRRRPRRNNsHLRDCXth qeaQ RR:Apmm Rqh:X=RRj<R3
j;RRRRRRRRPHNsNCLDR YhtQqae: RRmAmph qRR:=YRR<j;3j
RRRRRRRRsPNHDNLCqRepRz : R)q
p;RRRRLHCoMR
RRRRRR-R-RCBEOP	RN8DHHR0$FHVRM0bkRoNskMlC0R#
RRRRRRRRRHRRVYR5Rj=R3Rj20MEC
RRRRRRRRRRRRRRRR#RN#0CsRpwq1R 
RRRRRRRRRRRRRRRRRRRRRsRRCsbF0vR"mX75,3RjjH2R#MRk8HCVM"C8
RRRRRRRRRRRRRRRRRRRRRRRRP#CC0sH$)R );m)
RRRRRRRRRRRRRRRRCRs0MksRjj3;R
RRRRRRRRRRRRRCRM8H
V;
RRRRRRRRR--BbFlkR0CPkNDCR
RRRRRRVRHRX5Rhq ta QeR02RE
CMRRRRRRRRRRRRRRRRH5VRR YhtQqae2 RRC0EMR
RRRRRRRRRRRRRRRRRRRRRRqRepRz :X=RR5+Rwmpm)A5q125X/1qA52Y22A*q125Y;R
RRRRRRRRRRRRRRDRC#RC
RRRRRRRRRRRRRRRRRRRRReRRq pzRR:=XRR+5QB pA5q125X/1qA52Y22A*q125Y;R
RRRRRRRRRRRRRRMRC8VRH;R
RRRRRRDRC#RC
RRRRRRRRRRRRRHRRVRR5Yth qeaQ RR20MEC
RRRRRRRRRRRRRRRRRRRRRRRRpeqz: R=RRX-BR5 5Qpq5A1Xq2/AY152*22q5A1Y
2;RRRRRRRRRRRRRRRRCCD#
RRRRRRRRRRRRRRRRRRRRRRRRpeqz: R=RRX-wR5p)mm51qA5/X2q5A1Y222*1qA5;Y2
RRRRRRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMR;HV
R
RRRRRRCRs0MksRpeqz
 ;RRRRCRM8"7vm"
;

RRRRMVkOF0HM R)qqpvXXR5,RRY:MRHRq) pRR2skC0s)MR RqpHR#
RRRRR-RR-CR7#HOsbF0HMR:
RRRRR-RR-RRRRRRRRC1CRMVkOF0HMCR8OsDNNF0HMMRHR Q  0R18jR4(.n3-g4gnR
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRR2RNRq) pXvq5YX,2RR=XERICXMRRY=R
RRRRRRRR
--RRRRLHCoMR
RRRRRRVRHR>XR=RRY0MEC
RRRRRRRRRRRskC0sXMR;R
RRRRRRDRC#RC
RRRRRRRRRCRs0MksR
Y;RRRRRRRRCRM8H
V;RRRRCRM8)p qv;qX
R
RRkRVMHO0F)MR vqpQ5hRXY,RRH:RM R)q2pRR0sCkRsM)p qR
H#RRRRRRRR-7-RCs#OHHb0F
M:RRRRRRRR-R-RRRRRRCR1CkRVMHO0F8MRCNODsHN0FHMRM RQ 1 R048Rj3(n.g-4gRn
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRNRR2 R)qQpvh,5XY=2RRIXRERCMXRR=YR
RRRRRR-R-
RRRRoLCHRM
RRRRRHRRVRRX<Y=RRC0EMR
RRRRRRRRRR0sCkRsMXR;
RRRRRCRRD
#CRRRRRRRRRsRRCs0kM;RY
RRRRRRRR8CMR;HV
RRRR8CMRq) phvQ;


RRRRbOsFCs8kChRzQ)wmvN5PsLHND1CR 4 7, 1 7H.:M0FkR1umQeaQ N;PsLHNDXCR:0FkRq) pR2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRHR#
RRRRR-RR-CR7#HOsbF0HMR:
RRRRR-RR-RRRRRRRRC1CRMVkOF0HMCR8OsDNNF0HMMRHR Q  0R18jR4(.n3-g4gnR
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRR2RNR0)Ck#sMRjj3RRFMCFsssR
RRRRRR-R-
RRRRRRRRsPNHDNLC,RZRRi:Q hat; )
RRRRRRRRsPNHDNLC1Ra 4 7RQ:Rhta  :)R=hRQa  t)1'5 4 72R;
RRRRRPRRNNsHLRDCa 1 7:.RRaQh )t RR:=Q hat' )5 1 7;.2
RRRRoLCHRM
RRRRR-RR-ERBCRO	PHND8$H0RRFVNksol0CM#R
RRRRRRVRHR 1 7>4RRc.4(dcU6Rn.0MEC
RRRRRRRRRRRRRRRR#N#CRs0w1qp R
RRRRRRRRRRRRRRRRRRRRRRCRsb0FsR "1 R74>4R.cU(cd.6nRRHMzwhQm")v
RRRRRRRRRRRRRRRRRRRRRRRRP#CC0sH$)R );m)
RRRRRRRRRRRRRRRR:XR=3RjjR;
RRRRRRRRRRRRRsRRCs0kMR;
RRRRRCRRMH8RV
;
RRRRRRRRH1VR . 7R.>R4cc(UgddUER0CRM
RRRRRRRRRRRRRNRR#s#C0qRwp
1 RRRRRRRRRRRRRRRRRRRRRRRRsFCbs"0R17  .RR>.(4ccdUdgHURMhRzQ)wmvR"
RRRRRRRRRRRRRRRRRRRRR#RRCsPCHR0$ m)))R;
RRRRRRRRRRRRRXRRRR:=j;3j
RRRRRRRRRRRRRRRR0sCk;sM
RRRRRRRR8CMR;HV
R
RRRRRR-R-RlBFbCk0RIMCRC#C8NRPD#kCR8NMRCb#k-8Fs8NMFMlRkClLsR
RRRRRRRRi:a=R17  4d/6n;nU
RRRRRRRR a1 R74:c=Rjcj4R5*Ra 1 7-4RR*iRRn6dnRU2-RRi*.R4.;44
R
RRRRRRVRHR a1 R74<RRjRC0EMR
RRRRRRRRRRRRRR1Ra 4 7RR:=a 1 7+4RRc.4(dcU6;nd
RRRRRRRR8CMR;HV
R
RRRRRRRRi:a=R17  ../6(;(c
RRRRRRRR a1 R7.:c=Rj.ngR5*Ra 1 7-.RR*iRR(6.(Rc2-RRi*(Rdg
4;
RRRRRRRRRHVa 1 7<.RRRjR0MEC
RRRRRRRRRRRRRRRR a1 R7.:a=R17  .RR+.(4ccdUdg
g;RRRRRRRRCRM8H
V;
RRRRRRRR:ZR=1Ra 4 7Ra-R17  .R;
RRRRRHRRVRRZ<RR40MEC
RRRRRRRRRRRRRRRR:ZR=RRZ+4R.cU(cd.6n;R
RRRRRRMRC8VRH;R

RRRRR-RR-CRt0kRF00bkRDPNk
C#RRRRRRRR17  4=R:R1umQeaQ a'517  4
2;RRRRRRRR17  .=R:R1umQeaQ a'517  .
2;RRRRRRRRX=R:R R)qZp523*cnn6n4-dC4
j;RRRRCRM8zwhQm;)v



RRRRVOkM0MHFR)1TaXR5RH:RM R)q2pRR0sCkRsM)p qR
H#RRRRRRRR-7-RCs#OHHb0F
M:RRRRRRRR-R-RRRRRRCR1CkRVMHO0F8MRCNODsHN0FHMRM RQ 1 R048Rj3(n.g-4gRn
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRNRR2#RzC0#REhCRCFI0MN-)bFE#MbRNbGsFH0lNH:FM
RRRRRRRRR--RRRRRRRRRwRR54M+2RR=j*36rMw52RR+G5/wM
29RRRRRRRR-R-RRRRRR2RLR0)Ck#sMRjj3RRFMCFsssR
RRRRRR-R-
R
RRRRRRFROMN#0M 0Ru:1RRq) p=R:R1Aq u_ 1q*A1  _uR1;-B-RFCMPsMoCOVCRNFO0sR

RRRRRPRRNNsHLRDCQehQqRp:)p q;R
RRRRRRNRPsLHNDmCRpq7epRR:)p qRR;
RRRRRPRRNNsHLRDChe Wq:pRRq) p
R;RRRRRRRRPHNsNCLDRzBmh:aRRaQh )t RR:=4
;
RRRRLHCoMR
RRRRRR-R-RCBEOP	RN8DHHR0$FNVRslokC
M0RRRRRRRRH5VRR<XRRjj3R02RE
CMRRRRRRRRRRRRRRRRNC##sw0Rq p1
RRRRRRRRRRRRRRRRRRRRRRRRbsCFRs0"<XRRjj3RRHM1aT)5"X2
RRRRRRRRRRRRRRRRRRRRRRRRP#CC0sH$)R );m)
RRRRRRRRRRRRRRRR0sCkRsMj;3j
RRRRRRRR8CMR;HV
R
RRRRRR-R-R0tCRC0ERk#JNRsCs0FFRsVFRC#bODHNR#ONCR#
RRRRRHRRVRRX=3RjjER0CRM
RRRRRRRRRRRRRRRRR0sCkRsMj;3j
RRRRRRRR#CDCR
RRRRRRRRRRRRRRVRHRX5RR4=R32jRRC0EMR
RRRRRRRRRRRRRRRRRRRRRRCRs0MksRj43;R
RRRRRRRRRRRRRRMRC8VRH;R
RRRRRRMRC8VRH;R

RRRRR-RR-CRt0ER0CJR#kCNsRFsF0FRVsCRoMNCsDNRO#
C#RRRRRRRRQehQq:pR=XR um5pt25X*35j6;22RR--vEN0C0lNHDONDO$RFCssOL0RkH0RlCbsOCH#
RRRRRRRR7mpeRqp:Q=RhqQepR;
RRRRRhRR qWep=R:R/5Xmep7q+pRR7mpe2qp*6j3;R

RRRRR-RR-ERBCRO	VRFsRDsCNP0HCMRN8LRN#kFD0CCRsssFR8NMRGlNRkOFMR0
RRRRRIRRECHDRRR55qR5A515he Wq-pRmep7q/p2he WqRp2>uR 1m2R)R
RRRRRRRRRRRRRRRRRRA5q1 5hWpeqRm-Rpq7ep>2RR1 u2RR2q
h7RRRRRRRRRRRRRRRRR5RRBhmzaRR<v_qXBhmza22RRFRDFRb
RRRRRRRRRRRRRmRRpq7ep=R:RWh e;qp
RRRRRRRRRRRRRRRRWh eRqp:5=RXp/m7peqRm+Rpq7epj2*3
6;RRRRRRRRRRRRRRRRBhmza=R:RzBmh+aRR
4;RRRRRRRRCRM8DbFF;R
RRRRRRCRs0MksRWh e;qp
RRRR8CMR)1Ta
;
RRRRVOkM0MHFR)BAaXR5RH:RM R)q2pRR0sCkRsM)p qR
H#RRRRRRRR-7-RCs#OHHb0F
M:RRRRRRRR-R-RRRRRRCR1CkRVMHO0F8MRCNODsHN0FHMRM RQ 1 R048Rj3(n.g-4gRn
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRNRR2#RzC0#REhCRCFI0MN-)bFE#MbRNbGsFH0lNH:FM
RRRRRRRRR--RRRRRRRRRwRR54M+2RR=5d4/2.*r*Mw52RR+G5/wM*2*.
9;RRRRRRRR-R-
RRRRRORRF0M#NRM0 Ru1: R)q:pR=qRA1  _uA1*q_1  ;u1
R
RRRRRRNRPsLHNDQCRhqQep):R ;qp
RRRRRRRRsPNHDNLCpRXmpBqR):R Rqp:X=R;R
RRRRRRNRPsLHNDhCR atqQRe :mRAmqp h=R:R<XRRjj3;R
RRRRRRNRPsLHNDmCRpq7epRR:)p qRR;
RRRRRPRRNNsHLRDChe Wq:pRRq) p
R;RRRRRRRRPHNsNCLDRzBmh:aRRaQh )t RR:=4
;
RRRRLHCoMR

RRRRR-RR-FRBl0bkCFRsFV0RF#sRbHCONODRN##C
RRRRRRRRRHVXRR=jR3j0MEC
RRRRRRRRRRRRRRRR0sCkRsMj;3j
RRRRRRRR#CDH5VRR=XRRj43R02RE
CMRRRRRRRRRRRRRRRRskC0s4MR3
j;RRRRRRRRCCD#
RRRRRRRRRRRRRRRRRHVXRR=-j43RC0EMR
RRRRRRRRRRRRRRRRRRRRRRCRs0MksR3-4jR;
RRRRRRRRRRRRRCRRMH8RVR;
RRRRRCRRMH8RV
;
RRRRRRRR-B-RFklb0sCRFRF0VRFsoCCMsRNDOCN##R
RRRRRRVRHRth qeaQ ER0CRM
RRRRRRRRRRRRRXRRpqmBp=R:R;-X
RRRRRRRR8CMR;HV
R
RRRRRRhRQQpeqRR:= 5Xup5mtXBpmq/p25jd32R2;-v-RNC0ElHN0ODND$FROsOsC0kRL0R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-H-RlCbsOCH#
RRRRRRRR7mpeRqp:Q=RhqQepR;
RRRRRhRR qWep=R:Rp5XmpBq/p5m7peq*7mpe2qpR.+R3mj*pq7epd2/3
j;
RRRRRRRRR--BOEC	FRVsCRsDHN0PNCRMN8RLD#FkR0CCFsssN#RMl8RNOGRF0kM
RRRRRRRRHIED5CRRR5R51qA5 5hWpeqRp-m7peq2 /hWpeq2RR> Ru12)Rm
RRRRRRRRRRRRRRRRRRR51qA5Wh eRqp-pRm7peq2RR> Ru12RR2R7qh
RRRRRRRRRRRRRRRRRRR5mRBzRha<qRvXm_BzRha2RR2DbFF
RRRRRRRRRRRRRRRR7mpeRqp:h=R qWepR;
RRRRRRRRRRRRRhRR qWep=R:5mXpB/qp57mpe*qpmep7qRp2+3R.jp*m7peq23/djR;
RRRRRRRRRRRRRBRRmazhRR:=BhmzaRR+4R;
RRRRRCRRMD8RF;Fb
R
RRRRRRVRHRth qeaQ ER0CRM
RRRRRRRRRRRRRhRR qWep=R:R -hWpeq;R
RRRRRRMRC8VRH;R

RRRRRsRRCs0kM RhWpeq;R
RRMRC8ARB)
a;
RRRRMVkOF0HM*R"*5"RXRR:HQMRhta  R);YRR:H)MR 2qpR0sCkRsM)p qR
H#RRRRRRRR-7-RCs#OHHb0F
M:RRRRRRRR-R-RRRRRRCR1CkRVMHO0F8MRCNODsHN0FHMRM RQ 1 R048Rj3(n.g-4gRn
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRNRR2CR)0Mks#3RjjMRFRsCsFOsRFHM80MHF
R
RRCRLo
HMRRRRRRRR-B-RE	CORDPNH08H$VRFRoNskMlC0R
RRRRRRVRHR55RR<XRRRjR2MRN8RR5Y=R/Rjj3R22RRC0EMR
RRRRRRRRRRRRRR#RN#0CsRpwq1R 
RRRRRRRRRRRRRRRRRRRRRsRRCsbF0XR"Rj<RR8NMR/YR=3RjjMRHR*X*YR"
RRRRRRRRRRRRRRRRRRRRR#RRCsPCHR0$ m)))R;
RRRRRRRRRRRRRsRRCs0kM3RjjR;
RRRRRCRRMH8RV
;
RRRRRRRRH5VRRX5RRj=RRRR2NRM85RRY<j=R32jRR02RE
CMRRRRRRRRRRRRRRRRNC##sw0Rq p1
RRRRRRRRRRRRRRRRRRRRRRRRbsCFRs0"=XRRNjRMY8RRR<=jR3jHXMR*"*Y
RRRRRRRRRRRRRRRRRRRRRRRRP#CC0sH$)R );m)
RRRRRRRRRRRRRRRR0sCkRsMj;3j
RRRRRRRR8CMR;HV
R
RRRRRR-R-R0tCRDPNkVCRF#sRbHCONODRN##C
RRRRRRRRRHV5RRX=RRjR8NMRRRY>3RjjRR20MEC
RRRRRRRRRRRRRRRR0sCkRsMj;3j
RRRRRRRR8CMR;HV
R
RRRRRRVRHRX5RR4=RR02RE
CMRRRRRRRRRRRRRRRRskC0s4MR3
j;RRRRRRRRCRM8H
V;
RRRRRRRRRHV5RRY=3RjjMRN8RRX/j=RR02RE
CMRRRRRRRRRRRRRRRRskC0s4MR3
j;RRRRRRRRCRM8H
V;
RRRRRRRRRHV5RRY=3R4j02RE
CMRRRRRRRRRRRRRRRRskC0s5MR)p q52X2;R
RRRRRRMRC8VRH;R

RRRRR-RR-CRt0NRPDRkCVRFsoCCMsRNDOCN#
RRRRRRRR0sCkRsM RXu5*YRRtpmR 5)qXp52;22
RRRR8CMR*"*"
;
RRRRVOkM0MHFR*"*"XR5RH:RM R)qRp;YRR:H)MR 2qpR0sCkRsM)p qR
H#RRRRRRRR-7-RCs#OHHb0F
M:RRRRRRRR-R-RRRRRRCR1CkRVMHO0F8MRCNODsHN0FHMRM RQ 1 R048Rj3(n.g-4gRn
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRNRR2CR)0Mks#3RjjMRFRsCsFOsRFHM80MHF
R
RRCRLo
HMRRRRRRRR-B-RE	CORDPNH08H$VRFRoNskMlC0R
RRRRRRVRHR55RR<XRRjj3RRR2NRM85RRY/j=R32jRR02RE
CMRRRRRRRRRRRRRRRRNC##sw0Rq p1
RRRRRRRRRRRRRRRRRRRRRRRRbsCFRs0"<XRRjj3R8NMR/YR=3RjjMRHR*X*YR"
RRRRRRRRRRRRRRRRRRRRR#RRCsPCHR0$ m)))R;
RRRRRRRRRRRRRsRRCs0kM3RjjR;
RRRRRCRRMH8RV
;
RRRRRRRRH5VRRX5RRj=R3RjR2MRN8RR5Y=R<Rjj3R22RRC0EMR
RRRRRRRRRRRRRR#RN#0CsRpwq1R 
RRRRRRRRRRRRRRRRRRRRRsRRCsbF0XR"Rj=R3NjRMY8RRR<=jR3jHXMR*"*Y
RRRRRRRRRRRRRRRRRRRRRRRRP#CC0sH$)R );m)
RRRRRRRRRRRRRRRR0sCkRsMj;3j
RRRRRRRR8CMR;HV
R
RRRRRR-R-R0tCRDPNkVCRF#sRbHCONODRN##C
RRRRRRRRRHV5RRX=3RjjNRRMR8RYRR>jR3j2ER0CRM
RRRRRRRRRRRRRsRRCs0kM3RjjR;
RRRRRCRRMH8RV
;
RRRRRRRRH5VRR=XRRj43R02RE
CMRRRRRRRRRRRRRRRRskC0s4MR3
j;RRRRRRRRCRM8H
V;
RRRRRRRRRHV5RRY=3RjjMRN8RRX/j=R32jRRC0EMR
RRRRRRRRRRRRRRCRs0MksRj43;R
RRRRRRMRC8VRH;R

RRRRRHRRVRR5YRR=423jRC0EMR
RRRRRRRRRRRRRRCRs0MksR25X;R
RRRRRRMRC8VRH;R

RRRRR-RR-CRt0NRPDRkCVRFsoCCMsRNDOCN#
RRRRRRRR0sCkRsM RXu5*YRRtpmR25X2R;
RCRRM"8R*;*"
-
-ApzQazQh1R 7RVRRk0MOHRFM RXuRR5X:MRHRq) pRR2skC0s)MR RqpH-#
-QAzphaQz71 RRRRRRRR-7-RCs#OHHb0F
M:-z-AQQpah z17RRRRRRRRR--RRRRR1RRCVCRk0MOHRFM8DCON0sNHRFMHQMR R  1R084nj(34.-g
gn-z-AQQpah z17RRRRRRRRR--hCF0#-:
-QAzphaQz71 RRRRRRRR-R-RRRRRR2RNRHaE#kRVMHO0FOMRFklb0RC#0RECCFGbM0CMHRNDkM#HoER0CFRVDIDFH
Mo-z-AQQpah z17RRRRRRRRR--RRRRRRRRRCR#s#HC:-
-ApzQazQh1R 7RRRRR-RR-RRRRRRRRRRRRRRRRbCG5RG2=RR4+RRG+*RG*../!RR+Gd**/Rd!+3R33RR;|RG|<3R4j-
-ApzQazQh1R 7RRRRR-RR-RRRRRRRRRRRNRM8skC8ORC#Nksol0CMR0XRFNR0	NCR8MPN0CNoRRFVC5GbG2+$R-=
-QAzphaQz71 RRRRRRRR-R-RRRRRRRRRRbCG5*G2C5Gb$-2
-QAzphaQz71 RRRRRRRR---
-QAzphaQz71 RRRRRRRR-R-RRRRRR2RLRHaE#lRHblDCCNM00MHFRlDHHR0#XFR0RRLCD#C#RN0EMmRpt 5)q]p'Q2t]
A--zaQpQ1hz R7RRRRRR-R-RRRRRRRRR0RRFPRNFRH8FsPCVIDF3)RRCs0kM)#R 'qp]]QtRCIEMRRXsOCNERC#00EN
A--zaQpQ1hz R7RRRRRR-R-RRRRRRRRRDRRH0lH
A--zaQpQ1hz R7RRRRRR-R-
A--zaQpQ1hz R7RRRRRRFROMN#0M 0Ru:1RRq) p=R:R1Aq u_ 1q*A1  _uA1*q_1  ;u1-u-RsHCO#MHFRHOs0HCsN-
-ApzQazQh1
 7-z-AQQpah z17RRRRRRRRRRRRsPNHDNLC R)B)QumpBq:mRAmqp h=R:R<XRRjj3;R--BOEC	HR#oFMRVsRNoCklM-0
-QAzphaQz71 RRRRRRRRRRRRPHNsNCLDRmXpBRqp: R)q:pR=ARq125X;RRRRRRR-z-R#bCRF0#HHRPCPkNDC-
-ApzQazQh1R 7RRRRRRRRRPRRNNsHLRDCmep7qRp:)p qR-;
-QAzphaQz71 RRRRRRRRRRRRPHNsNCLDRzBmhRa:Q hatR );-
-ApzQazQh1R 7RRRRRRRRRPRRNNsHLRDChe WqRp:)p qR-;
-QAzphaQz71 RRRRRRRRRRRRPHNsNCLDR1pqa _a)Rv:)p qR-;
-QAzphaQz71 RRRRRRRRPHNsNCLDRBwqaRm): R)q:pR=3R4j-;
-QAzphaQz71 
A--zaQpQ1hz R7RRLRRCMoH
A--zaQpQ1hz R7RRRRRRRRRR-R-RlBFbCk0RDPNkVCRF#sRbHCONODRN##C
A--zaQpQ1hz R7RRRRRRVRHR=XRRjj3RC0EM-
-ApzQazQh1R 7RRRRRRRRRRRRRsRRCs0kM3R4j-;
-QAzphaQz71 RRRRRRRRCRM8H
V;-z-AQQpah z17-
-ApzQazQh1R 7RRRRRHRRVXRRpqmBpRR=4R3jRC0EM-
-ApzQazQh1R 7RRRRRRRRRRRRRHRRV R)B)QumpBqRC0EM-
-ApzQazQh1R 7RRRRRRRRRRRRRRRRRRRRRsRRCs0kMqRva4]__ me);_ 
A--zaQpQ1hz R7RRRRRRRRRRRRRRDRC#-C
-QAzphaQz71 RRRRRRRRRRRRRRRRRRRRRRRRskC0svMRq_a] -;
-QAzphaQz71 RRRRRRRRRRRRRRRRCRM8H
V;-z-AQQpah z17RRRRRRRR8CMR;HV
A--zaQpQ1hz -7
-QAzphaQz71 RRRRRRRRHRVRXBpmq=pRRj.3RER0C-M
-QAzphaQz71 RRRRRRRRRRRRRRRRH)VR uBQ)qmBpER0C-M
-QAzphaQz71 RRRRRRRRRRRRRRRRRRRRRRRRskC0s4MR3vj/q_a] ._u;-
-ApzQazQh1R 7RRRRRRRRRRRRRCRRD
#C-z-AQQpah z17RRRRRRRRRRRRRRRRRRRRRRRR0sCkRsMv]qa_u _.-;
-QAzphaQz71 RRRRRRRRRRRRRRRRCRM8H
V;-z-AQQpah z17RRRRRRRR8CMR;HV
A--zaQpQ1hz -7
-QAzphaQz71 RRRRRRRRHRVRXBpmq=pRR34jj0RRE
CM-z-AQQpah z17RRRRRRRRRRRRRRRRRHV)Q BuB)mq0pRE
CM-z-AQQpah z17RRRRRRRRRRRRRRRRRRRRRRRR0sCkRsM4/3jv]qa_u _4
j;-z-AQQpah z17RRRRRRRRRRRRRRRR#CDC-
-ApzQazQh1R 7RRRRRRRRRRRRRRRRRRRRRsRRCs0kMqRva ]__ju4;-
-ApzQazQh1R 7RRRRRRRRRRRRRCRRMH8RV-;
-QAzphaQz71 RRRRRRRRCRM8H
V;-z-AQQpah z17-
-ApzQazQh1R 7RRRRRHRRVpRXmpBqRp>Rm)t5 'qp]]Qt2ER0C-M
-QAzphaQz71 RRRRRRRRRRRRRRRRH)VR uBQ)qmBpER0C-M
-QAzphaQz71 RRRRRRRRRRRRRRRRRRRRRRRRskC0sjMR3
j;-z-AQQpah z17RRRRRRRRRRRRRRRR#CDC-
-ApzQazQh1R 7RRRRRRRRRRRRRRRRRRRRRNRR#s#C0qRwp
1 -z-AQQpah z17RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRbsCFRs0">XRRtpm5q) pQ']tR]2H MRXXu52-"
-QAzphaQz71 RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR#CCPs$H0Rahm -;
-QAzphaQz71 RRRRRRRRRRRRRRRRRRRRRRRRskC0s)MR 'qp]]Qt;-
-ApzQazQh1R 7RRRRRRRRRRRRRCRRMH8RV-;
-QAzphaQz71 RRRRRRRRCRM8H
V;-z-AQQpah z17-
-ApzQazQh1R 7RRRRR-RR-CR)8CkORoNskMlC0FR0R1qA5RX2<3R4j-
-ApzQazQh1R 7RRRRRIRRECHDRmXpBRqp>jR43DjRF
Fb-z-AQQpah z17RRRRRRRRRRRRRRRRmXpBRqp:X=RpqmBpRR-4jj3;-
-ApzQazQh1R 7RRRRRRRRRRRRRwRRqmBa)=R:RBwqa*m)v]qa_u _4
j;-z-AQQpah z17RRRRRRRR8CMRFDFb-;
-QAzphaQz71 
A--zaQpQ1hz R7RRRRRRERIHRDCXBpmq>pRRj43RFDFb-
-ApzQazQh1R 7RRRRRRRRRRRRRXRRpqmBp=R:RmXpBRqp-3R4j-;
-QAzphaQz71 RRRRRRRRRRRRRRRRwaqBm:)R=qRwB)am*avq];_ 
A--zaQpQ1hz R7RRRRRRMRC8FRDF
b;-z-AQQpah z17-
-ApzQazQh1R 7RRRRR-RR-FRBl0bkCNRPDRkCVRFsOCN#R<jRRmXpBRqp<
R4-z-AQQpah z17RRRRRRRR7mpeRqp:4=R3
j;-z-AQQpah z17RRRRRRRR1pqa _a):vR=pRXmpBq;-
-ApzQazQh1R 7RRRRRhRR qWepR:=mep7q+pRR1pqa _a)
v;-z-AQQpah z17RRRRRRRRzBmh:aR=;R.
A--zaQpQ1hz -7
-QAzphaQz71 RRRRRRRR-B-RE	CORsVFRDsCNP0HCMRN8LRN#kFD0CCRsssF#MRN8NRlGFROk
M0-z-AQQpah z17RRRRRRRRHIED5CRR55Rq5A15Wh eRqp-pRm7peq2 /hWpeq2RR> 2u1R
m)-z-AQQpah z17RRRRRRRRRRRRRRRR5RRq5A1he Wq-pRR7mpe2qpR >RuR122hRq7-
-ApzQazQh1R 7RRRRRRRRRRRRRRRRRm5BzRha<qRvXm_BzRha2RR2DbFF
A--zaQpQ1hz R7RRRRRRRRRRRRRRpRm7peqRR:=he Wq
p;-z-AQQpah z17RRRRRRRRRRRRRRRR1pqa _a):vR=qRp1aa_ *)v5mXpBRqp/)R5 5qpBhmza222;-
-ApzQazQh1R 7RRRRRRRRRRRRRhRR qWep=R:R7mpeRqp+qRp1aa_ ;)v
A--zaQpQ1hz R7RRRRRRRRRRRRRRmRBzRha:B=RmazhR4+R;-
-ApzQazQh1R 7RRRRRCRRMD8RF;Fb
A--zaQpQ1hz -7
-QAzphaQz71 RRRRRRRR-B-RFklb0VCRHDMNRDPNkkCR#oHMRbCG5$G+2RR=C5GbGC2*G$b52-
-ApzQazQh1R 7RRRRRhRR qWep=R:RWh e*qpwaqBm
);-z-AQQpah z17-
-ApzQazQh1R 7RRRRRHRRV R)B)QumpBqRC0EM-
-ApzQazQh1R 7RRRRRRRRRRRRRhRR qWep=R:Rj43/Wh e;qp
A--zaQpQ1hz R7RRRRRRMRC8VRH;-
-ApzQazQh1
 7-z-AQQpah z17RRRRRRRR0sCkRsMhe Wq
p;-z-AQQpah z17RRRRMRC8XR u
;

RRRR
--RRRR-q-RkDGHH$NsRMwkOF0HM0#RFFRBl0bkCmRptR
RR-R-
RRRRMVkOF0HMpRQm5tAXH:RM R)qRp2skC0sQMRhta  Q)R1R
RRRRRR-R-R#7CObsH0MHF:R
RRRRRR-R-RRRRRRRR)kC0sRM#MkR#O0ERERN0-<4R=ARq125X/M.^R.<R
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRRMhFCR

RRRRRPRRNNsHLRDChQ:Rhta  :)R=;Rj
RRRRRRRRsPNHDNLC:RYRq) p=R:R1qA5;X2
R
RRCRLo
HMRRRRRRRRHYV5R4=R3FjRsRRY=3Rjj02RE
CMRRRRRRRRRRRRRRRRskC0sjMR;R
RRRRRRMRC8VRH;R

RRRRRHRRVY5RR4>R3Rj20MEC
RRRRRRRRRRRRRRRRHIEDYCRRR>=.R3jDbFF
RRRRRRRRRRRRRRRRRRRRRRRR:YR=/RY.;3j
RRRRRRRRRRRRRRRRRRRRRRRR:hR=+Rh4R;
RRRRRRRRRRRRRCRRMD8RF;Fb
RRRRRRRRRRRRRRRR0sCkRsMhR;
RRRRRCRRMH8RV
;
RRRRRRRR-m-RRY<RR4<R
RRRRRRRRHIEDYCRR4<R3DjRF
FbRRRRRRRRRRRRRRRRY=R:R.Y*3
j;RRRRRRRRRRRRRRRRh=R:R-hR4R;
RRRRRCRRMD8RF;Fb
RRRRRRRR0sCkRsMhR;
RCRRMQ8RpAmt;R

RVRRk0MOHRFMpX7 u:5XRRHM)p q;:RhRRHMQ hat2 )Ra) zR)h)p qR
Q1RRRRRRRR-7-RCs#OHHb0F
M:RRRRRRRR-R-RRRRRRCR)0Mks#*RX.
^MRRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRRMhFCR
RRCRLo
HMRRRRRRRRskC0sXMR*35.j*R*R;h2
RRRR8CMR p7X
u;
A--zaQpQ1hz R7RRkRVMHO0FpMRm5tRXRR:H)MR Rqp2CRs0MksRq) p1RQ
A--zaQpQ1hz R7RRRRRR-R-R#7CObsH0MHF:-
-ApzQazQh1R 7RRRRR-RR-RRRRRRRRC1CRMVkOF0HMCR8OsDNNF0HMMRHR Q  0R18jR4(.n3-g4gn-
-ApzQazQh1R 7RRRRR-RR--
-ApzQazQh1R 7RRRRR-RR-FRh0:C#
A--zaQpQ1hz R7RRRRRR-R-RRRRRRRRN)2RCs0kM)#R 'qppRmWFCMRsssF
A--zaQpQ1hz R7RRRRRR-R-
A--zaQpQ1hz R7RRRRRR-R-RbBF$osHE50RO42RgRg.)CCoMR0#F0VREzCRMCHPs0#H$VRFRDBNHsVFM3HN
A--zaQpQ1hz R7RRRRRR-R-RDqDRosHER0#sCC#s8PC3-
-ApzQazQh1R 7RRRRR-RR--
-ApzQazQh1R 7RRRRR-RR-CR)80H#skHL0MHFR8NMRCk#RRHM#sFkONCRML8RHsMN$FRVs,l#R0IHEsRFR0IHE0Fk
A--zaQpQ1hz R7RRRRRR-R-R8lFHOVHNF0HMN,RsbCRCHsl080CRFbsPCH88ER0N00REVCRFFDDIoHMRMOF8HH0F
M#-z-AQQpah z17RRRRRRRRR--NRsCl:C0
A--zaQpQ1hz R7RRRRRR-R-RR43)HC8#H0sLHk0FRM#F#VRFOksCFRO8lCRkR#0sNC0H0MRENCRLCFPRbOF$osHE-0
-QAzphaQz71 RRRRRRRR-M-RFO0HC0,RERH#D0H#RRFVO8FMHF0HMN#RM08REVCRFFDDIoHMR#8HOHDNl3Cs
A--zaQpQ1hz R7RRRRRR-R-RR.3)HC8#H0sLHk0FRM#HLMRHsMN$FRVsllRkR#0ssCbFO8kCER0CLRNFRPCO$FbsEHo0-
-ApzQazQh1R 7RRRRR-RR-FRM0CHO,ER0HD#RHR#0FOVRFHM80MHF#MRN8ER0CFRVDIDFHRMo8OH#DlNHCHsRMER0C-
-ApzQazQh1R 7RRRRR-RR-FR8OCklM00NHRFMN/M8FFsR0sECR0lNCNsHDb#RsHFP8RC8IEH0RC0ER#8H0LsHkF0HM-3
-QAzphaQz71 RRRRRRRR-d-R3DRqD8RNP0CsHM#HoNRl0HCsNRD#l0CMHHFMMVoRCkN0sRC#FksR#FCRVER0H-#
-QAzphaQz71 RRRRRRRR-#-RFIV0NRsCl0k#R#8Hb$DNRC0ERDVFDHFIMNoROF	MI8DCoCClM
0:-z-AQQpah z17RRRRRRRRR--a#EHRFbs80kOROHMDCk8#FR#VN0Is8CRCDPCF8bCRRL$0RECzPMHCHs#0F$RV-
-ApzQazQh1R 7RRRRR-RR-NRBDFHVsNMH,CRAsD	CCN$RMH8R0O#RFsM0H0LkF3s#
A--zaQpQ1hz R7RRRRRR-R-RRc3h0CHERCs0RECMCNlRRFV0RECzPMHCHs#0M$RF0sREMCRN#lCRRFVH
0#-z-AQQpah z17RRRRRRRRR--O0FMskHL0#FsR$lNRRLCk8#CRR0FCFM8sR#CFbsRsFFl0bCRskF8OR0#8HCsP
C8-z-AQQpah z17RRRRRRRRR--VlsFRH0E#FR#VN0IsICRHF0Ek#0RbHCOVRHObFsHssRIHC00MCRbs#lH#MHF3-
-ApzQazQh1R 7RRRRR-RR--
-ApzQazQh1R 7RRRRR-RR-]RaQ11RmWwaqR) Qu1R)Qme7R 7AaYR]) R ht aq1RhB7Rm)haQaAzmR)1`1`qR'Q1'-
-ApzQazQh1R 7RRRRR-RR-hRq7hRqYXR u1) 1)RmRuQvp7Q R)Wq)aqhQ, 1RBQhpQz7hRt,ARzahRmapQQvaR 7a
m,-z-AQQpah z17RRRRRRRRR--aR] QpvuQR 7W)q)qQha m1Rw Rv)qB]hAaqQapQYhRq7QRwa1h 1mRw)
Rq-z-AQQpah z17RRRRRRRRR--uaq)QpBzqu)Rzm)u1q R)7 RQp1Bq Qv7Q3RhmRhR  eh1aR]pqpR a]Rt)  1haR
m)-z-AQQpah z17RRRRRRRRR--Bamh)zQAa1m)RRA pAQqpw Rmq)Rh7YRQB) aQ,Rh)7Q ,BaRBQhQh7 a,qpR 1uBpQq,-
-ApzQazQh1R 7RRRRR-RR-XR  pvuq,)YRRm)B1mh  TzhqaQpqR7v qt1QR5hzBp7tQh,zRAamRhaQRpv Qa7mRa,-
-ApzQazQh1R 7RRRRR-RR-)Rum)Bz hv awRmRA1z1aaQzRa t7mm1)RmR)1 e QB1p;RmR11mzwR1R ,7qqa,)Rm
A--zaQpQ1hz R7RRRRRR-R-Rmu)w1Qa;)RmR1AzQ1h 1hRQa) )zQuamRh2] mWeR )B1qz q7Rhm7RhhRqY]Ra Ym)
A--zaQpQ1hz R7RRRRRR-R-RRmwpAQqQapQYW,R]] a Q)RhmRBhqa)BRa,1Qa)BpaRQQqApYQa,)RmR)ama-
-ApzQazQh1R 7RRRRR-RR-QR5hzBp7tQhRth p QthRB mm)Ra)] W Q12)RqQh1QthRQRYqhRYWqRamzRRmwa
] -z-AQQpah z17RRRRRRRRR--zR1 mawR]RQ11amwW q),eR  QhRw7Rqe Q17wRmR a]R1um1QQApYQaRRmw1]zB
A--zaQpQ1hz R7RRRRRR-R-Rv7qq3t 
A--zaQpQ1hz R7RRRRRR-R-
A--zaQpQ1hz R7RRRRRR-R-Rahm a:RERH#ep]7RsPC#MHFR#INRMoCC0sNCk8R#oHMRC0ERPBRCHs#FFMRVER0C-
-ApzQazQh1R 7RRRRR-RR-RRRRRRRRsRFHMoHNVDRk0MOHRFML0$REQCR R  ep]7R0vNENCl0NHODNRuOo	NC-
-ApzQazQh1R 7RRRRR-RR-RRRRRRRRFRWsM	HosRtFRkb5/B1K
a2-z-AQQpah z17-
-ApzQazQh1R 7RRRRRORRF0M#NRM0hQ:Rhta  :)R=.R4U-;
-QAzphaQz71 
A--zaQpQ1hz R7RRRRRR-R-RLaNDFCRVFRDo[5w2RR=DwFo_NEC89r[RD+RF_ow0DNHr,[9RsVFRRw[=+R4[./4U-3
-QAzphaQz71 RRRRRRRR-z-R#RC8VRFsoCCMsHN0FFMRVGRC08CMRCbsOHH#FDMRFsoNHl0E#-3
-QAzphaQz71 RRRRRRRR-a-REOCRF0M#NRM0dU64c.d(jUUUdH.R#^R.cR6,#0FRE8CRH8PHC#RHRNCGO
03-z-AQQpah z17RRRRRRRRR--QC0RMs#kCO#RFCssOs0RCHN8MFoRVFRDoEw_C,N8RCCPMFRVsMRHNkOOsCN0
A--zaQpQ1hz R7RRRRRR-R-RO8CHDlN--0FLNHMsO$RFCMPsF#HMFRskM0HCR#35C PsF$L8o$RCR0#0
EC-z-AQQpah z17RRRRRRRRR--sEHo0MRN#sICRsVFRaQh )t #CRD#0#RERNM.d^63-2
-QAzphaQz71 RRRRRRRR-e-RNCDk#FRVsmRpt25wRsICCCRoMNCs0RC8kM#HosRCsRFs<jR4^(-6R#NLF0DkC-
-ApzQazQh1R 7RRRRR-RR-HRI00ERELCRODR-RObN	CNo3-
-ApzQazQh1
 7-z-AQQpah z17RRRRRRRRb0$C R)qep_ mBa)#RHRsNsN5$Rhzqa)RqpsoNMC>R<2VRFRq) p-;
-QAzphaQz71 
A--zaQpQ1hz R7RRRRRRFROMN#0Mq0R4 :)q:pR=3RjjdUdddddddddd(d4U(U.;-
-ApzQazQh1R 7RRRRRORRF0M#NRM0q).: Rqp:j=R3.j46jjjjjjjd4(((.cgd-;
-QAzphaQz71 RRRRRRRRO#FM00NMR:qd)p qRR:=jj3j...d4gdgU4(gg(ccU;jg
A--zaQpQ1hz R7RRRRRRFROMN#0Mq0Rc :)q:pR=3RjjcjjdUcU(((((nj(4(c6c
.;-z-AQQpah z17-
-ApzQazQh1R 7RRRRRORRF0M#NRM0pwmt_Qaqp):R _qpea Bmj)5RRamh:2R=
R5-z-AQQpah z17RRRRRRRRRRRRRRRRjj3,-
-ApzQazQh1R 7RRRRRRRRRRRRR-RRjj3jjjjjjjjjjjjj6.cd.dggUjc.j,cg
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rjjjjjjjjjjjjjj(j4.6(cng(cgn(j4-,
-QAzphaQz71 RRRRRRRRRRRRRRRR-jj3jjjjjjjjjjjj4dd.jU4(4.U.gd.d,-
-ApzQazQh1R 7RRRRRRRRRRRRR-RRjj3jjjjjjjjjj4jj466c..(nUg.UU,(.
A--zaQpQ1hz R7RRRRRRRRRRRRRRjR-3jjjjjjjjjjjjcjjn.n6ggcngd6Uj
j,-z-AQQpah z17RRRRRRRRRRRRRRRRjj3jjjjjjjjjjjj6U4cU6cg(U.n6jU4,-
-ApzQazQh1R 7RRRRRRRRRRRRR-RRjj3jjjjjjjjjj.jj64d.ncUgd(44c,c6
A--zaQpQ1hz R7RRRRRRRRRRRRRRjR-3jjjjjjjjjjjj.j64.dnjgnd46dnj
c,-z-AQQpah z17RRRRRRRRRRRRRRRR3-jjjjjjjjjjjjjj44Ugn6jjjjd4UnU4-,
-QAzphaQz71 RRRRRRRRRRRRRRRRjj3jjjjjjjjjjnjjdj.gn66gUc(.6,cc
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rjjjjjjjjjjjjjj4Unc.64gjdnU4(Uc-,
-QAzphaQz71 RRRRRRRRRRRRRRRR-jj3jjjjjjjjjjjj(6d6(.(j4dgc6Uj.,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3jjjjjjjjjjjjnjgdnUj(Un66.6.(
(,-z-AQQpah z17RRRRRRRRRRRRRRRRjj3jjjjjjjjjjjj(U6gn6dngg(4c44c,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3jjjjjjjjjjjj6j.(ggggU4.dgjng
j,-z-AQQpah z17RRRRRRRRRRRRRRRR3-jjjjjjjjjjjjjj6cncg(.(6c(gcUcc-,
-QAzphaQz71 RRRRRRRRRRRRRRRR-jj3jjjjjjjjjjjj(n66gn.jU6(c4ndd,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3jjjjjjjjjjjj44jgd6(6d..(cjU(
.,-z-AQQpah z17RRRRRRRRRRRRRRRR3-jjjjjjjjjjjjj44(dgcjdccjn.j.dn-,
-QAzphaQz71 RRRRRRRRRRRRRRRR-jj3jjjjjjjjjjjj(U(4jdj4d.nUUUjg,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3jjjjjjjjjjjjg4jU6j(cgjgU.66d
U,-z-AQQpah z17RRRRRRRRRRRRRRRR3-jjjjjjjjjjjjjjc.j(6.d(jUjcgn46-,
-QAzphaQz71 RRRRRRRRRRRRRRRR-jj3jjjjjjjjjjjjU.d(jjg4gdg.6.g4,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3jjjjjjjjjjjjj4cU.U4((gd4444d
6,-z-AQQpah z17RRRRRRRRRRRRRRRRjj3jjjjjjjjj4jj.gUnj44(6U(6U(.6,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3jjjjjjjjjjjj(4(U6UUjU((44gUj
n,-z-AQQpah z17RRRRRRRRRRRRRRRRjj3jjjjjjjjjjjjnjccU46n6gjnn4Ug,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3jjjjjjjjjjjj44nd..U.(nn.Ucj.
.,-z-AQQpah z17RRRRRRRRRRRRRRRR3-jjjjjjjjjjjjjjc(6jng46g446Un4U-,
-QAzphaQz71 RRRRRRRRRRRRRRRR-jj3jjjjjjjjjjjjjnjd64j(UdUU4j(g,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3jjjjjjjjjjjj4jg.djg(g.cgg4cU
c,-z-AQQpah z17RRRRRRRRRRRRRRRRjj3jjjjjjjjj4jjU(6n6g(j6gg(njj4,-
-ApzQazQh1R 7RRRRRRRRRRRRR-RRjj3jjjjjjjjjjdjj4.cgnn6j644gc,Ud
A--zaQpQ1hz R7RRRRRRRRRRRRRRjR-3jjjjjjjjjjjjdjgj6gcg6cg4UgnU
g,-z-AQQpah z17RRRRRRRRRRRRRRRRjj3jjjjjjjjj4jj(cg4dndUj.4dg(44,-
-ApzQazQh1R 7RRRRRRRRRRRRR-RRjj3jjjjjjjjjj4jjdgj.(4g((jddU,nn
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rjjjjjjjjjjjjj.gdj(6dU.64(Udngg-,
-QAzphaQz71 RRRRRRRRRRRRRRRRjj3jjjjjjjjjjdj.g6ggcUjcc4.4(,d(
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rjjjjjjjjjjjjj4g6ddn((4c(c6j6cU-,
-QAzphaQz71 RRRRRRRRRRRRRRRR-jj3jjjjjjjjjdjjnjU(cd.U4d6U(Un(,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3jjjjjjjjjjjjgdn.(jd6.jUjjUjU
g,-z-AQQpah z17RRRRRRRRRRRRRRRR3-jjjjjjjjjjjjjjUgdd(c4.n.dngdng-,
-QAzphaQz71 RRRRRRRRRRRRRRRRjj3jjjjjjjjjjgjjcdddgUU4g.64n,gj
A--zaQpQ1hz R7RRRRRRRRRRRRRR3RjjjjjjjjjjjjjcU4c4Ud4(.jc6nU6U-,
-QAzphaQz71 RRRRRRRRRRRRRRRR-jj3jjjjjjjjjjjjd.(gdc4nUjj.gcd4,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3jjjjjjjjjjjjcjUj6d4ncdj(cg..
c,-z-AQQpah z17RRRRRRRRRRRRRRRR3-jjjjjjjjjjjjjdnc..cgdd.cUU.6cg-,
-QAzphaQz71 RRRRRRRRRRRRRRRRjj3jjjjjjjjjjdjc(44.g64g(gc.4,c6
A--zaQpQ1hz R7RRRRRRRRRRRRRRjR-3jjjjjjjjjjjjc4j(66(jUj6(6(nc
4,-z-AQQpah z17RRRRRRRRRRRRRRRR3-jjjjjjjjjjjjj4444U4n(d6Ug6.gdd-,
-QAzphaQz71 RRRRRRRRRRRRRRRRjj3jjjjjjjjjj(jd66cg(6(.(g.6U,6d
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rjjjjjjjjjjjjj44dg.4Uc.44.gn(66-,
-QAzphaQz71 RRRRRRRRRRRRRRRRjj3jjjjjjjjjjjj4(((6cddj(.6(n,cj
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rjjjjjjjjjjjjj.ggd4gU64nU(cjUjj-,
-QAzphaQz71 RRRRRRRRRRRRRRRR-jj3jjjjjjjjjcjj.j(g6jjgnnjjjc((,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3jjjjjjjjjjjj(..((cjnc44j6dg6
6,-z-AQQpah z17RRRRRRRRRRRRRRRRjj3jjjjjjjjj4jjjgUc6nng.n.g(.g4,-
-ApzQazQh1R 7RRRRRRRRRRRRR-RRjj3jjjjjjjjjjdj.jU(djc4g66(j(,6U
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rjjjjjjjjjjjjj4n6(4d.j(g(dndgc6-,
-QAzphaQz71 RRRRRRRRRRRRRRRRjj3jjjjjjjjjjdjjd(c64nj.gc6cj,U.
A--zaQpQ1hz R7RRRRRRRRRRRRRRjR-3jjjjjjjjjjjj6c4.664Udjnc4dn.
d,-z-AQQpah z17RRRRRRRRRRRRRRRRjj3jjjjjjjjjdjj.6n6nUgUgjng(n4c,-
-ApzQazQh1R 7RRRRRRRRRRRRR-RRjj3jjjjjjjjjjcjc(.jcn46jj.c6c,cn
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rjjjjjjjjjjjjjd.c6((ncgj6.d(g(.-,
-QAzphaQz71 RRRRRRRRRRRRRRRR-jj3jjjjjjjjjjjj(Ujcgdn.gj.4gn(c,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3jjjjjjjjjjjj(44((ngU4(6d.ng4
c,-z-AQQpah z17RRRRRRRRRRRRRRRR3-jjjjjjjjjjjjj4(j(c4dccnn4j(g6U-,
-QAzphaQz71 RRRRRRRRRRRRRRRRjj3jjjjjjjjjj4j.Udndcgd.d6.4g,4j
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rjjjjjjjjjjjjj.dc4.gndcdg4ddd44-,
-QAzphaQz71 RRRRRRRRRRRRRRRRjj3jjjjjjjjjjgjdjc6(nj..gjUd(,jj
A--zaQpQ1hz R7RRRRRRRRRRRRRRjR-3jjjjjjjjjjjj6.n((jngd.j6(nj6
4,-z-AQQpah z17RRRRRRRRRRRRRRRRjj3jjjjjjjjjdjj(64d4gc44gg6.4j.,-
-ApzQazQh1R 7RRRRRRRRRRRRR-RRjj3jjjjjjjjjj(j44gnn.d4dn.jUc,d4
A--zaQpQ1hz R7RRRRRRRRRRRRRRjR-3jjjjjjjjjjjjn.U6UU.6(46gd4c6
d,-z-AQQpah z17RRRRRRRRRRRRRRRR3-jjjjjjjjjjjjj.4dU..6c.cndcjnUg-,
-QAzphaQz71 RRRRRRRRRRRRRRRRjj3jjjjjjjjjjnjj6n(n6ng(Uj6Uj,n.
A--zaQpQ1hz R7RRRRRRRRRRRRRRjR-3jjjjjjjjjjjj..U4cj4dnUc4.U4n
(,-z-AQQpah z17RRRRRRRRRRRRRRRRjj3jjjjjjjjj4jjj4(jg(d4n4.4cc.6,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3jjjjjjjjjjjj44U4cgdnndnc4c44
j,-z-AQQpah z17RRRRRRRRRRRRRRRRjj3jjjjjjjjjjjjgjUcc.n6(dU..(n.,-
-ApzQazQh1R 7RRRRRRRRRRRRR-RRjj3jjjjjjjjjjdjd44cg6Uj...(66,c.
A--zaQpQ1hz R7RRRRRRRRRRRRRRjR-3jjjjjjjjjjjjd4Uj6.U(nd6jnc4n
U,-z-AQQpah z17RRRRRRRRRRRRRRRR3-jjjjjjjjjjjjj4jn.(jcj4(6ncccgg-,
-QAzphaQz71 RRRRRRRRRRRRRRRRjj3jjjjjjjjjjUjcddjd4ccggd66.,j4
A--zaQpQ1hz R7RRRRRRRRRRRRRRjR-3jjjjjjjjjjjj6(4n6j6d.4(d4U.4
6,-z-AQQpah z17RRRRRRRRRRRRRRRRjj3jjjjjjjjjUjjU4U..6dg4(U646U6,-
-ApzQazQh1R 7RRRRRRRRRRRRR-RRjj3jjjjjjjjjjjjdg6jjU4j6dU.d.,cc
A--zaQpQ1hz R7RRRRRRRRRRRRRRjR-3jjjjjjjjjjjjjn4(6n64.g(Uc64g
n,-z-AQQpah z17RRRRRRRRRRRRRRRRjj3jjjjjjjjjdjj6gn6gnngncdd(jUd,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3jjjjjjjjjjjj(d6Ug.dn46g.d(nU
d,-z-AQQpah z17RRRRRRRRRRRRRRRR3-jjjjjjjjjjjjjc.n.n(jUj6j4c(c6U-,
-QAzphaQz71 RRRRRRRRRRRRRRRRjj3jjjjjjjjjj.jn.((gn4.g(6..4,6n
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rjjjjjjjjjjjjj(d.UU(gc.j(.nc6(4-,
-QAzphaQz71 RRRRRRRRRRRRRRRRjj3jjjjjjjjjjnj.Unjgc4nn64.4n,(d
A--zaQpQ1hz R7RRRRRRRRRRRRRRjR-3jjjjjjjjjjjjg4jn.jU6njcj.6g(
U,-z-AQQpah z17RRRRRRRRRRRRRRRRjj3jjjjjjjjjjjj.4d4gdcgUjdUj(6d,-
-ApzQazQh1R 7RRRRRRRRRRRRR-RRjj3jjjjjjjjjjUj6cjng6jUj6g.g.,c(
A--zaQpQ1hz R7RRRRRRRRRRRRRRjR-3jjjjjjjjjjjj4j.jcd(U4.64cccg
c,-z-AQQpah z17RRRRRRRRRRRRRRRR3-jjjjjjjjjjjjj..ddd.4Ug6c6Uj(cU-,
-QAzphaQz71 RRRRRRRRRRRRRRRR-jj3jjjjjjjjjcjj.dddn.gcUcU44ng4,-
-ApzQazQh1R 7RRRRRRRRRRRRR-RRjj3jjjjjjjjjjdjcggdddn(gg((dU,cc
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rjjjjjjjjjjjjjcc4d4(ncjU(ddn666-,
-QAzphaQz71 RRRRRRRRRRRRRRRRjj3jjjjjjjjjjnjjU(c4ncdn446gc,nn
A--zaQpQ1hz R7RRRRRRRRRRRRRR3RjjjjjjjjjjjjjcU(66c6djcjcdcjn4-,
-QAzphaQz71 RRRRRRRRRRRRRRRRjj3jjjjjjjjjjdjUnn(g((Unc((6n,g6
A--zaQpQ1hz R7RRRRRRRRRRRRRRjR-3jjjjjjjjjjjj(U6ndd(cnncnn6Uc
j,-z-AQQpah z17RRRRRRRRRRRRRRRRjj3jjjjjjjjj.jj4dg4..U4.cgdj.jg,-
-ApzQazQh1R 7RRRRRRRRRRRRR-RRjj3jjjjjjjjjj.jn.Uc.cd.6n4cd4,cU
A--zaQpQ1hz R7RRRRRRRRRRRRRRjR-3jjjjjjjjjjjjg4jUgd6c6d.ccdUd
j,-z-AQQpah z17RRRRRRRRRRRRRRRRjj3jjjjjjjjjnjj6jd4cdd4(d(nd4n6,-
-ApzQazQh1R 7RRRRRRRRRRRRR-RRjj3jjjjjjjjjj(jc64Ujg.gj4j(4(,ng
A--zaQpQ1hz R7RRRRRRRRRRRRRRjR-3jjjjjjjjjjjjUd(66c.46.ncj6(c
j,-z-AQQpah z17RRRRRRRRRRRRRRRRjj3jjjjjjjjjcjjjggd..dd4(UnUcnn,-
-ApzQazQh1R 7RRRRRRRRRRRRRjRR3jjjjjjjjjjjjcU(.Ucddcg4U.6Ug
4,-z-AQQpah z17RRRRRRRRRRRRRRRRjj3jjjjjjjjj.jj6U.44cUU6cnU..UU,-
-ApzQazQh1R 7RRRRRRRRRRRRR-RRjj3jjjjjjjjjjdjjn4jUdn4dj.c.6,6(
A--zaQpQ1hz R7RRRRRRRRRRRRRRjR-3jjjjjjjjjjjj66j46U66cg..gUjj
.,-z-AQQpah z17RRRRRRRRRRRRRRRRjj3jjjjjjjjj(jjUgngcdjd.6dd6(d4,-
-ApzQazQh1R 7RRRRRRRRRRRRR-RRjj3jjjjjjjjjj(jnjU.j(nng4ggcj,nj
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rjjjjjjjjjjjjj4jn4U66((g6dd6.cU-,
-QAzphaQz71 RRRRRRRRRRRRRRRRjj3jjjjjjjjjjUj664.(UdUcn4.66,jg
A--zaQpQ1hz R7RRRRRRRRRRRRRRjR-3jjjjjjjjjjjj.d6c6n(((.gg(jcg
4,-z-AQQpah z17RRRRRRRRRRRRRRRR3-jjjjjjjjjjjjj4(Ud.cjUcng6.6gjU-,
-QAzphaQz71 RRRRRRRRRRRRRRRRjj3jjjjjjjjjjUjUnnjnU4gUdccgg,4n
A--zaQpQ1hz R7RRRRRRRRRRRRRR3RjjjjjjjjjjjjjnUncnU.njc(4njU(j-,
-QAzphaQz71 RRRRRRRRRRRRRRRRjj3jjjjjjjjjjdjnUnd44(64jnnc6,4g
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rjjjjjjjjjjjjj.c64cj.d(d.U((nj.-,
-QAzphaQz71 RRRRRRRRRRRRRRRR-jj3jjjjjjjjj4jj(g.dc6cc.46nccUd2-;
-QAzphaQz71 
A--zaQpQ1hz R7RRRRRRFROMN#0Mp0Rm_tw]7 q: R)qep_ mBa)R5jahmR2=R:R-5
-QAzphaQz71 RRRRRRRRRRRRRRRRj,3j
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rjj(j(Uc.4j.ccjdnjUc4.n-,
-QAzphaQz71 RRRRRRRRRRRRRRRRj43j6c6j46Undn6gdn6.n,gc
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rjj4.dn6(jg4.U6nc(jjUcn-,
-QAzphaQz71 RRRRRRRRRRRRRRRRjd3jj4((nn6Unnn(6d.dn,c(
A--zaQpQ1hz R7RRRRRRRRRRRRRR3RjjddU4nUUc.dj4.c4nUccU-,
-QAzphaQz71 RRRRRRRRRRRRRRRRjc3j6gUj6jdndc4..c(4n,(j
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rjj.6dc4c6cU64Und(j6c66-,
-QAzphaQz71 RRRRRRRRRRRRRRRRjn3jjcn.nU.44UncnUg((,Un
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rjjgn(6njn4Ugj6g.6c6ccc-,
-QAzphaQz71 RRRRRRRRRRRRRRRRj(3j6d..c..4d.(6c6.dj,dg
A--zaQpQ1hz R7RRRRRRRRRRRRRR3RjjcU.cndngj.4gcUUcdn4U-,
-QAzphaQz71 RRRRRRRRRRRRRRRRjU3jg.n44n6UUng(jjngd,..
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rjj(gn..gnnUc6c(6cd44nU-,
-QAzphaQz71 RRRRRRRRRRRRRRRRjj34dn(g(ngdUn46(U6(c,nj
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rj4U4j4ncdnjdc.dnc4jc.d-,
-QAzphaQz71 RRRRRRRRRRRRRRRRj434(d(Ujnd66dncj4jjU,dn
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rj4(.cj(dcU46jjUd.j(6jj-,
-QAzphaQz71 RRRRRRRRRRRRRRRRjd344n6(d(6(U4Un(6d4.,dn
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rj4cdUj..d.gU6.dg...njg-,
-QAzphaQz71 RRRRRRRRRRRRRRRRjc346.4UjUjgc(c66(j(.,g6
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rj4g644cnj.6j.(4d.nd(6j-,
-QAzphaQz71 RRRRRRRRRRRRRRRRj634U6njj4dj(6nngnj6c,64
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rj4.n6c(g6.6UgdUgjUUd(n-,
-QAzphaQz71 RRRRRRRRRRRRRRRRj(344jU6.g6n.4n6U4dcj,nj
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rj4c(Uj6(n(.c(nnUgjcng(-,
-QAzphaQz71 RRRRRRRRRRRRRRRRjU34c.g.dcdUgddUcc4j4,6n
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rj4dg4g6cU.ggg6jn6ccnj(-,
-QAzphaQz71 RRRRRRRRRRRRRRRRjg34(6U.(dcd.6g(U.664,d6
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rj..jc4c664Uc.(dnnjnjnU-,
-QAzphaQz71 RRRRRRRRRRRRRRRRj43.jc6n(4ngj6(dj.jj(,c4
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rj.U4n(ddgUjdj64.d6cj.n-,
-QAzphaQz71 RRRRRRRRRRRRRRRRj.3.dd4c6d644.cjcjjUj,6n
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rj.d.g(jc44cjnUd((.c.n.-,
-QAzphaQz71 RRRRRRRRRRRRRRRRjd3.6n6njd(44n.Ujdjjn,(.
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rj.(c44dggnnUUgjnn.6c(U-,
-QAzphaQz71 RRRRRRRRRRRRRRRRjc3.(nUd4gndjgc6cn.U6,((
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rj.g6d4j6.gjgU(cd.(Uj.6-,
-QAzphaQz71 RRRRRRRRRRRRRRRRj63.g(g66c.cdUnnn4j(6,n(
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rj.gn6ncd6UncggjUcj(d6(-,
-QAzphaQz71 RRRRRRRRRRRRRRRRj(3.4dgd(c46U4cjjdcn4,4c
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rj.U((n6Uc4djjj4U(jd.c6-,
-QAzphaQz71 RRRRRRRRRRRRRRRRjU3.dU(n44(dddj(U.cd6,4g
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rj.nUgdgd...6UgdcUcg.Un-,
-QAzphaQz71 RRRRRRRRRRRRRRRRjg3.6ccn.U4.g.dc4djn4,gg
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rjd.j4nd4djU6(4(ggj(c4(-,
-QAzphaQz71 RRRRRRRRRRRRRRRRjj3d(6j.j.d6g.cU(jUd6,4.
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rjd(4.646(jcjj.6dg4.((g-,
-QAzphaQz71 RRRRRRRRRRRRRRRRj43dUdc6(4d44gUj(dcgU,gj
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rjd4.c4ngcUcn6d(4ndgd64-,
-QAzphaQz71 RRRRRRRRRRRRRRRRj.3dgd(6.dUn((.6gU4n6,.U
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rjddd66c664jg.(dn.dUccc-,
-QAzphaQz71 RRRRRRRRRRRRRRRRjc3djng.6gUn(6jcc4jUU,g.
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rjdccnnnn((ndc4Ujj.UdcU-,
-QAzphaQz71 RRRRRRRRRRRRRRRRj63d4ng(c4.d6UnUcn.nj,nd
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rjdc6(6U6UU.g..nd4(4gdn-,
-QAzphaQz71 RRRRRRRRRRRRRRRRjn3d.6gjcngdUcg4j.(4d,(n
A--zaQpQ1hz R7RRRRRRRRRRRRRR3RjddnU.n664U4664gg66(d.-,
-QAzphaQz71 RRRRRRRRRRRRRRRRj(3ddn(4c(jgg4dUcUU4U,cj
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rjdj(g(6Ud.cgdUU44c6ndd-,
-QAzphaQz71 RRRRRRRRRRRRRRRRjU3dc4c4nggU4gj.U.6Un,d.
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rjd(Ug46n(4j4ccccjn6cg4-,
-QAzphaQz71 RRRRRRRRRRRRRRRRjg3dcdggU.jUccj6.4c.4,4(
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rjc.jjcnd4c(4.c(6gc(g6g-,
-QAzphaQz71 RRRRRRRRRRRRRRRRjj3c66cn44jUj4(Ug64jc,gU
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rjcn4j6.ggc6gUdUdU(666U-,
-QAzphaQz71 RRRRRRRRRRRRRRRRj43c6(U.U4g6cgd6d64gU,.6
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rjcg.jngg.ccnc.dd((cg6d-,
-QAzphaQz71 RRRRRRRRRRRRRRRRj.3cncjUddg64Ujn4gc.n,g4
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rjc4d4(ndccUU44jdj4nccc-,
-QAzphaQz71 RRRRRRRRRRRRRRRRjd3cnn.d((nn(.c6(6cg(,.n
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rjc.c4(nc6j6Uj4gcjdUn.4-,
-QAzphaQz71 RRRRRRRRRRRRRRRRjc3cn(.U4nj..cUjUj4n4,4d
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rjc.64(ccncg4dn.dj66cdU-,
-QAzphaQz71 RRRRRRRRRRRRRRRRj63cn(.dccddU(4Uc(4(.,d.
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rjc4n4(46(6.4.c.jUgg4(j-,
-QAzphaQz71 RRRRRRRRRRRRRRRRjn3cngjU(g.g.dc6d(c6g,nj
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rjcg(j(4g(6g.4j4(d4Udg6-,
-QAzphaQz71 RRRRRRRRRRRRRRRRj(3c66UcgUjcn6gUncUgg,c(
A--zaQpQ1hz R7RRRRRRRRRRRRRR3RjcnUjU.U6g6dc6((j44c..-,
-QAzphaQz71 RRRRRRRRRRRRRRRRjU3c6(6jU(46Uj4n.dcj4,cg
A--zaQpQ1hz R7RRRRRRRRRRRRRR3RjcdgjjUdgU6jc6d.6.6gnd-,
-QAzphaQz71 RRRRRRRRRRRRRRRRjg3c6(j(.(nngdUjcd6c4,(4
A--zaQpQ1hz R7RRRRRRRRRRRRRR3RjcUgg.n(Ugn66nc44j.dU.-,
-QAzphaQz71 RRRRRRRRRRRRRRRRjj36cn66j(4j644g.d.6g,jU
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rj6.jgnj4g4j(g66.d6d.d6-,
-QAzphaQz71 RRRRRRRRRRRRRRRRj436d6gc(464jc4dnc4jc,j6
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rj6n4Ujn((cU.jdn6cd6(gU-,
-QAzphaQz71 RRRRRRRRRRRRRRRRj.36dU.c4(cdn664U.njj,dn
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rj6U.(nU(jgjn.c(U6U46c(-,
-QAzphaQz71 RRRRRRRRRRRRRRRRjd36.ccn(UgUn4g4cgj4g,jU
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rj6jd(cn4c6(Ugdgc64d6cn-,
-QAzphaQz71 RRRRRRRRRRRRRRRRjc364(6g.cU.d..44d6(g,c(
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rj64cndd.c((6gc.j(njjgg-,
-QAzphaQz71 RRRRRRRRRRRRRRRRj636j(nc4g4(6g.dc.4U(,gd
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rj6466cj46(j6cn.44jnjg6-,
-QAzphaQz71 RRRRRRRRRRRRRRRRj636g6n4(gU(dg6dgn6n(,((
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rj6jnc(dj4U6.UdnU(66nn4-,
-QAzphaQz71 RRRRRRRRRRRRRRRRjn36Uc6j(dd66U.ngg(c6,n4
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rj6g(.46g(d.6nj(4Uc.jg.-,
-QAzphaQz71 RRRRRRRRRRRRRRRRj(36(6d4djn6dc6.n4gc.,nj
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rj6nU4gd4(g6ndjUn4.j4gj-,
-QAzphaQz71 RRRRRRRRRRRRRRRRjU36ngjcjjc6jnd4c.(gc,dd
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rj6dgjUc(cn.nj4gj(6j(j6-,
-QAzphaQz71 RRRRRRRRRRRRRRRRjg36c((j4(j(c4n.ncgd4,(c
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rj6jggjUU4g6nc.ncnjg.6c-,
-QAzphaQz71 RRRRRRRRRRRRRRRRjj3ndj.gUc64dcUg4gUgn,U(
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rjn6j(666.jc..dn..nU.nU-,
-QAzphaQz71 RRRRRRRRRRRRRRRRj43n44Uj64c4j4nn64ddg,66
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rjnj4n.(gU(6.4nU.d6g66j-,
-QAzphaQz71 RRRRRRRRRRRRRRRRj.3njj.cc(jg6j4.ccc.6,d(
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rjnc.cdUd.U.j4ddngjddj.-,
-QAzphaQz71 RRRRRRRRRRRRRRRRj.3nUUnjnc6g.6.(.jnU.,6n
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rjn(d.nnnngj6(nc.Ud4(.d-,
-QAzphaQz71 RRRRRRRRRRRRRRRRjd3nn(gjc.n.dgn4c(gU(,U4
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rjnjc4d(44gjc.n4(gj(g44-,
-QAzphaQz71 RRRRRRRRRRRRRRRRjc3n6(4dgdn4(.dnj.(Ug,(U
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rjn.cg.c(gn6n.nj46j6ccj-,
-QAzphaQz71 RRRRRRRRRRRRRRRRj63nd4dj.j(.464gUcnc(,.6
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rjnd6(6(Uj.g(jj.djd4Ug4-,
-QAzphaQz71 RRRRRRRRRRRRRRRRjn3n4Udgc.U.cj6.d.g.6,j.
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rjncn6.d.n.c6c64j6(n(j6-,
-QAzphaQz71 RRRRRRRRRRRRRRRRjn3ngjcdng6dcU.g4c(dU,(4
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rjnc(d.(.n6..4dc6jcc44.-,
-QAzphaQz71 RRRRRRRRRRRRRRRRj(3n(UdgU6.dg.jgjdj(g,44
A--zaQpQ1hz R7RRRRRRRRRRRRRR3RjndU46.g.c(Uj..dUjnn.(-,
-QAzphaQz71 RRRRRRRRRRRRRRRRjU3n6cdjjjjdgUU.4j4jd,g.
A--zaQpQ1hz R7RRRRRRRRRRRRRR3Rjn.UgdUd.4U.d666(d4Uj(-,
-QAzphaQz71 RRRRRRRRRRRRRRRRjg3nd(4c46Ujn4j4(d(jU2n.;-
-ApzQazQh1
 7-z-AQQpah z17RRRRRRRRsPNHDNLC,RvRQK:hta  
);-z-AQQpah z17RRRRRRRRsPNHDNLC4Rw,.Rw,,RtRRT,zz,R.e,R: R)q
p;-z-AQQpah z17RRRRRRRRsPNHDNLC RZ)Rm:)p qRR:=j;3j-N-v8PCRNNsHLRDC#MFRFFROMN#0MV0RFHD8MFoROsOk#-
-ApzQazQh1R 7RRRRRPRRNNsHLRDCm:h Rq) p=R:Rj43;-R-vCN8RsPNHDNLCFR#RRMFO#FM00NMRDVF8oHMROFOk
s#-z-AQQpah z17-
-ApzQazQh1R 7RRRRR-RR-FR8kCLDRoDFL,52RCD8G2b5;-
-ApzQazQh1
 7-z-AQQpah z17RRRRRRRRsPNHDNLC4Rz:q) p-;
-QAzphaQz71 
A--zaQpQ1hz R7RRLRRCMoH
A--zaQpQ1hz -7
-QAzphaQz71 RRRRRRRR-B-RE	CORDPNH08H$VRFRoNskMlC0-
-ApzQazQh1R 7RRRRRHRRVRR5X=R<Rjj3R02RE
CM-z-AQQpah z17#--$EM0C##HRN0sMN#D0FC_V-V
-QAzphaQz71 RRRRRRRRRRRRRRRRNC##sw0Rq p1
A--zaQpQ1hz R7RRRRRRRRRRRRRRRRRRRRRRCRsb0FsRR"X<j=R3HjRMmRpt25X"-
-ApzQazQh1R 7RRRRRRRRRRRRRRRRRRRRR#RRCsPCHR0$ m)))-;
-QAzphaQz71 -$-#MC0E#RH#0MsN#0DNCM_F
A--zaQpQ1hz R7RRRRRRRRRRRRRRCRs0Mks5q) pm'pW
2;-z-AQQpah z17RRRRRRRR8CMR;HV
A--zaQpQ1hz -7
-QAzphaQz71 RRRRRRRR-B-RFklb0PCRNCDkRsVFRC#bODHNR#ONC-#
-QAzphaQz71 RRRRRRRRH5VRR=XRRj43R02RE
CM-z-AQQpah z17RRRRRRRRRRRRRRRR0sCkRsMj;3j
A--zaQpQ1hz R7RRRRRRMRC8VRH;-
-ApzQazQh1
 7-z-AQQpah z17RRRRRRRRRHV5RRX=qRva ]_R02RE
CM-z-AQQpah z17RRRRRRRRRRRRRRRR0sCkRsM4;3j
A--zaQpQ1hz R7RRRRRRMRC8VRH;-
-ApzQazQh1
 7-z-AQQpah z17RRRRRRRRR--qksol0CMR8sCkHO0FRM:4=R<R<oRRR.;G^/.lRR=o-;
-QAzphaQz71 RRRRRRRR-$-RRw=R*R54+/RVwV2RF|sRV<|R=^R.--U
-QAzphaQz71 
A--zaQpQ1hz R7RRRRRRRRv:Q=RpAmt5;X2
A--zaQpQ1hz R7RRRRRRRRt:p=R7u X5RX,-;v2
A--zaQpQ1hz R7RRRRRRRRK:Q=Rhta  ))5 5qph52*t3-4j;22RR--BFRO8NCR8R8#jR36VRFssMFk8oHM
A--zaQpQ1hz R7RRRRRR4RwRR:=5j43/q) p25h2RR*)p q5RK2+3R4j-;R-*w44R.UHN#RMhRQa  t)MRHR.r4U4,6.-9
-QAzphaQz71 RRRRRRRRw:.R=RRt-4Rw;-
-ApzQazQh1
 7-z-AQQpah z17RRRRRRRRR--qsbbFlGHNR0CCNGbMF#HMFRVsFRDo+54Vw./4~2R=RRk+
RJ-z-AQQpah z17RRRRRRRR:tR=3R4j./53wj*4.+w2-;
-QAzphaQz71 RRRRRRRRz=R:Rj.3**w.t-;
-QAzphaQz71 RRRRRRRRe=R:Rzz*;-
-ApzQazQh1R 7RRRRRTRRRR:=z**e5Rq4+*Re5Rq.+*Re5Rqd+*Req2c22-;
-QAzphaQz71 
A--zaQpQ1hz R7RRRRRR-R-R#BNC:R4RRk4=RRksMFk8RC80.FR^d-cR#NLF0DkC13RHCMOR<kRR-.^U-,
-QAzphaQz71 RRRRRRRR-R-RRRRRRRk4ERN#Nl0RFR#0dL6RH,0#R8NMR*w4kH4R#GRCN,O0RRN#wE4RN<#RRLURH30#
A--zaQpQ1hz R7RRRRRR-R-RRRRRQRR0DRN#NFR8R8#COGN0RD$0|FRlF*DoE._HRR+D_FowC_EN[8r9RR|<6R(j-3
-QAzphaQz71 RRRRRRRR---
-QAzphaQz71 RRRRRRRRH5VRR/KR=RRjFvsRRR/=j02RE
CM-z-AQQpah z17RRRRRRRRRRRRRRRRRz4:z=RR6+R4jd3;-
-ApzQazQh1R 7RRRRRRRRRRRRRzRR4=R:RRz4-4R6d;3j
A--zaQpQ1hz -7
-QAzphaQz71 RRRRRRRRRRRRRRRR-B-RNR#C.|:R4|-GR4<R/n.63ERaC-RlR8NMRR[-8CCbMM8C0CR0sRl#NRsCxFCs
A--zaQpQ1hz R7RRRRRRRRRRRRRR-R-RRRRRRRRk=4RR0kRFcR.R0LH#-3
-QAzphaQz71 RRRRRRRRRRRRRRRR---
-QAzphaQz71 RRRRRRRRCCD#
A--zaQpQ1hz R7RRRRRRRRRRRRRR4RzRR:=z-;
-QAzphaQz71 RRRRRRRRRRRRRRRR-)-az5hBz;42RQ--MRRO0#EHRRH#k=4RRF58kCLD2VR5D0FN2kR54-2
-QAzphaQz71 RRRRRRRRCRM8H
V;-z-AQQpah z17-
-ApzQazQh1R 7RRRRRzRR.=R:R35.jw*5.RR-wz4*4-2RR*z4wR.2*;Rt
A--zaQpQ1hz R7RRRRRR-R-RRk4+.RkR.=RV./5w2+VRR0FCsG0NsRbC#OHH3FM
A--zaQpQ1hz -7
-QAzphaQz71 RRRRRRRR-D-RFGo52RR=D5Fo.*^lw54*4.+V/2w42
R=-z-AQQpah z17RRRRRRRRR--5Dl*F_o.EpH+m_tw]7 q5+[2kR42+lR5*oDF.F_D+tpmwq_aQ[p522+J;-
-ApzQazQh1R 7RRRRR-RR-CR5G0NO2RR+5M0H$-2
-QAzphaQz71 
A--zaQpQ1hz R7RRRRRR4RzRR:=z+4RRq) p25v*tpmw _]qh752RR+pwmt_q] 725K;RRRRRRRRR-- OGN0-
-ApzQazQh1R 7RRRRRzRR.=R:R.5zRp+Rm_twapqQ52K2RT+R;RRRRRRRRR--a$HM
A--zaQpQ1hz R7RRRRRR.RzRR:=z+.RRtpmwq_aQhp52 *)qvp52-;
-QAzphaQz71 RRRRRRRRskC0s5MRz+4RR2z.;-
-ApzQazQh1R 7RCRRMp8Rm
t;
R
RRkRVMHO0FpMRmRt.5RX:H)MR 2qpR0sCkRsM)p qR
H#RRRRRRRR-7-RCs#OHHb0F
M:RRRRRRRR-R-RRRRRRCR1CkRVMHO0F8MRCNODsHN0FHMRM RQ 1 R048Rj3(n.g-4gRn
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRNRR2CR)0Mks# R)qpp'mFWRMsRCs
FsRRRRLHCoMR
RRRRRR-R-RCBEOP	RN8DHHR0$FNVRslokC#M0
RRRRRRRRRHV5RRX<j=R32jRRER0C-M
-M#$0#ECH0#Rs#NMDCN0_VFV
RRRRRRRRRRRRRRRR#N#CRs0w1qp R
RRRRRRRRRRRRRRRRRRRRRRCRsb0FsRR"X<j=R3HjRMmRptX.52R"
RRRRRRRRRRRRRRRRRRRRR#RRCsPCHR0$ m)))-;
-M#$0#ECH0#Rs#NMDCN0_
FMRRRRRRRRRRRRRRRRskC0s)M5 'qpp2mW;R
RRRRRRMRC8VRH;R

RRRRR-RR-FRBl0bkCNRPDRkCVRFs#ObCHRNDOCN##R
RRRRRRVRHRX5RR4=R32jRRC0EMR
RRRRRRRRRRRRRRCRs0MksRjj3;R
RRRRRRMRC8VRH;R

RRRRRHRRVRR5XRR=.R3j2ER0CRM
RRRRRRRRRRRRRsRRCs0kM3R4jR;
RRRRRCRRMH8RV
;
RRRRRRRR-B-RFklb0PCRNCDkRsVFRMoCCDsNR#ONCR
RRRRRRCRs0MksRv5Rq_a]p.mt__mw m*pt25XR
2;RRRRCRM8p.mt;


RRRRVOkM0MHFRtpm45jRXH:RM R)qRp2skC0s)MR RqpHR#
RRRRR-RR-CR7#HOsbF0HMR:
RRRRR-RR-RRRRRRRRC1CRMVkOF0HMCR8OsDNNF0HMMRHR Q  0R18jR4(.n3-g4gnR
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRR2RNR0)Ck#sMRq) pm'pWMRFRsCsFRs
RLRRCMoH
RRRRRRRRR--BOEC	NRPDHH80F$RVsRNoCklM
0#RRRRRRRRH5VRR<XR=3RjjRR2RC0EM-
-#0$MEHC##sR0NDM#N_0CF
VVRRRRRRRRRRRRRRRRRNRR#s#C0qRwp
1 RRRRRRRRRRRRRRRRRRRRRRRRsFCbs"0RX=R<Rjj3RRHMp4mtj25X"R
RRRRRRRRRRRRRRRRRRRRRRCR#PHCs0 $R)))m;-
-#0$MEHC##sR0NDM#N_0CFRM
RRRRRRRRRRRRRRRRRCRs0Mks5q) pm'pW
2;RRRRRRRRCRM8H
V;
RRRRRRRRR--BbFlkR0CPkNDCFRVsbR#CNOHDNRO#
C#RRRRRRRRH5VRR=XRRj43R02RE
CMRRRRRRRRRRRRRRRRskC0sjMR3
j;RRRRRRRRCRM8H
V;
RRRRRRRRRHV5RRX=jR432jRRC0EMR
RRRRRRRRRRRRRRCRs0MksRj43;R
RRRRRRMRC8VRH;R

RRRRR-RR-FRBl0bkCNRPDRkCVRFsoCCMsRNDOCN#
RRRRRRRR0sCkRsM5qRvap]_mjt4__mw m*pt25XR
2;RRRRCRM8p4mtj
;

RRRRMVkOF0HMmRptXR5:MRHRq) pA;Rq:1 RRHM)p q2CRs0MksRq) p#RH
RRRRRRRRR--7OC#s0HbH:FM
RRRRRRRRR--RRRRR1RRCVCRk0MOHRFM8DCON0sNHRFMHQMR R  1R084nj(34.-g
gnRRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRN)2RCs0kM)#R 'qppRmWFCMRsssF
RRRRoLCHRM
RRRRR-RR-ERBCRO	PHND8$H0RRFVNksol0CM#R
RRRRRRVRHRX5RRR<=jR3j20RRE
CM-$-#MC0E#RH#0MsN#0DNCV_FVR
RRRRRRRRRRRRRRNRR#s#C0qRwp
1 RRRRRRRRRRRRRRRRRRRRRRRRsFCbs"0RX=R<Rjj3RRHMp5mtXA,Rq21 "R
RRRRRRRRRRRRRRRRRRRRRRCR#PHCs0 $R)))m;-
-#0$MEHC##sR0NDM#N_0CFRM
RRRRRRRRRRRRRRRRskC0s)M5 'qpp2mW;R
RRRRRRMRC8VRH;R

RRRRRHRRVRR5A q1RR<=jR3jFAsRqR1 =3R4jRR2RC0EMR
RRRRRRRRRRRRRRNRR#s#C0qRwp
1 RRRRRRRRRRRRRRRRRRRRRRRRsFCbs"0RA q1RR<=jR3jFAsRqR1 =3R4jMRHRtpm5RX,A q12R"
RRRRRRRRRRRRRRRRRRRRR#RRCsPCHR0$ m)))R;
RRRRRRRRRRRRRRRRskC0s)M5 'qpp2mW;R
RRRRRRMRC8VRH;R

RRRRR-RR-FRBl0bkCNRPDRkCVRFs#ObCHRNDOCN##R
RRRRRRVRHRX5RR4=R32jRRC0EMR
RRRRRRRRRRRRRRCRs0MksRjj3;R
RRRRRRMRC8VRH;R

RRRRRHRRVRR5XRR=A q1R02RE
CMRRRRRRRRRRRRRRRRskC0s4MR3
j;RRRRRRRRCRM8H
V;
RRRRRRRRR--BbFlkR0CPkNDCFRVsCRoMNCsDNRO#RC
RRRRRsRRCs0kMRR5p5mtXp2/mAt5q21 2R;
RCRRMp8Rm
t;
-
-RRRRVOkM0MHFRQR1hXR5RH:RM R)q2pRR0sCkRsM)p qR
H#-R-RRRRRR-R-R#7CObsH0MHF:-
-RRRRRRRR-R-RRRRRR1RRCVCRk0MOHRFM8DCON0sNHRFMHQMR R  1R084nj(34.-g
gn-R-RRRRRR-R-R0hFC
#:-R-RRRRRR-R-RRRRRRRRRRN215Qh-RX2=1R-QXh52-
-RRRRRRRR-R-RRRRRRLRR2QR1h25XRX=RRRHVq5A1X<2RR1 u
R--RRRRR-RR-RRRRRRRR2RORh1Q5RX2=RRX-*RX*dd/!VRHR1 uRq<RAX152RR<A q1_1 u
R--RRRRR-RR-RRRRRRRR2R8Rh1Q5avq]Q_u_ me)R_.-2RXRB=RmX152-
-RRRRRRRR-R-RRRRRRCRR2mRB125XR4=R3-jRR6j3**X*.VRHR1qA5RX2<uR 1-
-RRRRRRRR-R-RRRRRRVRR2mRB125XR4=R3-jRR6j3**X*.RR+5*X*cc2/!VRH
R--RRRRR-RR-RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRuR 1q<RAX152AR<q_1  
u1---
-RRRRRRRRMOF#M0N0uR 1RR:)p qRR:=A q1_1 u*1Aq u_ 1-;R-FRBMsPCoOCMCsROHs0CH-N
--
-RRRRRRRRPHNsNCLDR:hRRaQh )t ;-
-RRRRRRRRPHNsNCLDRth qeaQ RR:Apmm Rqh:X=RRj<R3
j;-R-RRRRRRNRPsLHNDXCRpqmBpRR:)p qRR:=q5A1X;2R
R--RRRRRPRRNNsHLRDCezqp ):R ;qp
R--RRRRRPRRNNsHLRDCau vR):R ;qp

---R-RRCRLo
HM-R-RRRRRR-R-R	vNCpRXmpBqRv<Rq_a].Q_u
R--RRRRRHRRVpRXmpBqRv>Rq_a].Q_uRC0EM-
-RRRRRRRRRRRRRRRRau vRR:=wmpm)p5XmpBq/avq]__.u;Q2
R--RRRRRRRRRRRRRXRRpqmBp=R:RmXpBRqp- Ravvu*q_a].Q_u;-
-RRRRRRRRCRM8H
V;---
-RRRRRRRRRHVXBpmq<pRRjj3RC0EM-
--$-#MC0E#RH#0MsN#0DNCV_FV-
-RRRRRRRRRRRRRRRRNC##sw0Rq p1
R--RRRRRRRRRRRRRRRRRRRRRsRRCsbF0XR"pqmBp=R<Rjj3R0NVCssRCO8k0MHFRRHM15QhX
2"-R-RRRRRRRRRRRRRRRRRRRRRRCR#PHCs0 $R)))m;-
--$-#MC0E#RH#0MsN#0DNCM_F
R--RRRRRRRRRRRRRXRRpqmBp=R:Rp-XmpBq;-
-RRRRRRRRCRM8H
V;---
-RRRRRRRRR--BbFlkR0CPkNDCFRVsbR#CNOHDNRO#
C#-R-RRRRRRVRHRmXpBRqp=3RjjFRRspRXmpBqRv=Rq_a].Q_uRRFsXBpmq=pRRavq]Q_uRER0C-M
-RRRRRRRRRRRRRRRR0sCkRsMj;3j
R--RRRRRCRRMH8RV-;
--
-RRRRRRRRHRVRXBpmq=pRRavq]Q_u_ me)R_.0MEC
R--RRRRRRRRRRRRRHRRV RhtQqae0 RE
CM-R-RRRRRRRRRRRRRRRRRRRRRRCRs0MksR3-4j-;
-RRRRRRRRRRRRRRRR#CDC-
-RRRRRRRRRRRRRRRRRRRRRRRRskC0s4MR3
j;-R-RRRRRRRRRRRRRRMRC8VRH;-
-RRRRRRRRCRM8H
V;---
-RRRRRRRRRHVRmXpBRqp=qRvad]___uQm)e _0.RE
CM-R-RRRRRRRRRRRRRRVRHRth qeaQ ER0C-M
-RRRRRRRRRRRRRRRRRRRRRRRR0sCkRsM4;3j
R--RRRRRRRRRRRRRCRRD
#C-R-RRRRRRRRRRRRRRRRRRRRRRCRs0MksR3-4j-;
-RRRRRRRRRRRRRRRR8CMR;HV
R--RRRRRCRRMH8RV-;
--
-RRRRRRRRHXVRpqmBpRR< Ru10MEC
R--RRRRRRRRRRRRRHRRV RhtQqae0 RE
CM-R-RRRRRRRRRRRRRRRRRRRRRRCRs0MksRp-XmpBq;-
-RRRRRRRRRRRRRRRRCCD#
R--RRRRRRRRRRRRRRRRRRRRRsRRCs0kMpRXmpBq;-
-RRRRRRRRRRRRRRRRCRM8H
V;-R-RRRRRRDRC#-C
-RRRRRRRRRRRRRRRRRHVXBpmq<pRR1Aq u_ 1ER0C-M
-RRRRRRRRRRRRRRRRRRRRRRRRva u=R:RmXpBRqp-XR5pqmBpp*XmpBq*mXpB2qp/jn3;-
-RRRRRRRRRRRRRRRRRRRRRRRRHhVR atqQRe 0MEC
R--RRRRRRRRRRRRRRRRRRRRRRRRRRRRRsRRCs0kMaR- ;vu
R--RRRRRRRRRRRRRRRRRRRRRCRRD
#C-R-RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRCRs0MksRva u-;
-RRRRRRRRRRRRRRRRRRRRRRRR8CMR;HV
R--RRRRRRRRRRRRRCRRMH8RV-;
-RRRRRRRR8CMR;HV

---R-RRRRRR Rav:uR=qRvau]_QRR-XBpmq
p;-R-RRRRRRVRHR1qA5va u<2RR1 uRC0EM-
-RRRRRRRRRRRRRRRRHhVR atqQRe 0MEC
R--RRRRRRRRRRRRRRRRRRRRRsRRCs0kMaR- ;vu
R--RRRRRRRRRRRRRCRRD
#C-R-RRRRRRRRRRRRRRRRRRRRRRCRs0MksRva u-;
-RRRRRRRRRRRRRRRR8CMR;HV
R--RRRRRCRRD
#C-R-RRRRRRRRRRRRRRVRHR1qA5va u<2RR1Aq u_ 1ER0C-M
-RRRRRRRRRRRRRRRRRRRRRRRRva u=R:Rva uRR-5va u *avau* 2vu/jn3;-
-RRRRRRRRRRRRRRRRRRRRRRRRHhVR atqQRe 0MEC
R--RRRRRRRRRRRRRRRRRRRRRRRRRRRRRsRRCs0kMaR- ;vu
R--RRRRRRRRRRRRRRRRRRRRRCRRD
#C-R-RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRCRs0MksRva u-;
-RRRRRRRRRRRRRRRRRRRRRRRR8CMR;HV
R--RRRRRRRRRRRRRCRRMH8RV-;
-RRRRRRRR8CMR;HV

---R-RRRRRR Rav:uR=qRva.]__RuQ-pRXmpBq;-
-RRRRRRRRHqVRAa15 2vuR <Ru01RE
CM-R-RRRRRRRRRRRRRRVRHRth qeaQ ER0C-M
-RRRRRRRRRRRRRRRRRRRRRRRR0sCkRsMau v;-
-RRRRRRRRRRRRRRRRCCD#
R--RRRRRRRRRRRRRRRRRRRRRsRRCs0kMaR- ;vu
R--RRRRRRRRRRRRRCRRMH8RV-;
-RRRRRRRR#CDC-
-RRRRRRRRRRRRRRRRHqVRAa15 2vuRA<Rq_1  Ru10MEC
R--RRRRRRRRRRRRRRRRRRRRRaRR Rvu:a=R Rvu-aR5 *vuau v*va un2/3
j;-R-RRRRRRRRRRRRRRRRRRRRRRVRHRth qeaQ ER0C-M
-RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR0sCkRsMau v;-
-RRRRRRRRRRRRRRRRRRRRRRRRCCD#
R--RRRRRRRRRRRRRRRRRRRRRRRRRRRRRsRRCs0kMaR- ;vu
R--RRRRRRRRRRRRRRRRRRRRRCRRMH8RV-;
-RRRRRRRRRRRRRRRR8CMR;HV
R--RRRRRCRRMH8RV-;
--
-RRRRRRRRau vRR:=q5A1v]qa__uQm)e _-.RRmXpB2qp;-
-RRRRRRRRHaVR Rvu<uR 1ER0C-M
-RRRRRRRRRRRRRRRRva u=R:Rj43Ra-R *vuau v*6j3;-
-RRRRRRRRRRRRRRRRHhVR atqQRe 0MEC
R--RRRRRRRRRRRRRRRRRRRRRsRRCs0kMaR- ;vu
R--RRRRRRRRRRRRRCRRD
#C-R-RRRRRRRRRRRRRRRRRRRRRRCRs0MksRva u-;
-RRRRRRRRRRRRRRRR8CMR;HV
R--RRRRRCRRD
#C-R-RRRRRRRRRRRRRRVRHRva uRR<A q1_1 uRC0EM-
-RRRRRRRRRRRRRRRRRRRRRRRRau vRR:=4R3j-va u *avju*3+6RRva u *avau* *vuau v/3.cj-;
-RRRRRRRRRRRRRRRRRRRRRRRRRHVhq ta QeRC0EM-
-RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRskC0s-MRau v;-
-RRRRRRRRRRRRRRRRRRRRRRRRCCD#
R--RRRRRRRRRRRRRRRRRRRRRRRRRRRRRsRRCs0kM Rav
u;-R-RRRRRRRRRRRRRRRRRRRRRRMRC8VRH;-
-RRRRRRRRRRRRRRRRCRM8H
V;-R-RRRRRRMRC8VRH;-
-
R--RRRRRaRR Rvu:q=RAv15q_a]dQ_u_ me)R_.-pRXmpBq2-;
-RRRRRRRRRHVau vR <Ru01RE
CM-R-RRRRRRRRRRRRRR Rav:uR=3R4jRR-au v*va u3*j6-;
-RRRRRRRRRRRRRRRRRHVhq ta QeRC0EM-
-RRRRRRRRRRRRRRRRRRRRRRRRskC0saMR ;vu
R--RRRRRRRRRRRRRCRRD
#C-R-RRRRRRRRRRRRRRRRRRRRRRCRs0MksR -av
u;-R-RRRRRRRRRRRRRRMRC8VRH;-
-RRRRRRRRCCD#
R--RRRRRRRRRRRRRHRRV Rav<uRR1Aq u_ 1ER0C-M
-RRRRRRRRRRRRRRRRRRRRRRRRva u=R:Rj43R -avau* *vujR36+ Ravau* *vuau v*va uc/.3
j;-R-RRRRRRRRRRRRRRRRRRRRRRVRHRth qeaQ ER0C-M
-RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR0sCkRsMau v;-
-RRRRRRRRRRRRRRRRRRRRRRRRCCD#
R--RRRRRRRRRRRRRRRRRRRRRRRRRRRRRsRRCs0kMaR- ;vu
R--RRRRRRRRRRRRRRRRRRRRRCRRMH8RV-;
-RRRRRRRRRRRRRRRR8CMR;HV
R--RRRRRCRRMH8RV-;
--
-RRRRRRRR-B-RFklb0PCRNCDkRsVFRMoCCDsNR#ONC-#
-RRRRRRRRRHV5p5XmpBqRv<Rq_a]umQ_e_ ).RR2NRM85mXpBRqp>3RjjR220MEC
S--SRSSezqp R:=PF_OsO8H_8lFCF_s0HN0FRM5iRB,j,3jRRG,.R(,4
2;-R-RRRRRRRRRRRRRR-RR-qRep:z =BRRmQ)7Bi5RBj,R3Rj,G.,R(),RmaaqQ2mh5;42
R--RRRRRCRRMH8RV-;
--
-RRRRRRRRh=R:RaQh )t Rw5Rp)mm5mXpB/qpv]qa__uQm)e _2.2;-
-RRRRRRRROCN#RqTz7h)qah5RR8lFRRc2H-#
-RRRRRRRRRRRIMECR=jR>-
-SSSSezqp R:=PF_OsO8H_8lFCF_s0HN0FRM5iRB,j,3jRmXpB,qpR,.(R;42
R--RRRRRRRRRRRRR-RR-peqz: R=mRB)B7Q5BRi,3RjjX,RpqmBp.,R(),RmaaqQ2mh5;42
R--RRRRRRRRRERIC4MRR
=>-S-SSqSep:z =_RPO8FsHlO_F_8CsNF00MHF5BRi,3RjjX,RpqmBpRR-v]qa__uQm)e _R.,.R(,j
2;-R-RRRRRRRRRRRRRR-R-ezqp =R:R)Bm75QBR,iBRjj3,pRXmpBqRv-Rq_a]umQ_e_ )..,R(-,
-RRRRRRRRRRRRRRRRR--RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR)RRmaaqQ2mh5;j2
R--RRRRRRRRRERIC.MRR
=>-S-SSqSep:z =PR-_sOF8_HOlCF8_0sFNF0HMi5RBj,R3Rj,XBpmq-pRRavq]Q_u,(R.,2R4;-
-RRRRRRRRRRRRRRRR-q-epRz :-=RB7m)QRB5iRB,j,3jRmXpBRqp-qRvau]_Q.,R(),RmaaqQ2mh5;42
R--RRRRRRRRRERICdMRR
=>-S-SRSRRSpeqz= :R_-PO8FsHlO_F_8CsNF00MHF5BRi,3RjjX,RpqmBpRR-v]qa_ud_Qe_m .)_,(R.,2Rj;-
-RRRRRRRRRRRRRRRR-q-epRz :-=RB7m)QRB5iRB,j,3jRmXpBRqp-qRvad]___uQm)e _R.,.
(,-R-RRRRRRRRRRRRRR-R-RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR)qmaahQm225j;-
-RRRRRRRRCRM8OCN#;-
-
R--RRRRRHRRV RhtQqae0 RE
CM-R-RRRRRRRRRRRRRRCRs0MksRq-ep;z 
R--RRRRRCRRD
#C-R-RRRRRRRRRRRRRRCRs0MksRpeqz
 ;-R-RRRRRRMRC8VRH;-
-RRRRCRM81;Qh
-

-RRRVOkM0MHFR1BmRR5X:MRHRq) ps2RCs0kM R)qHpR#-
-RRRRRRRR-7-RCs#OHHb0F
M:-R-RRRRRR-R-RRRRRRRR1RCCVOkM0MHFRO8CDNNs0MHFRRHMQ   R810R(4jn-3.4ngg
R--RRRRR-RR-FRh0:C#
R--RRRRR-RR-RRRRRRRRRN2B5m1-RX2=mRB125X
R--RRRRR-RR-RRRRRRRRRL2B5m1X=2RRh1Q5avq]Q_u_ me)R_.-2RX
R--RRRRR-RR-RRRRRRRRRO2B5m1v]qa_RuQ+2RXRRR=-1Bm5
X2-R-RRRRRR-R-RRRRRRRR8B2RmX152RR=4R3j-*RXX3/.jVRHR1qA5RX2<uR 1-
-RRRRRRRR-R-RRRRRR2RCR1Bm5RX2=3R4jRR-j*36X.**R5+RXc**2!/cR
HV-R-RRRRRR-R-RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR RRuR1<q5A1X<2RA q1_1 u
R--RRRRR-RR--
-RRRRRRRRO#FM00NMR1 uR):R Rqp:A=Rq_1  *u1A q1_1 u;-
-
R--RRRRRPRRNNsHLRDCXBpmq:pRRq) p=R:R1qA5;X2
R--RRRRRPRRNNsHLRDCezqp ):R ;qp
R--RRRRRPRRNNsHLRDCau vR):R ;qp

---R-RRCRLo
HM-R-RRRRRR-R-R	vNCpRXmpBqRv<Rq_a].Q_u
R--RRRRRHRRVpRXmpBqRv>Rq_a].Q_uRC0EM-
-RRRRRRRRRRRRRRRRau vRR:=wmpm)p5XmpBq/avq]__.u;Q2
R--RRRRRRRRRRRRRXRRpqmBp=R:RmXpBRqp- Ravvu*q_a].Q_u;-
-RRRRRRRRCRM8H
V;---
-RRRRRRRRRHVXBpmq<pRRjj3RC0EM-
--$-#MC0E#RH#0MsN#0DNCV_FV-
-RRRRRRRRRRRRRRRRNC##sw0Rq p1
R--RRRRRRRRRRRRRRRRRRRRRsRRCsbF0XR"pqmBp=R<Rjj3R0NVCssRCO8k0MHFRRHMB5m1X
2"-R-RRRRRRRRRRRRRRRRRRRRRRCR#PHCs0 $R)))m;-
--$-#MC0E#RH#0MsN#0DNCM_F
R--RRRRRRRRRRRRRXRRpqmBp=R:Rp-XmpBq;-
-RRRRRRRRCRM8H
V;---
-RRRRRRRRR--BbFlkR0CPkNDCFRVsbR#CNOHDNRO#
C#-R-RRRRRRVRHRmXpBRqp=3RjjFRRspRXmpBqRv=Rq_a].Q_uRC0EM-
-RRRRRRRRRRRRRRRRskC0s4MR3
j;-R-RRRRRRMRC8VRH;-
-
R--RRRRRHRRVXRRpqmBpRR=v]qa_RuQ0MEC
R--RRRRRRRRRRRRRsRRCs0kM4R-3
j;-R-RRRRRRMRC8VRH;-
-
R--RRRRRHRRVpRXmpBqRv=Rq_a]umQ_e_ ).sRFRmXpBRqp=qRvad]___uQm)e _0.RE
CM-R-RRRRRRRRRRRRRRCRs0MksRjj3;-
-RRRRRRRRCRM8H
V;---
-RRRRRRRRva u=R:R1qA5mXpB2qp;-
-RRRRRRRRH5VRRva uRR< 2u1RC0EM-
-RRRRRRRRRRRRRRRRskC0s5MR4R3j-3Rj6 *avau* 2vu;-
-RRRRRRRRCCD#
R--RRRRRRRRRRRRRHRRVaR5 Rvu<qRA1  _uR120MEC
R--RRRRRRRRRRRRRRRRRRRRRsRRCs0kM4R53-jRj*36au v*va uRR+au v*va u *avau* /vu.jc32-;
-RRRRRRRRRRRRRRRR8CMR;HV
R--RRRRRCRRMH8RV-;
--
-RRRRRRRRau vRR:=q5A1XBpmq-pRv]qa_u._Q
2;-R-RRRRRRVRHRa5R Rvu<uR 102RE
CM-R-RRRRRRRRRRRRRRCRs0MksR354jRR-j*36au v*va u
2;-R-RRRRRRDRC#-C
-RRRRRRRRRRRRRRRRRHV5va uRR<A q1_1 u2ER0C-M
-RRRRRRRRRRRRRRRRRRRRRRRR0sCkRsM5j43R3-j6 *avau* Rvu+ Ravau* *vuau v*va uc/.3;j2
R--RRRRRRRRRRRRRCRRMH8RV-;
-RRRRRRRR8CMR;HV

---R-RRRRRR Rav:uR=ARq1XR5pqmBpRR-v]qa_2uQ;-
-RRRRRRRRHaVR Rvu<uR 1ER0C-M
-RRRRRRRRRRRRRRRR0sCkRsM53-4jRR+j*36au v*va u
2;-R-RRRRRRDRC#-C
-RRRRRRRRRRRRRRRRRHV5va uRR<A q1_1 u2ER0C-M
-RRRRRRRRRRRRRRRRRRRRRRRR0sCkRsM53-4jjR+3a6* *vuau vRa-R *vuau v*va u *av.u/c23j;-
-RRRRRRRRRRRRRRRRCRM8H
V;-R-RRRRRRMRC8VRH;-
-
R--RRRRR-RR-FRBl0bkCNRPDRkCVRFsoCCMsRNDOCN##-
-RRRRRRRRskC0s1MRQvh5q_a]umQ_e_ ).RR-XBpmq;p2
R--RMRC8mRB1
;
RVRRk0MOHRFMaRqh5:XRRRHM)p q2CRs0MksRq) p#RH
RRRRRRRRR--7OC#s0HbH:FM
RRRRRRRRR--RRRRR1RRCVCRk0MOHRFM8DCON0sNHRFMHQMR R  1R084nj(34.-g
gnRRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRNa2Rqjh53Rj2=3RjjR
RRRRRR-R-RRRRRRRRLa2Rq-h5X=2RRq-ah25X
RRRRRRRRR--RRRRRORR2CR)0Mks# R)qpp'mFWRMsRCsRFsHXVRRj<R3Rj
RRRRR-RR-RRRRRRRRR82)kC0sRM#)p q't]Q]MRFRsCsFHsRVRRX>3RjjR

RRRRRPRRNNsHLRDChq ta QeRA:Rm mpq:hR=RRX<3RjjR;
RRRRRPRRNNsHLRDCXBpmq:pRRq) p=R:R1qA5RX2;R
RRRRRRNRPsLHNDeCRq pz: R)q
p;RRRRRRRRPHNsNCLDRva uRR:)p q;R

RLRRCMoH
RRRRRRRRR--vCN	Rjj3RR<=XBpmq<pR=qRva.]__
uQRRRRRRRRHXVRpqmBpRR>v]qa_u._QER0CRM
RRRRRRRRRRRRRaRR Rvu:w=Rp)mm5mXpB/qpv]qa_u._Q
2;RRRRRRRRRRRRRRRRXBpmq:pR=pRXmpBqRa-R *vuv]qa_u._QR;
RRRRRCRRMH8RV
;
RRRRRRRRHXVRpqmBpRR<jR3j0MEC
#--$EM0C##HRN0sMN#D0FC_VRV
RRRRRRRRRRRRRNRR#s#C0qRwp
1 RRRRRRRRRRRRRRRRRRRRRRRRsFCbs"0RXBpmq<pR=3RjjVRN0RCsskC8OF0HMMRHRhaq5"X2
RRRRRRRRRRRRRRRRRRRRRRRRP#CC0sH$)R );m)
#--$EM0C##HRN0sMN#D0FC_MR
RRRRRRRRRRRRRRpRXmpBqRR:=-mXpB;qp
RRRRRRRR8CMR;HV
R
RRRRRR-R-RCBEOP	RN8DHHR0$FNVRslokC
M0RRRRRRRRHXVRpqmBpRR=v]qa__uQm)e _0.RE
CMRRRRRRRRRRRRRRRRNC##sw0Rq p1
RRRRRRRRRRRRRRRRRRRRRRRRbsCFRs0"HXR#RRNl0kDHCbDRRFVv]qa__uQm)e _H.RMqRah25X"R
RRRRRRRRRRRRRRRRRRRRRRCR#PHCs0 $R)))m;R
RRRRRRRRRRRRRRVRHRth qeaQ ER0CRM
RRRRRRRRRRRRRRRRRRRRRsRRCs0kM 5)qpp'm;W2
RRRRRRRRRRRRRRRR#CDCR
RRRRRRRRRRRRRRRRRRRRRRCRs0Mks5q) pQ']t;]2
RRRRRRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMR;HV
R
RRRRRRVRHRmXpBRqp=qRvad]___uQm)e _0.RE
CMRRRRRRRRRRRRRRRRNC##sw0Rq p1
RRRRRRRRRRRRRRRRRRRRRRRRbsCFRs0"HXR#RRNl0kDHCbDRRFVv]qa_ud_Qe_m .)_RRHMa5qhX
2"RRRRRRRRRRRRRRRRRRRRRRRR#CCPs$H0R) )m
);RRRRRRRRRRRRRRRRHhVR atqQRe 0MEC
RRRRRRRRRRRRRRRRRRRRRRRR0sCk5sM)p q't]Q]
2;RRRRRRRRRRRRRRRRCCD#
RRRRRRRRRRRRRRRRRRRRRRRR0sCk5sM)p q'Wpm2R;
RRRRRRRRRRRRRCRRMH8RVR;
RRRRRCRRMH8RV
;
RRRRRRRR-B-RFklb0PCRNCDkRsVFRC#bODHNR#ONCR#
RRRRRHRRVpRXmpBqRj=R3FjRspRXmpBqRv=Rq_a]u0QRE
CMRRRRRRRRRRRRRRRRskC0sjMR3
j;RRRRRRRRCRM8H
V;
RRRRRRRRR--BbFlkR0CPkNDCFRVsCRoMNCsDNRO#
C#RRRRRRRRezqp =R:Rh1Q5mXpB2qp/1Bm5mXpB2qp;R
RRRRRRVRHRth qeaQ ER0CRM
RRRRRRRRRRRRRsRRCs0kMeR-q pz;R
RRRRRRDRC#RC
RRRRRRRRRRRRRsRRCs0kMqRep;z 
RRRRRRRR8CMR;HV
RRRCRM8a;qh
R
RRMVkOF0HM)RqBh1QRR5X:MRHRq) pRR2skC0s)MR RqpHR#
RRRRR-RR-CR7#HOsbF0HMR:
RRRRR-RR-RRRRRRRRC1CRMVkOF0HMCR8OsDNNF0HMMRHR Q  0R18jR4(.n3-g4gnR
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRR2RNRBq)15Qh-RX2=qR-)QB1h25X
RRRRRRRRR--RRRRRLRR2CR)0Mks#RRXFCMRsssF
R
RRRRRRNRPsLHNDhCR atqQRe :mRAmqp h=R:R<XRRjj3;R
RRRRRRNRPsLHNDXCRpqmBpRR:)p qRR:=q5A1X
2;RRRRRRRRPHNsNCLDRpeqz: RRq) p
;
RLRRCMoH
RRRR-RR-ERBCRO	PHND8$H0RRFVNksol0CM#R
RRRRRHXVRpqmBpRR>4R3j0MEC
RRRRRRRR#RN#0CsRpwq1R 
RRRRRRRRRRRRRsRRCsbF0qR"AX152RR>4R3jHqMR)QB1h25X"R
RRRRRRRRRRRRRRCR#PHCs0 $R)))m;R
RRRRRRsRRCs0kM;RX
RRRRCRRMH8RV
;
RRRRR-R-RlBFbCk0RDPNkVCRF#sRbHCONODRN##C
RRRRHRRVpRXmpBqRj=R30jRE
CMRRRRRRRRR0sCkRsMj;3j
RRRRCRRDV#HRmXpBRqp=3R4jER0CRM
RRRRRRRRHhVR atqQRe 0MEC
RRRRRRRRRRRRRRRR0sCkRsM-avq]Q_u_ me);_.
RRRRRRRRDRC#RC
RRRRRRRRRRRRRsRRCs0kMqRvau]_Qe_m .)_;R
RRRRRRCRRMH8RVR;
RRRRR8CMR;HV
R
RRRRR-B-RFklb0PCRNCDkRsVFRMoCCDsNR#ONCR#
RRRRRRHVXBpmq<pRRgj3RC0EMR
RRRRRReRRq pzRR:=qa)BqXh5pqmBp1/5T5)a4R3j-pRXmpBq*mXpB2qp2
2;RRRRRDRC#RC
RRRRRRRRezqp =R:Ravq]Q_u_ me)R_.-)RqBhaq5)1Ta354jRR-XBpmqXp*pqmBpX2/pqmBp
2;RRRRRMRC8VRH;R

RRRRRRHVhq ta QeRC0EMR
RRRRRReRRq pzRR:=-peqz
 ;RRRRRMRC8VRH;R

RRRRR0sCkRsMezqp R;
RMRC8)RqBh1Q;R

RkRVMHO0FqMR)mBB1XR5RH:RM R)qRp2skC0s)MR RqpHR#
RRRRR-RR-CR7#HOsbF0HMR:
RRRRR-RR-RRRRRRRRC1CRMVkOF0HMCR8OsDNNF0HMMRHR Q  0R18jR4(.n3-g4gnR
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRR2RNRBq)B5m1-RX2=qRvau]_QRR-qB)BmX152R
RRRRRR-R-RRRRRRRRL)2RCs0kMX#RRRFMCFsssR

RRRRRPRRNNsHLRDChq ta QeRA:Rm mpq:hR=RRX<3RjjR;
RRRRRPRRNNsHLRDCXBpmq:pRRq) p=R:R1qA5;X2
RRRRRRRRsPNHDNLCqRepRz : R)q
p;
RRRLHCoMR
RRRRR-B-RE	CORDPNH08H$VRFRoNskMlC0R
RRRRRHXVRpqmBpRR>4R3j0MEC
RRRRRRRR#RN#0CsRpwq1R 
RRRRRRRRRRRRRsRRCsbF0qR"AX152RR>4R3jHqMR)mBB125X"R
RRRRRRRRRRRRRRCR#PHCs0 $R)))m;R
RRRRRRsRRCs0kM;RX
RRRRCRRMH8RV
;
RRRRR-R-RlBFbCk0RDPNkVCRF#sRbHCONODRN##C
RRRRHRRVRRX=3R4jER0CRM
RRRRRRRRskC0sjMR3
j;RRRRRDRC#RHVXRR=jR3j0MEC
RRRRRRRRCRs0MksRavq]Q_u_ me);_.
RRRRCRRDV#HR=XRR3-4jER0CRM
RRRRRRRRskC0svMRq_a]u
Q;RRRRRMRC8VRH;R

RRRRRR--BbFlkR0CPkNDCFRVsCRoMNCsDNRO#
C#RRRRRVRHRmXpBRqp>3RjgER0CRM
RRRRRRRRezqp =R:RBq)a5qh1aT)5j43RX-RpqmBpp*XmpBq2p/XmpBq2R;
RRRRR#CDCR
RRRRRReRRq pzRR:=v]qa__uQm)e _-.RRBq)a5qhXBpmq1p/T5)a4R3j-pRXmpBq*mXpB2qp2R;
RRRRR8CMR;HV
R

RRRRRRHVhq ta QeRC0EMR
RRRRRReRRq pzRR:=v]qa_RuQ-qRep;z 
RRRRCRRMH8RV
;
RRRRRCRs0MksRpeqz
 ;RCRRMq8R)mBB1
;

RRRVOkM0MHFRBq)aRqh5:YRRRHM)p q2CRs0MksRq) p#RH
RRRRRRRRR--7OC#s0HbH:FM
RRRRRRRRR--RRRRR1RRCVCRk0MOHRFM8DCON0sNHRFMHQMR R  1R084nj(34.-g
gnRRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRNq2R)qBahY5-2RR=-Bq)a5qhYR2
RRRRR-RR-RRRRRRRRRL2qa)BqYh52RR=-Bq)a5qh4/3jY+2RRavq]Q_u_ me)R_.VRFs|RY|>3R4jR
RRRRRR-R-RRRRRRRROq2R)qBah25YRY=RRsVFR||YR <Ru
1
RRRRRRRRO#FM00NMR1 uR):R Rqp:A=Rq_1  *u1A q1_1 u*1Aq u_ 1
;
RRRRRRRRPHNsNCLDRth qeaQ RR:Apmm Rqh:Y=RRj<R3
j;RRRRRRRRPHNsNCLDRB) Qmu)BRqp:mRAmqp hR;
RRRRRPRRNNsHLRDCYBpmq:pRRq) p=R:R1qA5;Y2
RRRRRRRRsPNHDNLCqRepRz : R)q
p;
RRRLHCoMR
RRRRR-v-RNR	CNksol0CMR||YR4<=3Rj
RRRRRRHVYBpmq>pRRj43RC0EMR
RRRRRRRRRRRRRRpRYmpBqRR:=4/3jYBpmq
p;RRRRRRRRRRRRRRRR)Q BuB)mq:pR=)Raz
 ;RRRRRDRC#RC
RRRRRRRRRRRRR)RR uBQ)qmBp=R:Rpwq1
 ;RRRRRMRC8VRH;R

RRRRRR--BbFlkR0CPkNDCFRVsbR#CNOHDNRO#
C#RRRRRVRHRmYpBRqp=3RjjER0CRM
RRRRRRRRH)VR uBQ)qmBpER0CRM
RRRRRRRRRRRRRHRRV RhtQqae0 RE
CMRRRRRRRRRRRRRRRRRRRRRRRRskC0s5MR-avq]Q_u_ me)2_.;R
RRRRRRRRRRRRRRDRC#RC
RRRRRRRRRRRRRRRRRRRRRsRRCs0kMvR5q_a]umQ_e_ ).
2;RRRRRRRRRRRRRRRRCRM8H
V;RRRRRRRRR#CDCR
RRRRRRRRRRRRRRCRs0MksRjj3;R
RRRRRRCRRMH8RVR;
RRRRR8CMR;HV
R
RRRRRHYVRpqmBpRR< Ru10MEC
RRRRRRRRVRHRth qeaQ ER0CRM
RRRRRRRRRRRRRHRRV R)B)QumpBqRC0EMR
RRRRRRRRRRRRRRRRRRRRRRCRs0MksRv5-q_a]umQ_e_ ).RR+YBpmq;p2
RRRRRRRRRRRRRRRR#CDCR
RRRRRRRRRRRRRRRRRRRRRRCRs0MksRp-YmpBq;R
RRRRRRRRRRRRRRMRC8VRH;R
RRRRRRCRRD
#CRRRRRRRRRRRRRRRRH)VR uBQ)qmBpER0CRM
RRRRRRRRRRRRRRRRRRRRRsRRCs0kMvR5q_a]umQ_e_ ).RR-YBpmq;p2
RRRRRRRRRRRRRRRR#CDCR
RRRRRRRRRRRRRRRRRRRRRRCRs0MksRmYpB;qp
RRRRRRRRRRRRRRRR8CMR;HV
RRRRRRRRMRC8VRH;R
RRRRRCRM8H
V;
RRRR-RR-FRBl0bkCNRPDRkCVRFsoCCMsRNDOCN##R
RRRRRezqp =R:RmRB)B7Q53R4jY,RpqmBpj,R3Rj,.R(,ea Bmh)Qt5R2.
2;
RRRRHRRV R)B)QumpBqRC0EMR
RRRRRReRRq pzRR:=v]qa__uQm)e _-.RRpeqz
 ;RRRRRMRC8VRH;R

RRRRRRHVhq ta QeRC0EMR
RRRRRRqRepRz :-=Rezqp R;
RRRRR8CMR;HV
R
RRRRRskC0seMRq pz;R
RR8CMRBq)a;qh
R

RkRVMHO0FqMR)qBahYR5RH:RM R)qRp;XRR:H)MR 2qpR0sCkRsM)p qR
H#RRRRRRRR-7-RCs#OHHb0F
M:RRRRRRRR-R-RRRRRRCR1CkRVMHO0F8MRCNODsHN0FHMRM RQ 1 R048Rj3(n.g-4gRn
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRRRRN)2RCs0kMj#R3FjRMsRCs
Fs
RRRRRRRRsPNHDNLCpRYmpBqR):R ;qp
RRRRRRRRsPNHDNLCqRepRz : R)q
p;RLRRCMoH
R
RR-RR-ERBCRO	PHND8$H0RRFVNksol0CM#R
RRHRRVYR5Rj=R3NjRMX8RRj=R32jRRC0EMR
RRRRRRRRRR#N#CRs0w1qp CRsb0Fs
RRRRRRRRRRRRRRRR)"qBhaq5jj3,3RjjH2R#MRk8CC0sMlHC
8"RRRRRRRRRRRRRRRR#CCPs$H0R) )m
);RRRRRRRRRsRRCs0kM3RjjR;
RRRRCRM8H
V;
RRRR-R-RlBFbCk0RDPNkVCRF#sRbHCONODRN##C
RRRRVRHR=YRRjj3RC0EMR
RRRRRRVRHR>XRRjj3RC0EMR
RRRRRRRRRR0sCkRsMj;3j
RRRRRRRR#CDCR
RRRRRRRRRR0sCkRsMv]qa_;uQ
RRRRRRRR8CMR;HV
RRRRMRC8VRH;R

RRRRHXVRRj=R30jRE
CMRRRRRRRRHYVRRj>R30jRE
CMRRRRRRRRRsRRCs0kMqRvau]_Qe_m .)_;R
RRRRRRDRC#RC
RRRRRRRRRCRs0MksRq-vau]_Qe_m .)_;R
RRRRRRMRC8VRH;R
RRCRRMH8RV
;

RRRR-R-RlBFbCk0RDPNkVCRFosRCsMCNODRN##C
RRRRpRYmpBqRR:=q5A1Y2/X;R

RRRRezqp =R:RBq)a5qhYBpmq;p2
R
RRHRRVRRX<3RjjER0CRM
RRRRRRRRezqp =R:Ravq]Q_uRe-Rq pz;R
RRCRRMH8RV
;
RRRRRRHVYRR<jR3j0MEC
RRRRRRRRqRepRz :-=Rezqp R;
RRRRCRM8H
V;
RRRRCRs0MksRpeqz
 ;RCRRMq8R)qBah
;

RRRRMVkOF0HMQR1h5]RXRR:H)MR 2qpR0sCkRsM)p qR
H#RRRRRRRR-7-RCs#OHHb0F
M:RRRRRRRR-R-RRRRRRCR1CkRVMHO0F8MRCNODsHN0FHMRM RQ 1 R048Rj3(n.g-4gRn
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRNRR2CR)0Mks# R5XXu52RR- 5Xu-2X2/j.3
RRRRRRRRR--RRRRRLRR2QR1h-]5X=2RRh1Q]25X
R
RRRRRRNRPsLHNDhCR atqQRe :mRAmqp h=R:R<XRRjj3;R
RRRRRRNRPsLHNDXCRpqmBpRR:)p qRR:=q5A1X
2;RRRRRRRRPHNsNCLDRva uRR:)p q;R
RRRRRRNRPsLHNDeCRq pzR):R ;qp
R
RRCRLo
HMRRRRRRRR-B-RFklb0PCRNCDkRsVFRC#bODHNR#ONCR#
RRRRRHRRVpRXmpBqRj=R30jRE
CMRRRRRRRRRRRRRRRRskC0sjMR3
j;RRRRRRRRCRM8H
V;
RRRRRRRRR--BbFlkR0CPkNDCFRVsCRoMNCsDNRO#
C#RRRRRRRRau vRR:= 5XuXBpmq;p2
RRRRRRRRpeqz: R=aR5 Rvu-3R4j /av*u2j;36
R
RRRRRRHRRV RhtQqae0 RE
CMRRRRRRRRRRRRRRRRezqp =R:Rq-ep;z 
RRRRRRRR8CMR;HV
R
RRRRRRCRs0MksRpeqz
 ;RRRRCRM81]Qh;R

RVRRk0MOHRFMR1Bm]XR5RH:RM R)qRp2skC0s)MR RqpHR#
RRRRR-RR-CR7#HOsbF0HMR:
RRRRR-RR-RRRRRRRRC1CRMVkOF0HMCR8OsDNNF0HMMRHR Q  0R18jR4(.n3-g4gnR
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRR2RNR0)Ck#sMRX5 u25XR +RX-u5X/22.
3jRRRRRRRR-R-RRRRRR2RLR1Bm]X5-2RR=B]m15
X2
RRRRRRRRsPNHDNLCpRXmpBqR):R Rqp:q=RAX152R;
RRRRRPRRNNsHLRDCau vR):R ;qp
RRRRRRRRsPNHDNLCqRepRz : R)q
p;RRRRLHCoMR
RRRRRR-R-RlBFbCk0RDPNkVCRF#sRbHCONODRN##C
RRRRRRRRRHVXBpmq=pRRjj3RC0EMR
RRRRRRRRRRRRRRCRs0MksRj43;R
RRRRRRMRC8VRH;


RRRRRRRR-B-RFklb0PCRNCDkRsVFRMoCCDsNR#ONCR#
RRRRRaRR Rvu: =RXXu5pqmBp
2;RRRRRRRRezqp =R:R 5av+uRRj43/va uj2*3
6;
RRRRRRRR0sCkRsMezqp R;
RCRRMB8Rm;1]
R
RRkRVMHO0FRMRa]qhRR5X:MRHRq) ps2RCs0kM R)qHpR#R
RRRRRR-R-R#7CObsH0MHF:R
RRRRRR-R-RRRRRRRR1RCCVOkM0MHFRO8CDNNs0MHFRRHMQ   R810R(4jn-3.4ngg
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRRRN2)kC0sRM#5u X5RX2-XR uX5-252/ 5XuX+2RRu X52-X2R
RRRRRR-R-RRRRRRRRLa2Rq5h]-RX2=aR-q5h]X
2
RRRRRRRRPHNsNCLDRth qeaQ RR:Apmm Rqh:X=RRj<R3
j;RRRRRRRRPHNsNCLDRmXpBRqp: R)q:pR=ARq125X;R
RRRRRRNRPsLHNDaCR Rvu: R)q
p;RRRRRRRRPHNsNCLDRpeqz: RRq) p
;
RRRRLHCoMR
RRRRRR-R-RlBFbCk0RDPNkVCRF#sRbHCONODRN##C
RRRRRRRRRHVXBpmq=pRRjj3RC0EMR
RRRRRRRRRRRRRRCRs0MksRjj3;R
RRRRRRMRC8VRH;R

RRRRR-RR-FRBl0bkCNRPDRkCVRFsoCCMsRNDOCN##R
RRRRRR Rav:uR=XR up5XmpBq2R;
RRRRReRRq pzRR:=5va uRR-4/3jau v2a/5 Rvu+3R4j /av;u2
R
RRRRRRVRHRth qeaQ ER0CRM
RRRRRRRRRsRRCs0kMeR-q pz;R
RRRRRRDRC#RC
RRRRRRRRRsRRCs0kMqRep;z 
RRRRRRRR8CMR;HV
RRRR8CMRhaq]
;
RRRRVOkM0MHFRBq)1]QhRR5X:MRHRq) ps2RCs0kM R)qHpR#R
RRRRRR-R-R#7CObsH0MHF:R
RRRRRR-R-RRRRRRRR1RCCVOkM0MHFRO8CDNNs0MHFRRHMQ   R810R(4jn-3.4ngg
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRRRN2)kC0sRM#p5mtR+XRR)1TaX5R*+XRRj432
2
RRRRLHCoMR
RRRRRR-R-RlBFbCk0RDPNkVCRF#sRbHCONODRN##C
RRRRRRRRRHVXRR=jR3j0MEC
RRRRRRRRRRRRRRRR0sCkRsMj;3j
RRRRRRRR8CMR;HV
R
RRRRRR-R-RlBFbCk0RDPNkVCRFosRCsMCNODRN##C
RRRRRRRR0sCkRsM5mRptX5RR1+RT5)aRXX*R4+R32j2R
2;RRRRCRM8q1)BQ;h]



RVRRk0MOHRFMqB)BmR1]5:XRRRHM)p q2CRs0MksRq) p#RH
RRRRRRRRR--7OC#s0HbH:FM
RRRRRRRRR--RRRRR1RRCVCRk0MOHRFM8DCON0sNHRFMHQMR R  1R084nj(34.-g
gnRRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRN)2RCs0kMp#RmRt5XRR+1aT)5*RXXRR-423j2R;RR>XR=3R4jR
RRRRRR-R-RRRRRRRRL)2RCs0kMX#RRRFMCFsssR

RLRRCMoH
RRRRRRRRR--BOEC	NRPDHH80F$RVsRNoCklM
0#RRRRRRRRHXVRR4<R30jRE
CMRRRRRRRRRRRRRRRRR#N#CRs0w1qp R
RRRRRRRRRRRRRRRRRRRRRRCRsb0FsRR"X<3R4jMRHRBq)B]m15"X2
RRRRRRRRRRRRRRRRRRRRRRRRP#CC0sH$)R );m)
RRRRRRRRRRRRRRRRCRs0MksR
X;RRRRRRRRCRM8H
V;
RRRRRRRRR--BbFlkR0CPkNDCFRVsbR#CNOHDNRO#
C#RRRRRRRRHXVRR4=R30jRE
CMRRRRRRRRRRRRRRRRskC0sjMR3
j;RRRRRRRRCRM8H
V;
RRRRRRRRR--BbFlkR0CPkNDCFRVsCRoMNCsDNRO#
C#RRRRRRRRskC0s5MRRtpm5RRX+TR1)Ra5XR*X-3R4j222;R
RRMRC8)RqB1Bm]
;
RRRRVOkM0MHFRBq)a]qhRR5X:MRHRq) ps2RCs0kM R)qHpR#R
RRRRRR-R-R#7CObsH0MHF:R
RRRRRR-R-RRRRRRRR1RCCVOkM0MHFRO8CDNNs0MHFRRHMQ   R810R(4jn-3.4ngg
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRRRN2)kC0sRM#5tpm54R53+jRR/X25j43RX-R2/22.R3j;RR|XRR|<3R4jR
RRRRRR-R-RRRRRRRRL)2RCs0kMX#RRRFMCFsssR
RRCRLo
HMRRRRRRRR-B-RE	CORDPNH08H$VRFRoNskMlC0R#
RRRRRHRRVARq125XRR>=4R3j0MEC
RRRRRRRRRRRRRRRR#N#CRs0w1qp R
RRRRRRRRRRRRRRRRRRRRRRCRsb0FsRA"q125XRR>=4R3jHqMR)qBahX]52R"
RRRRRRRRRRRRRRRRRRRRR#RRCsPCHR0$ m)))R;
RRRRRRRRRRRRRsRRCs0kM;RX
RRRRRRRR8CMR;HV
R
RRRRRR-R-RlBFbCk0RDPNkVCRF#sRbHCONODRN##C
RRRRRRRRRHVXRR=jR3j0MEC
RRRRRRRRRRRRRRRR0sCkRsMj;3j
RRRRRRRR8CMR;HV
R
RRRRRR-R-RlBFbCk0RDPNkVCRFosRCsMCNODRN##C
RRRRRRRR0sCk5sMR6j3*tpm54R53Xj+24/53Xj-2RR22R;
RCRRMq8R)qBah
];
8CMRqRva)]_ ;qp
