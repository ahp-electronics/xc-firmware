--
@ER--B$FbsEHo0OR52gR4g-cRRj.jd$R1MHbDO$H0ROQM
R--fN]C8:CsR#//$DMbH0OH$N/lb0DN.Uj4J4.b/blNb#Cs/0N0/LDH/MoC_OFsN/cCs_NlsPI3E48yR-f
-


---
--
-Rl1HbRDC)RqvIEH0RM#HoRDCq)77 R11VRFss8CNR8NMRHIs0-C
-NRas0oCRp:RkMOC0RR-mq)BR
c -D-
HNLssH$RC;CC
Ck#RCHCC03#8F_Do_HO4c4n3DND;#
kCCRHC#C30D8_FOoH_o#HM3C8N;DD
Ck#RCHCC03#8F_Do_HON0sHED3ND-;
-LDHs$NsROFsN
c;-#-kCsRFO3NcFNsOObFl3DND;-
-Ns00H0LkC$R#MD_LN_O	LRFGF)VRB. dX:cRRlOFbCFMMH0R#sR0k
C;
0CMHR0$)_qv)HWR#R
RRCRoMHCsO
R5RRRRRRRRVHNlDR$:#H0sM:oR=MR"F"MC;R
RRRRRRHRI8R0E:MRH0CCos=R:RR(;
RRRRRRRR8N8s8IH0:ERR0HMCsoCRR:=(R;RRRRRR-R-RoLHRFCMkRoEVRFs80CbER
RRRRRRCR8bR0E:MRH0CCos=R:R.R4UR;
RRRRR8RRF_k0sRCo:FRLFNDCM=R:RDVN#RC;RRRR-E-RNF#Rkk0b0CRsoR
RRRRRRHR8MC_soRR:LDFFCRNM:V=RNCD#;RRRR-RR-NRE#NR80HNRM0bkRosC
RRRRRRRR8N8sC_soRR:LDFFCRNM:V=RNCD#RRRRR-R-R8ENRNsC88RN8#sC#CRsoR
RRRRRR;R2
RRRRsbF0
R5RRRRRRRR7amzRRR:FRk0#_08DHFoOC_POs0F58IH04E-RI8FMR0Fj
2;RRRRRRRR7RQhRRR:HRMR#_08DHFoOC_POs0F58IH04E-RI8FMR0Fj
2;RRRRRRRRq)77RRR:HRMR#_08DHFoOC_POs0F58N8s8IH04E-RI8FMR0Fj
2;RRRRRRRRWR RRRR:HRMR#_08DHFoOR;RRRRRRR--I0sHCMRCNCLDRsVFRlsN
RRRRRRRRiBpR:RRRRHMR8#0_oDFHRO;RRRRR-R-RFODOV	RFssRNRl,Ns88,HR8MR
RRRRRRBRmpRiR:MRHR0R#8F_DoRHORRRRR-RR-bRF0DROFRO	VRFs80Fk
RRRRRRRR
2;CRM8CHM00)$Rq)v_W
;
---
-HRwsR#0HDlbCMlC0HN0FlMRkR#0LOCRNCDD8sRNO
Ej-N-
sHOE00COkRsCNEsOjVRFRv)q_R)WHO#
FFlbM0CMRh1q7RU
b0FsRR5
RRRq:MRHR8#0_oDFH
O;RARRRH:RM0R#8F_Do;HO
RRRBRR:H#MR0D8_FOoH;R
RR:7RRRHM#_08DHFoOR;
RRR :MRHR8#0_oDFH
O;RwRRRH:RM0R#8F_Do;HO
RRRtRR:H#MR0D8_FOoH;R
RR:]RRRHM#_08DHFoOR;
RRRZ:kRF00R#8F_Do
HOR
2;CRM8ObFlFMMC0O;
FFlbM0CMRh1q7Rn
b0FsRR5
RRRq:MRHR8#0_oDFH
O;RARRRH:RM0R#8F_Do;HO
RRRBRR:H#MR0D8_FOoH;R
RR:7RRRHM#_08DHFoOR;
RRR :MRHR8#0_oDFH
O;RwRRRH:RM0R#8F_Do;HO
RRRZRR:FRk0#_08DHFoO2
R;M
C8FROlMbFC;M0
lOFbCFMM10Rqch7
FRbs50R
RRRqRR:H#MR0D8_FOoH;R
RR:ARRRHM#_08DHFoOR;
RRRB:MRHR8#0_oDFH
O;R7RRRH:RM0R#8F_Do;HO
RRRZRR:FRk0#_08DHFoO2
R;M
C8FROlMbFC;M0
lOFbCFMM10Rq.h7
FRbs50R
RRRqRR:H#MR0D8_FOoH;R
RR:ARRRHM#_08DHFoOR;
RRRZ:kRF00R#8F_Do
HOR
2;CRM8ObFlFMMC0
;
ObFlFMMC0qR1hj74
FRbs50R
RRRqRR:H#MR0D8_FOoH;R
RR:ARRRHM#_08DHFoOR;
RRRB:MRHR8#0_oDFH
O;R7RRRH:RM0R#8F_Do;HO
RRR RR:H#MR0D8_FOoH;R
RR:wRRRHM#_08DHFoOR;
RRRt:MRHR8#0_oDFH
O;R]RRRH:RM0R#8F_Do;HO
RRRQRR:H#MR0D8_FOoH;R
RR:KRRRHM#_08DHFoOR;
RRRZ:kRF00R#8F_Do
HOR
2;CRM8ObFlFMMC0O;
FFlbM0CMR )Bdc.X
FRbs50R
RRRqR7j:MRHR8#0_oDFH
O;RqRR7:4RRRHM#_08DHFoOR;
R7Rq.RR:H#MR0D8_FOoH;R
RRdq7RH:RM0R#8F_Do;HO
RRRqR7c:MRHR8#0_oDFH
O;R7RRQ:jRRRHM#_08DHFoOR;
RQR74RR:H#MR0D8_FOoH;R
RR.7QRH:RM0R#8F_Do;HO
RRR7RQd:MRHR8#0_oDFH
O;RBRRiRR:H#MR0D8_FOoH;R
RR)t1RH:RM0R#8F_Do;HO
RRRWh) RH:RM0R#8F_Do;HO
RRRWju RH:RM0R#8F_Do;HO
RRRW4u RH:RM0R#8F_Do;HO
RRR7Rmj:kRF00R#8F_Do;HO
RRR7Rm4:kRF00R#8F_Do;HO
RRR7Rm.:kRF00R#8F_Do;HO
RRR7Rmd:kRF00R#8F_Do;HO
RRRTj7mRF:Rk#0R0D8_FOoH;R
RRmT74RR:FRk0#_08DHFoOR;
R7RTm:.RR0FkR8#0_oDFH
O;RTRR7Rmd:kRF00R#8F_Do
HOR
2;CRM8ObFlFMMC0O;
F0M#NRM0M_klODCD#C_8C:bRR0HMCsoCRR:=5C58bR0E-2R4/2d.;RRRRRRRR-R-RFyRVFRsIF#RVBR) Xd.cCRODRD#M8CCCO8
F0M#NRM0M_klODCD#H_I8:CRR0HMCsoCRR:=5H5I8R0E-2R4/;c2RRRRRRRRR-R-RFyRVFRODMkl#VRFR )Bdc.XRDOCDM#RCCC88$
0bFCRkL0_k0#_$RbCHN#Rs$sNRk5MlC_OD_D#8bCCRI8FMR0Fj5,RM_klODCD#H_I8cC*2R+d8MFI0jFR2VRFR8#0_oDFH
O;#MHoNFDRkL0_kR#RRF:RkL0_k0#_$;bCRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RVFR8k50RHkMb0FR0RH0s-N#002C#
o#HMRNDF_k0CRMRRRR:#_08DHFoOC_POs0F5lMk_DOCD8#_CRCb8MFI0jFR2R;R-C-RMDNLCV#RF0sRs#H-0CN0#H
#oDMNRCIbjM_CR:RRR8#0_oDFHPO_CFO0sk5MlC_OD_D#8bCCRI8FMR0FjR2;RR--I0sHCMRCNCLD#FRVsNRCOsERFFIRVqR)vCROD
D##MHoNIDRb_C4CRMRR#:R0D8_FOoH_OPC05FsM_klODCD#C_8C8bRF0IMF2Rj;-RR-sRIHR0CCLMNDRC#VRFsCENORIsFRRFV)RqvODCD#H
#oDMNR_HMsRCoR:RRR8#0_oDFHPO_CFO0sH5I8+0EdFR8IFM0R;j2RRRRRRRRRR--k8#CRR0FsHCo#s0CRh7QRH
#oDMNR0Fk_osCR:RRR8#0_oDFHPO_CFO0sH5I8+0EdFR8IFM0R;j2RRRRRRRRRR--k8#CRR0FsHCo#s0CRz7maH
#oDMNR_HMs4CoR:RRR8#0_oDFHPO_CFO0sH5I8+0EdFR8IFM0R;j2RRRR
o#HMRNDNs8_CRoRRRR:#_08DHFoOC_POs0F58N8s8IH04E-RI8FMR0FjR2;RRRR-k-R#RC80sFRC#oH0RCsq)77
o#HMRNDD_FINs88RRR:#_08DHFoOC_POs0F58cRF0IMF2Rj;RRRRRRRRRRRRRRR-N-R8R8sL#H0RbHMk00RFqR)vCRODRD#5L6RHR0#skCJH8sC2$
0b0CRlNb_8_8s0C$bRRH#NNss$MR5kOl_C#DD_C8CbFR8IFM0RRj2F#VR0D8_FOoH_OPC0RFs58gRF0IMF2Rj;H
#oDMNRb0l_8N8s:RRRb0l_8N8s$_0b
C;
oLCH
M
RRRR-Q-RV8RN8HsI8R0E<RR6NH##o'MRj0'RFMRkk8#CR0LH#R
RR4RzRRR:H5VRNs88I0H8ERR=4o2RCsMCN
0CRRRRRRRRD_FINs88RR<="jjjj&"RR_N8s5Coj
2;RRRRCRM8oCCMsCN0R;z4
RRRRRz.RH:RVNR58I8sHE80R.=R2CRoMNCs0RC
RRRRRDRRFNI_8R8s<"=Rj"jjRN&R8C_soR548MFI0jFR2R;
RCRRMo8RCsMCNR0Cz
.;RRRRzRdR:VRHR85N8HsI8R0E=2RdRMoCC0sNCR
RRRRRRFRDI8_N8<sR=jR"j&"RR_N8s5Co.FR8IFM0R;j2
RRRR8CMRMoCC0sNCdRz;R
RRcRzRRR:H5VRNs88I0H8ERR=co2RCsMCN
0CRRRRRRRRD_FINs88RR<='Rj'&8RN_osC58dRF0IMF2Rj;R
RRMRC8CRoMNCs0zCRcR;
RzRR6:RRRRHV58N8s8IH0>ERRRc2oCCMsCN0
RRRRRRRRIDF_8N8s=R<R_N8s5CocFR8IFM0R;j2
RRRR8CMRMoCC0sNC6Rz;R

R-RR-VRQRH58MC_sos2RC#oH0RCs7RQhkM#HopRBiR
RRnRzRRR:H5VR8_HMs2CoRMoCC0sNCR
RRRRRRsRbF#OC#BR5pRi,72QhRoLCHRM
RRRRRRRRRHRRVBR5p=iRR''4R8NMRiBp'CCPMR020MEC
RRRRRRRRRRRRRRRR_HMsRCo<5=R"jjjj&"RRh7Q2R;
RRRRRRRRRCRRMH8RVR;
RRRRRCRRMb8RsCFO#
#;RRRRCRM8oCCMsCN0R;zn
RRRRRz(RH:RVMR5F80RHsM_CRo2oCCMsCN0
RRRRRRRRRRRR_HMsRCo<5=R"jjjj&"RRh7Q2R;
RCRRMo8RCsMCNR0Cz
(;
RRRRR--Q5VRNs88_osC2CRso0H#CqsR7R7)kM#HopRBiR
RR4Rz.:RRRRHV58N8sC_soo2RCsMCN
0CRRRRRRRRbOsFCR##5iBp,7Rq7R)2LHCoMR
RRRRRRRRRRVRHRp5BiRR='R4'NRM8B'piCMPC002RE
CMRRRRRRRRRRRRRRRRNs8_C<oR=7Rq7N)58I8sHE80-84RF0IMF2Rj;R
RRRRRRRRRRMRC8VRH;R
RRRRRRMRC8sRbF#OC#R;
RCRRMo8RCsMCNR0Cz;4.
R
RR4RzdRR:H5VRMRF0Ns88_osC2CRoMNCs0RC
RRRRRRRRRNRR8C_so=R<R7q7)85N8HsI8-0E4FR8IFM0R;j2
RRRR8CMRMoCC0sNC4Rzd
;
RRRRzR.nRH:RV8R5F_k0s2CoRMoCC0sNCR
RRRRRRsRbF#OC#mR5B,piR0Fk_osC2CRLo
HMRRRRRRRRRRRRH5VRmiBpR'=R4N'RMm8RB'piCMPC002RE
CMRRRRRRRRRRRRRRRR7amzRR<=F_k0s5CoI0H8ER-48MFI0jFR2R;
RRRRRRRRRCRRMH8RVR;
RRRRRCRRMb8RsCFO#
#;RRRRCRM8oCCMsCN0Rnz.;R

R-RR-CRtMNCs00CRE#CRCODC0FRDo
HORRRRzR4c:FRVsRRHHMMRkOl_C#DD_C8CbFR8IFM0RojRCsMCN
0CRRRR-A-Rk8HDR0FkbRk0CLMND#CRCODC0FRDo
HORRRRRRRR-Q-RVNR58I8sHE80R4>R682RF0M'RCk#RQ1pBCROD
D#RRRRRRRRmn 4RH:RVNR58I8sHE80R4>R6o2RCsMCN
0CRRRRRRRRRRRRRRRRF_k0CHM52=R<R''4RCIEMNR58C_so85N8HsI8-0E4FR8IFM0RR62=2RHR#CDCjR''R;
RRRRRCRRMo8RCsMCNR0Cmn 4;R
RRRRRR-R-RRQV58N8s8IH0>ERRR62qRh758N8s8IH0<ER=6R42#RkCpR1QOBRC#DD
RRRRRRRR4m 6RR:H5VRNs88I0H8ERR=4R62oCCMsCN0
RRRRRRRRRRRRRRRRb0l_8N8s25H58gRF0IMF2RjRR<=h5maOPFM_8#0_oDFHPO_CFO0s,5HR24j2mRX)8RN_osC58N8s8IH04E-RI8FMR0F6
2;RRRRRRRRRRRRRRRR17qh_R46:qR1hj74RsbF0NRlbqR5RR=>0_lbNs8855H2jR2,A>R=Rb0l_8N8s25H5,42R=BR>lR0b8_N8Hs5225.,RR7=0>RlNb_858sHd252R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR =0>RlNb_858sHc252w,RRR=>0_lbNs8855H26R2,t>R=Rb0l_8N8s25H5,n2R=]R>lR0b8_N8Hs5225(,RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRQ=0>RlNb_858sHU252K,RRR=>0_lbNs8855H2gR2,Z>R=R0Fk_5CMH;22
RRRRRRRR8CMRMoCC0sNC Rm4
6;RRRRRRRRmc 4RH:RVNR58I8sHE80R4=Rco2RCsMCN
0CRRRRRRRRRRRRRRRR0_lbNs8855H2UFR8IFM0RRj2<h=RmOa5F_MP#_08DHFoOC_POs0F5RH,gR22XRm)Ns8_CNo58I8sHE80-84RF0IMF2R6;R
RRRRRRRRRRRRRRqR1h47_cRR:17qh4bjRFRs0lRNb5=qR>lR0b8_N8Hs5225j,RRA=0>RlNb_858sH4252B,RRR=>0_lbNs8855H2.R2,7>R=Rb0l_8N8s25H5,d2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR >R=Rb0l_8N8s25H5,c2R=wR>lR0b8_N8Hs52256,RRt=0>RlNb_858sHn252],RRR=>0_lbNs8855H2(R2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRQ>R=Rb0l_8N8s25H5,U2R=KR>4R''Z,RRR=>F_k0CHM52
2;RRRRRRRRCRM8oCCMsCN0R4m cR;
RRRRRmRR R4d:VRHR85N8HsI8R0E=dR42CRoMNCs0RC
RRRRRRRRRRRRR0RRlNb_858sH(25RI8FMR0Fj<2R=mRhaF5OM#P_0D8_FOoH_OPC05FsHU,R2X2RmN)R8C_so85N8HsI8-0E4FR8IFM0R;62
RRRRRRRRRRRRRRRRh1q7d_4R1:RqUh7RFRbsl0RN5bRq>R=Rb0l_8N8s25H5,j2R=AR>lR0b8_N8Hs52254,RRB=0>RlNb_858sH.2527,RRR=>0_lbNs8855H2d
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR RRRR=>0_lbNs8855H2cR2,w>R=Rb0l_8N8s25H5,62R=tR>lR0b8_N8Hs5225n,RR]=0>RlNb_858sH(252
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRZRRRR=>F_k0CHM52
2;RRRRRRRRCRM8oCCMsCN0R4m dR;
RRRRRmRR R4.:VRHR85N8HsI8R0E=.R42CRoMNCs0RC
RRRRRRRRRRRRR0RRlNb_858sHn25RI8FMR0Fj<2R=mRhaF5OM#P_0D8_FOoH_OPC05FsH(,R2X2RmN)R8C_so85N8HsI8-0E4FR8IFM0R;62
RRRRRRRRRRRRRRRRh1q7._4R1:RqUh7RFRbsl0RN5bRq>R=Rb0l_8N8s25H5,j2R=AR>lR0b8_N8Hs52254,RRB=0>RlNb_858sH.2527,RRR=>0_lbNs8855H2d
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR RRRR=>0_lbNs8855H2cR2,w>R=Rb0l_8N8s25H5,62R=tR>lR0b8_N8Hs5225n,RR]='>R4R',
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRZ>R=R0Fk_5CMH;22
RRRRRRRR8CMRMoCC0sNC Rm4
.;RRRRRRRRm4 4RH:RVNR58I8sHE80R4=R4o2RCsMCN
0CRRRRRRRRRRRRRRRR0_lbNs8855H26FR8IFM0RRj2<h=RmOa5F_MP#_08DHFoOC_POs0F5RH,nR22XRm)Ns8_CNo58I8sHE80-84RF0IMF2R6;R
RRRRRRRRRRRRRRqR1h47_4RR:17qhnbRRFRs0lRNb5=qR>lR0b8_N8Hs5225j,RRA=0>RlNb_858sH4252B,RRR=>0_lbNs8855H2.R2,7>R=Rb0l_8N8s25H5,d2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR >R=Rb0l_8N8s25H5,c2R=wR>lR0b8_N8Hs52256,RRZ=F>RkC0_M25H2R;
RRRRRCRRMo8RCsMCNR0Cm4 4;R
RRRRRR Rm4:jRRRHV58N8s8IH0=ERR24jRMoCC0sNCR
RRRRRRRRRRRRRRlR0b8_N8Hs52R5c8MFI0jFR2=R<Rahm5MOFP0_#8F_Do_HOP0COFHs5,2R62mRX)8RN_osC58N8s8IH04E-RI8FMR0F6
2;RRRRRRRRRRRRRRRR17qh_R4j:qR1hR7nRsbF0NRlbqR5RR=>0_lbNs8855H2jR2,A>R=Rb0l_8N8s25H5,42R=BR>lR0b8_N8Hs5225.,RR7=0>RlNb_858sHd252R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR =0>RlNb_858sHc252w,RRR=>',4'R=ZR>kRF0M_C52H2;R
RRRRRRMRC8CRoMNCs0mCR ;4j
RRRRRRRRgm RRR:H5VRNs88I0H8ERR=go2RCsMCN
0CRRRRRRRRRRRRRRRR0_lbNs8855H2dFR8IFM0RRj2<h=RmOa5F_MP#_08DHFoOC_POs0F5RH,cR22XRm)Ns8_CNo58I8sHE80-84RF0IMF2R6;R
RRRRRRRRRRRRRRqR1hg7_R1:Rqch7RbRRFRs0lRNb5=qR>lR0b8_N8Hs5225j,RRA=0>RlNb_858sH4252B,RRR=>0_lbNs8855H2.R2,7>R=Rb0l_8N8s25H5,d2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRZ>R=R0Fk_5CMH;22
RRRRRRRR8CMRMoCC0sNC RmgR;
RRRRRmRR RUR:VRHR85N8HsI8R0E=2RURMoCC0sNCR
RRRRRRRRRRRRRRlR0b8_N8Hs52R5.8MFI0jFR2=R<Rahm5MOFP0_#8F_Do_HOP0COFHs5,2Rd2mRX)8RN_osC58N8s8IH04E-RI8FMR0F6
2;RRRRRRRRRRRRRRRR17qh_:URRh1q7RcRRsbF0NRlbqR5RR=>0_lbNs8855H2jR2,A>R=Rb0l_8N8s25H5,42R=BR>lR0b8_N8Hs5225.,RR7='>R4
',RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRZRRRR=>F_k0CHM52
2;RRRRRRRRCRM8oCCMsCN0RUm ;R
RRRRRR Rm(:RRRRHV58N8s8IH0=ERRR(2oCCMsCN0
RRRRRRRRRRRRRRRRb0l_8N8s25H584RF0IMF2RjRR<=h5maOPFM_8#0_oDFHPO_CFO0s,5HR2.2R)XmR_N8s5CoNs88I0H8ER-48MFI06FR2R;
RRRRRRRRRRRRR1RRq_h7(RR:17qh.RRRb0FsRblNRR5q=0>RlNb_858sHj252A,RRR=>0_lbNs8855H24R2,Z>R=R0Fk_5CMH;22
RRRRRRRR8CMRMoCC0sNC Rm(R;
RRRRRmRR RnR:VRHR85N8HsI8R0E=2RnRMoCC0sNCR
RRRRRRRRRRRRRRkRF0M_C5RH2<'=R4I'RERCM5_N8s5Co6=2RRMOFP0_#8F_Do_HOP0COFHs5,542jR22CCD#R''j;R
RRRRRRMRC8CRoMNCs0mCR 
n;RRRR-Q-RVNR58I8sHE80RR<=6M2RFkRF00bkRNCMLRDC#CCDOD0RFOoHRCMC8RC8/NRlbHR8s0COD0$RFqR)vR'#Ns88CR##DCHM#R
RRRRRR Rm6RR:H5VRNs88I0H8E=R<RR62oCCMsCN0
RRRRRRRRRRRRRRRR0Fk_5CMH<2R=4R''R;
RRRRRCRRMo8RCsMCNR0Cm; 6
R
RR-R-RRQV58N8s8IH0>ERRRg2kR#CWju RR0F8FCO8NCR8C8s#L#RHR0#nER0soFkERRgNRM8W4u RR0F8FCO8LCRHR0#4+jR
RRRRRRRR4W jRR:H5VRNs88I0H8ERR>go2RCsMCN
0CRRRRRRRRRRRRRRRRIjbC_5CMH<2R=4R''ERIC5MRNs8_CUo5RI8FMR0F6=2RRMOFP0_#8F_Do_HOP0COFHs5,2.j58dRF0IMF2Rj2DRC#'CRj
';RRRRRRRRRRRRRRRRI4bC_5CMH<2R=4R''ERIC5MRNs8_CNo58I8sHE80-84RF0IMF2RgRO=RF_MP#_08DHFoOC_POs0F5.H,jN258I8sHE80-8nRF0IMF2Rc2DRC#'CRj
';RRRRRRRRRRRRCRM8oCCMsCN0R4W jR;
R-RR-VRQR85N8HsI8R0E=RRUFgsR2#RkCuRW 0jRFCR8OCF8R8N8s#C#R0LH#RRn0FEskRoEgR
RRRRRR RWg:RRRRHV585N8HsI8R0E=2RURRm)58N8s8IH0=ERR2g2RMoCC0sNCR
RRRRRRRRRRRRRRbRICCj_M25HRR<='R4'IMECR85N_osC58N8s8IH04E-RI8FMR0F6=2RRRH2CCD#R''j;R
RRRRRRRRRRRRRRbRICC4_M25HRR<=';4'
RRRRRRRRRRRR8CMRMoCC0sNC RWgR;
R-RR-VRQR85N8HsI8R0E=2R(RCk#R WujFR0RO8CFR8C0RECnR0ENs88CR##LRH0&uRW 04RFCR8OCF8RC0ERE(0R8N8s#C#R0LH
RRRRRRRR(W RRR:H5VRNs88I0H8ERR=(o2RCsMCN
0CRRRRRRRRRRRRRRRRIjbC_5CMH<2R=4R''ERIC5MRNs8_C6o52RR=OPFM_8#0_oDFHPO_CFO0s,5H.j252C2RDR#C';j'
RRRRRRRRRRRRRRRRCIb4M_C5RH2<'=R4I'RERCM5_N8s5Con=2RRMOFP0_#8F_Do_HOP0COFHs5,5.24R22CCD#R''j;R
RRRRRRMRC8CRoMNCs0WCR 
(;RRRR-Q-RVNR58I8sHE80Rn=R2#RkCuRW 0jRFCR8OCF8RC0EREn0R8N8s#C#R0LH
RRRRRRRRnW RRR:H5VRNs88I0H8ERR=no2RCsMCN
0CRRRRRRRRRRRRRRRRIjbC_5CMH<2R=4R''ERIC5MRNs8_C6o52RR=OPFM_8#0_oDFHPO_CFO0s,5H4j252C2RDR#C';j'
RRRRRRRRRRRRRRRRCIb4M_C5RH2<'=R4
';RRRRRRRRCRM8oCCMsCN0RnW ;R
RR-R-RRQV58N8s8IH0<ER=2R6RRMFI0sHCMRCNCLDRD#CCRO0DHFoOCRMC88C
RRRRRRRR6W RRR:H5VRNs88I0H8E=R<RR62oCCMsCN0
RRRRRRRRRRRRRRRRCIbjM_C5RH2<'=R4
';RRRRRRRRRRRRRRRRI4bC_5CMH<2R=4R''R;
RRRRRCRRMo8RCsMCNR0CW; 6
R
RRMRC8CRoMNCs0zCR4
c;
RRRR6z.RH:RVMR5F80RF_k0s2CoRMoCC0sNCR
RRRRRR4Rz(R4:bOsFCR##50Fk_osC2R
RRRRRRCRLo
HMRRRRRRRRRRRR7amzRR<=F_k0s5CoI0H8ER-48MFI0jFR2R;
RRRRRCRRMb8RsCFO#z#R4;(4
RRRR8CMRMoCC0sNC.Rz6
;
RRRR-t-RCsMCNR0C0REC)RqvODCD#HRI00ERs#H-0CN0#R
RR4Rz6RR:VRFsHMRHRlMk_DOCD8#_CRCb8MFI0jFRRMoCC0sNCR
RRRRRR4Rz(RR:VRFs[MRHRlMk_DOCDI#_HR8C8MFI0jFRRMoCC0sNCR
RRRRRRRRRR)RzqRv:)dB .RXc
RRRRRRRRRRRRRRRRsbF0NRlb7R5Q=jR>MRH_osC5*5[c,22R47QRR=>HsM_C5o5[2*c+,42R.7QRR=>HsM_C5o5[2*c+,.2Rd7QRR=>HsM_C5o5[2*c+,d2R)t1RR=>',4'RR
RRRRRRRRRRRRRRRRRRRRRRRRRqR7j=D>RFNI_858sjR2,qR74=D>RFNI_858s4R2,qR7.=D>RFNI_858s.R2,qR7d=D>RFNI_858sdR2,qR7c=D>RFNI_858scR2,
R--RRRRRRRRRRRRRRRRRRRRRRRRR W)h>R=R,W R Wuj>R=RCIbjM_C5,H2R Wu4>R=RCIb4M_C5,H2RRBi=h>RmBaRpRi,
RRRRRRRRRRRRRRRRRRRRRRRRWRR)R h=W>R W,RuR j=I>Rb_CjCHM52W,RuR 4=I>Rb_C4CHM52B,Ri>R=RiBp,RR
RRRRRRRRRRRRRRRRRRRRRRRRRj7mRR=>F_k0L5k#H[,5*2c2,mR74>R=R0Fk_#Lk55H,[2*c+,42R.7mRR=>F_k0L5k#H[,5*+c2.R2,7Rmd=F>RkL0_kH#5,*5[cd2+2
2;RRRRRRRRRRRRRRRRF_k0s5Co5c[*2<2R=kRF0k_L#,5H5c[*2I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co5c[*22+4RR<=F_k0L5k#H[,5*+c24I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co5c[*22+.RR<=F_k0L5k#H[,5*+c2.I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co5c[*22+dRR<=F_k0L5k#H[,5*+c2dI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRCRM8oCCMsCN0R(z4;R
RRRRRRMRC8CRoMNCs0zCR4
6;
R--RUz.RH:RV8R5F_k0s2CoRMoCC0sNC-
-RRRRRRRRzR4n:FRVsRRHHMMRkOl_C#DD_C8CbFR8IFM0RojRCsMCN
0C-R-RRRRRR4RzURR:VRFs[MRHRlMk_DOCDI#_HR8C8MFI0jFRRMoCC0sNC-
-RRRRRRRRRRRRzv)q:BR) Xd.c-R
-RRRRRRRRRRRRRRRRsbF0NRlb7R5Q=jR>MRH_osC5*5[c,22R47QRR=>HsM_C5o5[2*c+,42R.7QRR=>HsM_C5o5[2*c+,.2Rd7QRR=>HsM_C5o5[2*c+,d2
R--RRRRRRRRRRRRRRRRRRRRRRRRRjq7RR=>D_FINs885,j2R4q7RR=>D_FINs885,42R.q7RR=>D_FINs885,.2Rdq7RR=>D_FINs885,d2Rcq7RR=>D_FINs885,c2
R--RRRRRRRRRRRRRRRRRRRRRRRRR W)h>R=R,W R Wuj>R=RCIbjM_C5,H2R Wu4>R=RCIb4M_C5,H2RRBi=h>RmBaRpRi,
R--RRRRRRRRRRRRRRRRRRRRRRRRRmT7j>R=R0Fk_#Lk55H,[2*c2T,R7Rm4=F>RkL0_kH#5,*5[c42+2T,R7Rm.=F>RkL0_kH#5,*5[c.2+2T,R7Rmd=F>RkL0_kH#5,*5[cd2+2
2;-R-RRRRRRRRRRRRRRkRF0C_so[55*2c2RR<=F_k0L5k#H[,5*2c2RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;-
-RRRRRRRRRRRRRRRRF_k0s5Co5c[*22+4RR<=F_k0L5k#H[,5*+c24I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';-R-RRRRRRRRRRRRRRkRF0C_so[55*+c2.<2R=kRF0k_L#,5H5c[*22+.RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;-
-RRRRRRRRRRRRRRRRF_k0s5Co5c[*22+dRR<=F_k0L5k#H[,5*+c2dI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';-R-RRRRRRRRRRMRC8CRoMNCs0zCR4
U;-R-RRRRRR8CMRMoCC0sNC4Rzn-;
-RRRR8CMRMoCC0sNC.RzU
;
-R-RRRRRk:URRRHV5k8F0C_soo2RCsMCN
0C-R-RRRRRRRRR7amzRR<=F_k0s5CoI0H8ER-48MFI0jFR2-;
-CRRMo8RCsMCNR0Ck
U;RRRRRRRRRRRRRRRRRM
C8sRNO0EHCkO0sNCRsjOE;