--
@ER--RbBF$osHE50RO42RgRgg1b$MDHHO0R$,Q3MO
R--RDqDRosHER0#sCC#s8PC3-
-

---f-R]8CNCRs:/$/#MHbDO$H0/blND.N0jJ4U./b4lbNbC/s#O8bD/LDH/MoC_0DN0CHO/bOl_3D0PyE84
Rf-
-
DsHLNRs$HCCC;#
kCCRHC#C30D8_FOoH_n44cD3NDk;
#HCRC3CC#_08DHFoOs_NH30EN;DD
0CMHR0$ObFlN_sCNkOOlH_L0#RH
FSbs
05SCSbJRR:H#MR0D8_FOoH;S
SbRD0:MRHR8#0_oDFH
O;S0SDHRR:H#MR0D8_FOoH;S
SCRJH:MRHR8#0_oDFH
O;S0SDRF:Rk#0R0D8_FOoH;S
SC:JRR0FkR8#0_oDFHSO
2C;
MO8RFNlbsNC_OlOk_0LH;N

sHOE00COkRsCLDFFCRNMFOVRFNlbsNC_OlOk_0LHR
H#LHCoMC
SJ=R<RJbCR8NMRHCJ;D
S0=R<R0bDRCIEMJRCHRR='R4'CCD#RHD0;M
C8FRLFNDCM
;
-N-ROlOkk0DNCER0C0RDR#sCkRD0VlsFRC0ERCbsPkHF#CRDPRCDObFlN#sC
LDHs$NsRCHCCk;
#HCRC3CC#_08DHFoO4_4nNc3D
D;kR#CHCCC38#0_oDFHNO_sEH03DND;M
C0$H0RlOFbCNs_ONOkHlR#o
SCsMCH5OR
#SSHRxC:MRH0CCos2
S;b
SF5s0
DSS0:HRRRHM#_08DHFoOC_POs0F5x#HCR-48MFI0jFR2S;
SHCJRH:RM0R#8F_Do_HOP0COF#s5H-xC4FR8IFM0R;j2
DSS0RR:FRk0#_08DHFoOS;
SRCJ:kRF00R#8F_Do
HOS
2;CRM8ObFlN_sCNkOOl
;
NEsOHO0C0CksRFLFDMCNRRFVObFlN_sCNkOOl#RH
HS#oDMNR0DDR#:R0D8_FOoH_OPC05Fs#CHxRI8FMR0Fj
2;So#HMRNDDRCJ:0R#8F_Do_HOP0COF#s5HRxC8MFI0jFR2S;
ObFlFMMC0FROlsbNCO_NO_klLRH0HS#
SsbF0S5
SCSbJRR:H#MR0D8_FOoH;S
SS0bDRH:RM0R#8F_Do;HO
SSSDR0H:MRHR8#0_oDFH
O;SCSSJ:HRRRHM#_08DHFoOS;
S0SDRF:Rk#0R0D8_FOoH;S
SSRCJ:kRF00R#8F_Do
HOS;S2
MSC8FROlMbFC;M0
oLCH
MRS0DD5Rj2<'=Rj
';SJDC5Rj2<'=R4
';SRp:VRFsMMRHR0jRFHR#x4C-RMoCC0sNCS
SOO:RFNlbsNC_OlOk_0LHRsbF0NRlb
R5SbSSC=JR>CRDJ25M,S
SSHCJRR=>C5JHM
2,SbSSD=0R>DRD025M,S
SSHD0RR=>D50HM
2,SCSSJ>R=RJDC54M+2S,
S0SDRR=>D5D0M2+4
2SS;C
SMo8RCsMCN;0C
0SDRR<=D5D0#CHx2S;
C<JR=CRDJH5#x;C2
8CMRFLFDMCN;D

HNLssH$RC;CC
Ck#RCHCC03#8F_Do_HO4c4n3DND;#
kCCRHC#C30D8_FOoH_HNs0NE3D
D;CHM00O$RFNlbsLC_HH0R#b
SF5s0
NSSRH:RM0R#8F_Do;HO
LSSRH:RM0R#8F_Do;HO
DSS0:HRRRHM#_08DHFoOS;
SHCJRH:RM0R#8F_Do;HO
DSS0RR:FRk0#_08DHFoOS;
SRCJ:kRF00R#8F_Do
HOS
2;CRM8ObFlN_sCL;H0
s
NO0EHCkO0sLCRFCFDNFMRVFROlsbNCH_L0#RH
oLCH
MRSRCJ<C=RJNHRMM8RF50RNFRGs2RL;D
S0=R<RILRERCM5GNRFLsR2RR='R4'CCD#RHD0;M
C8FRLFNDCM
;
DsHLNRs$HCCC;#
kCCRHC#C30D8_FOoH_n44cD3NDk;
#HCRC3CC#_08DHFoOs_NH30EN;DD
0CMHR0$ObFlNRsCHS#
oCCMsRHO5x#HCRR:HCM0oRCs2S;
b0FsRS5
S:NRRRHM#_08DHFoOC_POs0F5x#HCR-48MFI0jFR2S;
S:LRRRHM#_08DHFoOC_POs0F5x#HCR-48MFI0jFR2S;
SRD0:kRF00R#8F_Do;HO
CSSJRR:FRk0#_08DHFoO2
S;M
C8FROlsbNC
;
NEsOHO0C0CksRFLFDMCNRRFVObFlNRsCHS#
#MHoNbDRDR0,bRCJ:0R#8F_Do_HOP0COF#s5HRxC8MFI0jFR2S;
ObFlFMMC0FROlsbNCH_L0#RH
bSSF5s0
SSSNRR:H#MR0D8_FOoH;S
SS:LRRRHM#_08DHFoOS;
S0SDHRR:H#MR0D8_FOoH;S
SSHCJRH:RM0R#8F_Do;HO
SSSD:0RR0FkR8#0_oDFH
O;SCSSJRR:FRk0#_08DHFoOS
S2S;
CRM8ObFlFMMC0L;
CMoH
CSbJ25jRR<=';4'
DSb025jRR<=';j'
:StRsVFRHMRMRRj0#FRH-xC4CRoMNCs0
CRS:SORlOFbCNs_0LHRS
SSsbF0NRlb
R5SSSSNN=>5,M2RS
SS=SL>ML52
,RSSSSD=0H>0bD5,M2RS
SSJSCHb=>CMJ52
,RSSSSD>0=b5D0M2+4,SR
SCSSJb=>CMJ5+
42S2SS;C
SMo8RCsMCN;0C
0SDRR<=b5D0#CHx2S;
C<JR=CRbJH5#x;C2
8CMRFLFDMCN;D

HNLssH$RC;CC
Ck#RCHCC03#8F_Do_HO4c4n3DND;#
kCCRHC#C30D8_FOoH_HNs0NE3D
D;CHM00B$Rvpu_a#RH
RRRRMoCCOsH58IH0:ERR0HMCsoCRR:=U;j2RR--[
NoRRRRb0Fs5Rq:H#MR0D8_FOoH_OPC05FsI0H8E4R-RI8FMR0Fj
2;RRRRRRRRRRA:H#MR0D8_FOoH_OPC05FsI0H8E4R-RI8FMR0Fj
2;RRRRRRRRRRpa:kRF00R#8F_Do2HO;M
C8vRBua_p;N

sHOE00COkRsCLDFFCRNMFOVRlDb_0#RH
kSVMHO0FOMRNODOM50RO#FM00NMR,#xRNDCVR#x:MRH0CCoss2RCs0kMMRH0CCos#RH
NSPsLHNDDCRC0NVlsb,ORM0:MRH0CCosS;
LHCoMS
SDVCN0Rlb:#=RxRR/DVCN#
x;SVSHR#55xFRl8CRDNxV#2RR=j02RE
CMSsSSORM0:D=RC0NVl;bR
CSSDR#C
SSSs0OMRR:=5NDCVb0lR4+R2S;
S8CMR;HV
sSSCs0kMORsM
0;S8CMRDONO0OM;S

O#FM00NMRXvqBRvu:MRH0CCos=R:R
c;SMOF#M0N0CRDNHV#x:CRR0HMCsoCRR:=vBqXv
u;SMOF#M0N0lROb0OMRH:RMo0CC:sR=NRODMOO0H5I8,0EDVCN#CHx2S;

kSVMHO0FlMRNHGL0OR5F0M#NRM0MRR:HCM0o2CsR0sCkRsMHCM0oRCsHS#
PHNsNCLDRGlNRH:RMo0CC
s;SoLCHSM
SGlNRR:=54M+2C*DNHV#x-CRR
4;SVSHRN5lG=R>R8IH0RE20MEC
SSSlRNG:I=RHE80-
4;SMSC8VRH;S
SskC0slMRN
G;S8CMRGlNL;H0
#
SHNoMDDRo0RR:#_08DHFoOC_POs0F5bOlO-M04FR8IFM0R;j2
HS#oDMNRJoCR#:R0D8_FOoH_OPC05FsOOlbM40-RI8FMR0Fj
2;
FSOlMbFCRM0ObFlNRsCHS#
SMoCCOsHRH5#x:CRR0HMCsoC2S;
SsbF0
R5SNSSRH:RM0R#8F_Do_HOP0COF#s5H-xC4FR8IFM0R;j2
SSSLRR:H#MR0D8_FOoH_OPC05Fs#CHx-84RF0IMF2Rj;S
SSRD0:kRF00R#8F_Do;HO
SSSC:JRR0FkR8#0_oDFHSO
S
2;S8CMRlOFbCFMM
0;SlOFbCFMMO0RFNlbsNC_OlOkR
H#SCSoMHCsO
R5S#SSHRxC:MRH0CCosS
S2S;
SsbF0S5
S0SDHRR:H#MR0D8_FOoH_OPC05Fs#CHx-84RF0IMF2Rj;S
SSHCJRH:RM0R#8F_Do_HOP0COF#s5H-xC4FR8IFM0R;j2
SSSD:0RR0FkR8#0_oDFH
O;SCSSJRR:FRk0#_08DHFoOS
S2S;
CRM8ObFlFMMC0
;
So#HMRNDC:JRR8#0_oDFH
O;
oLCHSM
-k-R#NCRRF0I-PDCCDDRFNF	E8CNRE#OC
lCSRA:H5VRI0H8ERR>vBqXvRu2oCCMsCN0RS
StV:RFMsRRRHMOOlbM40-RI8FMR0FjCRoMNCs0SC
SFSOMN#0Ml0RGRL0:MRH0CCos=R:RGlNL5H0M
2;SOSSF0M#NRM0l0MLRH:RMo0CC:sR=*RMDVCN#CHx;S
SLHCoMS
SSRB:ObFlNRsCoCCMsRHOlRNb5x#HC>R=Rl4+G-L0l0ML2S
SSFSbsl0RN5bR
SSSSRSN=N>R5LlG0FR8IFM0RLlM0
2,SSSSS=LR>5RLl0GLRI8FMR0Fl0ML2S,
SSSSD>0=R0oD5,M2
SSSSJSC=o>RCMJ52S
SS;S2
CSSMo8RCsMCN;0C
S
SNO:RFNlbsNC_OlOkRS
SSMoCCOsHRblNRS5
S#SSHRxC=O>RlMbO0S
SSS2
SFSbsl0RN5bR
SSSSHD0RR=>o,D0
SSSSHCJRR=>o,CJ
SSSSRD0=D>R0S,
SCSSJ>R=R
CJS2SS;C
SMo8RCsMCN;0C
-
S-#RkCRRNsbHbDOCRFNlbsSC
1H:RVIR5HE80RR<=vBqXvRu2oCCMsCN0
BSS:FROlsbNCCRoMHCsONRlb#R5H=xC>8IH0
E2SbSSFRs0lRNb5S
SSRSN=N>R,S
SSRSL=L>R,S
SS0SD=D>R0S,
SCSSJR=>CSJ
S;S2
MSC8CRoMNCs0
C;
8CMRFLFDMCN;



