-- $Header: //synplicity/maplat2018q2p1/mappers/lattice/lib/gen_lava1/inc.vhd#1 $
@ER--H
MO
LDHs$NsR Q  k;
#QCR 3  #_08DHFoO4_4nNc3D
D;
-
-----------------------------------------------------RC

M00H$hRQB#RHRo

CsMCHMO5RH:RMo0CC=s:426c;
R
b0Fs5
R
qRR:H#MR0D8_FOoH_OPC05FsMR-48MFI0jFR2
;R
:1RR0FkR8#0_oDFHPO_CFO0s-5M4FR8IFM0RRj2
;
2RC

MQ8RhRB;
s
NO0EHCkO0spCReh_QBVRFRBQhR
H#
lOFbCFMMe0RBRB
RFRbs
05RRRRRRRXRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR:RFRk0RaR17m_ptRQB:'=R4;'2
8CMRlOFbCFMM
0;
lOFbCFMMt0RhR7
RFRbs
05RRRRRRRXRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR:RFRk0RaR17m_ptRQB:'=Rj;'2
8CMRlOFbCFMM
0;
lOFbCFMMB0RBqz_7R7
RFRbs
05RRRRRjRqRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR:RHRMRRaR17m_pt;QB
RRRRARRjRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR:RRHMR1RRap7_mBtQ;R
RRRRRBRQhRRRRRRRRRRRRRRRRRRRRRRRRR:RRRMRHRRRR1_a7pQmtBR;
RRRRRR1jRRRRRRRRRRRRRRRRRRRRRRRRRRRR:FRRkR0RR71a_tpmQ
B;RRRRRmRBzRaRRRRRRRRRRRRRRRRRRRRRRRRRRR:RFRk0RaR17m_pt2QB;M
C8FROlMbFC;M0
#

HNoMDNROsRs$RRR:#_08DHFoOC_POs0F5-RM4FR8IFM0R2jR;H
#oDMNRMOF#40_R#:R0D8_FOoH;H
#oDMNRMOF#j0_R#:R0D8_FOoH;L

CMoH
4Sz:BReBmRu)vaRqRu5XR=>O#FM02_4;z
S.t:Rhu7RmR)avRqu5=XR>FROM_#0j
2;RRRRRRRRzRd:B_BzqR77uam)Ruvq55RqjR2,O#FM0,_jRMOF#40_,5R1jR2,OsNs$25j2R;
RRRRRzRRcV:RFHsRRRHM4FR0R4M-RMoCC0sNCR
RRRRRRRRRRRRRR.Rz_Rp4:BRBz7_q7mRu)vaRqRu5q25H,FROM_#0jO,RN$ss54H-21,R5,H2RsONsH$52
2;RRRRRRRRCRM8oCCMsCN0;C

Mp8Reh_QB
;

