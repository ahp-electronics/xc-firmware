--
@ER--B$FbsEHo0OR52gR4g-cRRj.jd$R1MHbDO$H0ROQM
R--fN]C8:CsR#//$DMbH0OH$N/lb0DN.Uj4J4.b/blNb#Cs/DGHH/MGD/HLoCCMs/HOo_CMoCCMs/HOs_Nls_IbsE3P8Ry4f-
-
-
--R--Bp pRqX)vXd.4-7R----
LDHs$NsRCHCCk;
#HCRC3CC#_08DHFoO4_4nNc3D
D;kR#CHCCC38#0_oDFH#O_HCoM8D3NDD;
HNLssk$RMHH#lk;
#kCRMHH#lO3PFFlbM0CM#D3ND
;
CHM00X$R)dqv.7X4R
H#RFRbs50R
RRRRRRRRm7uR:RRR0FkR8#0_FkDo;HORRRRRRRR
RRRRRRRRm1uR:RRR0FkR8#0_FkDo;HO
R
RRRRRRjRqRRRR:MRHR8#0_FkDo;HO
RRRRRRRRRq4R:RRRRHM#_08koDFH
O;RRRRRRRRqR.RRRR:H#MR0k8_DHFoOR;
RRRRRqRRdRRRRH:RM0R#8D_kFOoH;R
RRRRRRcRqRRRR:MRHR8#0_FkDo;HO
RRRRRRRRR7RR:RRRRHM#_08koDFH
O;RRRRRRRR7qu)jRR:H#MR0k8_DHFoOR;
RRRRR7RRu4)qRH:RM0R#8D_kFOoH;R
RRRRRRuR7)Rq.:MRHR8#0_FkDo;HO
RRRRRRRR)7uq:dRRRHM#_08koDFH
O;RRRRRRRR7qu)cRR:H#MR0k8_DHFoOR;
RRRRRWRRBRpiRH:RM0R#8D_kFOoH;RRRRRRRRR
RRRRRR RWRRRR:MRHR8#0_FkDo
HORRRRR2RR;
RRCRM8Xv)qd4.X7N;
sHOE00COkRsCXv)qd4.X7R_eFXVR)dqv.7X4R
H#R#RSHNoMDCRIjI,RCR4,#,FjR4#F,FR8j8,RFR4:#_08DHFoOL;
CMoH
uS7m=R<Rj8FRCIEM7R5uc)qR'=RjR'2CCD#R48F;1
Su<mR=FR#jERIC5MRq=cRR''j2DRC##CRF
4;SjICRR<=WN RM58RMRF0q;c2
CSI4=R<RRW NRM8q
c;RjSzR):Rqnv4XR47
RRRRRRRRRRRRRRRRsbF0NRlb7R5RR=>7q,Rj>R=R,qjRRq4=q>R4q,R.>R=R,q.RRqd=q>RdR,
S7SSuj)qRR=>7qu)j7,Ru4)qRR=>7qu)47,Ru.)qRR=>7qu).7,Rud)qRR=>7qu)d
,RSWSS >R=RjIC,BRWp=iR>BRWpRi,7Rum=8>RFRj,1Rum=#>RF;j2
zRS4RR:)4qvn7X4RR
RRRRRRRRRRRRRRFRbsl0RN5bR7>R=RR7,q=jR>jRq,4RqRR=>qR4,q=.R>.Rq,dRqRR=>q
d,RSSS7qu)j>R=R)7uqRj,7qu)4>R=R)7uqR4,7qu).>R=R)7uqR.,7qu)d>R=R)7uqRd,
SSSW= R>CRI4W,RBRpi=W>RB,piRm7uRR=>8,F4Rm1uRR=>#2F4;M
C8)RXq.vdX_47e
;
----- RBpXpR)nqvc7X4R----D-
HNLssH$RC;CC
Ck#RCHCC03#8F_Do_HO4c4n3DND;#
kCCRHC#C30D8_FOoH_o#HM3C8N;DD
LDHs$NsRHkM#;Hl
Ck#RHkM#3HlPlOFbCFMM30#N;DD
M
C0$H0RqX)vXnc4H7R#R
Rb0FsRR5
RRRRR7RRuRmRRF:Rk#0R0k8_DHFoOR;RRRRRRRR
RRRRR1RRuRmRRF:Rk#0R0k8_DHFoO
;
RRRRRRRRqRjRRRR:H#MR0k8_DHFoOR;
RRRRRqRR4RRRRH:RM0R#8D_kFOoH;R
RRRRRR.RqRRRR:MRHR8#0_FkDo;HO
RRRRRRRRRqdR:RRRRHM#_08koDFH
O;RRRRRRRRqRcRRRR:H#MR0k8_DHFoOR;
RRRRRqRR6RRRRH:RM0R#8D_kFOoH;R
RRRRRRRR7RRRR:MRHR8#0_FkDo;HO
RRRRRRRR)7uq:jRRRHM#_08koDFH
O;RRRRRRRR7qu)4RR:H#MR0k8_DHFoOR;
RRRRR7RRu.)qRH:RM0R#8D_kFOoH;R
RRRRRRuR7)Rqd:MRHR8#0_FkDo;HO
RRRRRRRR)7uq:cRRRHM#_08koDFH
O;RRRRRRRR7qu)6RR:H#MR0k8_DHFoOR;
RRRRRWRRBRpiRH:RM0R#8D_kFOoH;RRRRRRRRR
RRRRRR RWRRRR:MRHR8#0_FkDo
HORRRRR2RR;
RRCRM8Xv)qn4cX7N;
sHOE00COkRsCXv)qn4cX7R_eFXVR)nqvc7X4R
H#R#RSHNoMDCRIjI,RCR4,I,C.RdIC,FR#j#,RFR4,#,F.Rd#F,FR8j8,RFR4,8,F.Rd8F:0R#8F_Do;HO
oLCHSM
7Rum<R=R8RFjIMECRu57)Rq6=jR''MRN8uR7)Rqc=jR''C2RDR#C
8SSFI4RERCM5)7uq=6RR''jR8NMR)7uq=cRR''42DRC#
CRSFS8.ERIC5MR7qu)6RR='R4'NRM87qu)cRR='2j'R#CDCSR
Sd8F;1
Su<mR=#RRFIjRERCM5Rq6=jR''MRN8cRqR'=RjR'2CCD#RS
S#RF4IMECR65qR'=RjN'RMq8RcRR='24'R#CDCSR
S.#FRCIEMqR56RR='R4'NRM8q=cRR''j2DRC#
CRSFS#dS;
IRCj<W=R MRN8MR5Fq0R6N2RM58RMRF0q;c2
CSI4=R<RRW NRM850MFR2q6R8NMR;qc
CSI.=R<RRW NRM8qN6RM58RMRF0q;c2
CSId=R<RRW NRM8qN6RMq8RcR;
SRzj:qR)vX4n4
7RRRRRRRRRRRRRRRRRb0FsRblNRR57=7>R,jRqRR=>qRj,q=4R>4Rq,.RqRR=>qR.,q=dR>dRq,S
RSuS7)Rqj=7>Ruj)q,uR7)Rq4=7>Ru4)q,uR7)Rq.=7>Ru.)q,uR7)Rqd=7>Rud)q,SR
S SWRR=>I,CjRpWBi>R=RpWBi7,Ru=mR>FR8j1,Ru=mR>FR#j
2;R4SzR):Rqnv4XR47
RRRRRRRRRRRRRRRRsbF0NRlb7R5RR=>7q,Rj>R=R,qjRRq4=q>R4q,R.>R=R,q.RRqd=q>RdR,
S7SSuj)qRR=>7qu)j7,Ru4)qRR=>7qu)47,Ru.)qRR=>7qu).7,Rud)qRR=>7qu)d
,RSWSS >R=R4IC,BRWp=iR>BRWpRi,7Rum=8>RFR4,1Rum=#>RF;42
zRS.RR:)4qvn7X4RR
RRRRRRRRRRRRRRFRbsl0RN5bR7>R=RR7,q=jR>jRq,4RqRR=>qR4,q=.R>.Rq,dRqRR=>q
d,RSSS7qu)j>R=R)7uqRj,7qu)4>R=R)7uqR4,7qu).>R=R)7uqR.,7qu)d>R=R)7uqRd,
SSSW= R>CRI.W,RBRpi=W>RB,piRm7uRR=>8,F.Rm1uRR=>#2F.;S
Rz:dRRv)q44nX7RR
RRRRRRRRRRRRRbRRFRs0lRNb5=7R>,R7RRqj=q>Rjq,R4>R=R,q4RRq.=q>R.q,Rd>R=R,qd
SRSS)7uq=jR>uR7),qjR)7uq=4R>uR7),q4R)7uq=.R>uR7),q.R)7uq=dR>uR7),qdRS
SSRW =I>RCRd,WiBpRR=>WiBp,uR7m>R=Rd8F,uR1m>R=Rd#F2C;
MX8R)nqvc7X4_
e;

-----
-HR1lCbDRv)qR0IHEHR#MCoDR7q7)1 1RsVFR0LFECRsNN8RMI8RsCH0
R--aoNsC:0RRDXHH
MG-
-
DsHLNRs$HCCC;#
kCCRHC#C30D8_FOoH_n44cD3NDk;
#HCRC3CC#_08DHFoOH_#o8MC3DND;H
DLssN$MRkHl#H;#
kCMRkHl#H3FPOlMbFC#M03DND;M
C0$H0Rv)q_u)W_H)R#o
SCsMCH5OR
RSRRNRVl$HDR#:R0MsHo=R:RF"MM;C"
ISSHE80RH:RMo0CC:sR=;R4RS
SNs88I0H8ERR:HCM0oRCs:n=R;RRRRRRRRR--LRHoCkMFoVERF8sRCEb0
8SSCEb0RH:RMo0CC:sR=URc;S
Ssk8F0C_soRR:LDFFCRNM:V=RNCD#;RRRR-RR-NRE#kRF00bkRosC
ISS80Fk_osCRL:RFCFDN:MR=NRVD;#CS-S-R#ENR0FkbRk0s
CoSHS8MC_soRR:LDFFCRNM:V=RNCD#;RRRRRRRRR--ERN#8NN0RbHMks0RCSo
S8sN8ss_C:oRRFLFDMCNRR:=V#NDCR;RRRRR-E-RNs#RCRN8Ns88CR##s
CoSNSI8_8ssRCo:FRLFNDCM:RR=NRVDR#CRRRRRR--ERN#I0sHC8RN8#sC#CRsoS
S2S;
b0FsRS5
S7)_m:zaR0FkR8#0_oDFHPO_CFO0sH5I8-0E4FR8IFM0R;j2
WSS_z7maRR:FRk0#_08DHFoOC_POs0F58IH04E-RI8FMR0Fj
2;SqS)7R7):MRHR8#0_oDFHPO_CFO0s85N8HsI8-0E4FR8IFM0R;j2
7SSQRhR:MRHR8#0_oDFHPO_CFO0sH5I8-0E4FR8IFM0R;j2
WSSq)77RH:RM0R#8F_Do_HOP0COFNs58I8sHE80-84RF0IMF2Rj;S
SWR R:MRHR8#0_oDFHRO;RRRRR-R-RHIs0CCRMDNLCFRVsNRslS
SBRpi:MRHR8#0_oDFHRO;RRRRR-R-RFODOV	RFssRNRl,Ns88,HR8MS
S)B_mp:iRRRHM#_08DHFoOR;RRRRRRR--FRb0OODF	FRVs_Rs80Fk
WSS_pmBiRR:H#MR0D8_FOoHR-R-FRb0VRFsIF_8kS0
S
2;CRM8CHM00)$Rq)v_W)u_;-

--
-RswH#H0RlCbDl0CMNF0HMkRl#L0RCNROD8DCRONsE-j
-s
NO0EHCkO0sLCRD	FO_lsNRRFV)_qv)_Wu)#RH
lOFbCFMMX0R)dqv.7X4RbRRFRs05R
RRRRRRuR7mRRR:kRF00R#8D_kFOoH;RRRRRRRRR
RRRRRRuR1mRRR:kRF00R#8D_kFOoH;R

RRRRRqRRjRRRRH:RM0R#8D_kFOoH;R
RRRRRR4RqRRRR:MRHR8#0_FkDo;HO
RRRRRRRRRq.R:RRRRHM#_08koDFH
O;RRRRRRRRqRdRRRR:H#MR0k8_DHFoOR;
RRRRRqRRcRRRRH:RM0R#8D_kFOoH;R
RRRRRRRR7RRRR:MRHR8#0_FkDo;HO
RRRRRRRR)7uq:jRRRHM#_08koDFH
O;RRRRRRRR7qu)4RR:H#MR0k8_DHFoOR;
RRRRR7RRu.)qRH:RM0R#8D_kFOoH;R
RRRRRRuR7)Rqd:MRHR8#0_FkDo;HO
RRRRRRRR)7uq:cRRRHM#_08koDFH
O;RRRRRRRRWiBpRRR:H#MR0k8_DHFoOR;RRRRRRRR
RRRRRWRR RRRRH:RM0R#8D_kFOoH
RRRRRRR2R;R
8CMRlOFbCFMM
0;ObFlFMMC0)RXqcvnXR47RFRbs50R
RRRRRRRRm7uR:RRR0FkR8#0_FkDo;HORRRRRRRR
RRRRRRRRm1uR:RRR0FkR8#0_FkDo;HO
R
RRRRRRjRqRRRR:MRHR8#0_FkDo;HO
RRRRRRRRRq4R:RRRRHM#_08koDFH
O;RRRRRRRRqR.RRRR:H#MR0k8_DHFoOR;
RRRRRqRRdRRRRH:RM0R#8D_kFOoH;R
RRRRRRcRqRRRR:MRHR8#0_FkDo;HO
RRRRRRRRRq6R:RRRRHM#_08koDFH
O;RRRRRRRR7RRRRRR:H#MR0k8_DHFoOR;
RRRRR7RRuj)qRH:RM0R#8D_kFOoH;R
RRRRRRuR7)Rq4:MRHR8#0_FkDo;HO
RRRRRRRR)7uq:.RRRHM#_08koDFH
O;RRRRRRRR7qu)dRR:H#MR0k8_DHFoOR;
RRRRR7RRuc)qRH:RM0R#8D_kFOoH;R
RRRRRRuR7)Rq6:MRHR8#0_FkDo;HO
RRRRRRRRpWBi:RRRRHM#_08koDFHRO;RRRRR
RRRRRRRRRRWR RRRR:H#MR0k8_DHFoOR
RRRRRRR2;RM
C8FROlMbFC;M0
MVkOF0HMkRVMHO_M5H0LRR:LDFFC2NMR0sCkRsM#H0sMHoR#C
Lo
HMRVRHR25LRC0EMR
RRCRs0Mks52"";R
RCCD#
RRRR0sCk5sM"kBFDM8RFH0RlCbDl0CMRFADO)	RqRv3Q0#REsCRCRN8Ns88CR##sHCo#s0CCk8R#oHMRC0ERl#NCDROFRO	N0#RE)CRq"v?2R;
R8CMR;HV
8CMRMVkOM_HH
0;VOkM0MHFR0oC_8CM_b8C0#E5HRxC:MRH0CCosRR;80CbERR:HCM0o2CsR0sCkRsMHCM0oRCsHP#
NNsHLRDCl_HM#CHxRH:RMo0CC:sR=;Rj
oLCHRM
RMlH_x#HC=R:Rb8C0
E;RVRHRH5#x<CRRb8C0RE20MEC
RRRRMlH_x#HC=R:Rx#HCR;
R8CMR;HV
sRRCs0kMHRlMH_#x
C;CRM8o_C0C_M880CbEN;
0H0sLCk0RMoCC0sNFss_CsbF0RR:#H0sM
o;Ns00H0LkCCRoMNCs0_FssFCbsF0RVDRLF_O	sRNl:sRNO0EHCkO0sHCR#kRVMHO_M5H0s8N8sC_so
2;-L-RCMoHRFLDOs	RNHlRlCbDl0CMNF0HMHR#oDMN#$
0bHCRMN0_s$sNRRH#NNss$jR5RR0F6F2RVMRH0CCosO;
F0M#NRM0I0H8Es_NsRN$:MRH0s_NsRN$:5=R4.,R,,RcRRg,4RU,d;n2
MOF#M0N0CR8b_0ENNss$RR:H_M0NNss$=R:Rn54d,UcRgU4.c,Rj,gnRc.jU4,Rj,.cR.642O;
F0M#NRM08dHP.RR:HCM0oRCs:5=RI0H8E2-4/;dn
MOF#M0N0HR8PR4n:MRH0CCos=R:RH5I8-0E442/UO;
F0M#NRM08UHPRH:RMo0CC:sR=IR5HE80-/42gO;
F0M#NRM08cHPRH:RMo0CC:sR=IR5HE80-/42cO;
F0M#NRM08.HPRH:RMo0CC:sR=IR5HE80-/42.O;
F0M#NRM084HPRH:RMo0CC:sR=IR5HE80-/424
;
O#FM00NMRFLFD:4RRFLFDMCNRR:=5P8H4RR>j
2;O#FM00NMRFLFD:.RRFLFDMCNRR:=5P8H.RR>j
2;O#FM00NMRFLFD:cRRFLFDMCNRR:=5P8HcRR>j
2;O#FM00NMRFLFD:URRFLFDMCNRR:=5P8HURR>j
2;O#FM00NMRFLFDR4n:FRLFNDCM=R:RH58PR4n>2Rj;F
OMN#0ML0RFdFD.RR:LDFFCRNM:5=R8dHP.RR>j
2;
MOF#M0N0HR8Pd4nU:cRR0HMCsoCRR:=5b8C04E-2n/4d;Uc
MOF#M0N0HR8PgU4.RR:HCM0oRCs:5=R80CbE2-4/gU4.O;
F0M#NRM08cHPjRgn:MRH0CCos=R:RC58b-0E4c2/j;gn
MOF#M0N0HR8Pc.jURR:HCM0oRCs:5=R80CbE2-4/c.jUO;
F0M#NRM084HPjR.c:MRH0CCos=R:RC58b-0E442/j;.c
MOF#M0N0HR8P.64RH:RMo0CC:sR=8R5CEb0-/426;4.
F
OMN#0ML0RF6FD4:.RRFLFDMCNRR:=5P8H6R4.>2Rj;F
OMN#0ML0RF4FDjR.c:FRLFNDCM=R:RH58P.4jcRR>j
2;O#FM00NMRFLFDc.jURR:LDFFCRNM:5=R8.HPjRcU>2Rj;F
OMN#0ML0RFcFDjRgn:FRLFNDCM=R:RH58PgcjnRR>j
2;O#FM00NMRFLFDgU4.RR:LDFFCRNM:5=R8UHP4Rg.>2Rj;F
OMN#0ML0RF4FDncdURL:RFCFDN:MR=8R5HnP4dRUc>2Rj;O

F0M#NRM0#_klI0H8ERR:HCM0oRCs:A=Rm mpqbh'FL#5F4FD2RR+Apmm 'qhb5F#LDFF.+2RRmAmph q'#bF5FLFDRc2+mRAmqp hF'b#F5LF2DURA+Rm mpqbh'FL#5F4FDn
2;O#FM00NMRl#k_b8C0:ERR0HMCsoCRR:=6RR-5mAmph q'#bF5FLFD.642RR+Apmm 'qhb5F#LDFF4cj.2RR+Apmm 'qhb5F#LDFF.Ujc2RR+Apmm 'qhb5F#LDFFcnjg2RR+Apmm 'qhb5F#LDFFU.4g2
2;
MOF#M0N0_RIOHEFOIC_HE80RH:RMo0CC:sR=HRI8_0ENNss$k5#lH_I820E;F
OMN#0MI0R_FOEH_OC80CbERR:HCM0oRCs:8=RCEb0_sNsN#$5kIl_HE802O;
F0M#NRM08E_OFCHO_8IH0:ERR0HMCsoCRR:=I0H8Es_Ns5N$#_kl80CbE
2;O#FM00NMRO8_EOFHCC_8bR0E:MRH0CCos=R:Rb8C0NE_s$sN5l#k_b8C0;E2
F
OMN#0MI0R_8IH0ME_kOl_C#DDRH:RMo0CC:sR=IR5HE80-/42IE_OFCHO_8IH0+ERR
4;O#FM00NMR8I_CEb0_lMk_DOCD:#RR0HMCsoCRR:=5b8C04E-2_/IOHEFO8C_CEb0R4+R;O

F0M#NRM08H_I8_0EM_klODCD#RR:HCM0oRCs:5=RI0H8E2-4/O8_EOFHCH_I8R0E+;R4
MOF#M0N0_R880CbEk_MlC_ODRD#:MRH0CCos=R:RC58b-0E482/_FOEH_OC80CbERR+4
;
O#FM00NMR#I_HRxC:MRH0CCos=R:RII_HE80_lMk_DOCD*#RR8I_CEb0_lMk_DOCD
#;O#FM00NMR#8_HRxC:MRH0CCos=R:RI8_HE80_lMk_DOCD*#RR88_CEb0_lMk_DOCD
#;
MOF#M0N0FRLF8D_RL:RFCFDN:MR=8R5_x#HCRR-IH_#x<CR=2Rj;F
OMN#0ML0RF_FDIRR:LDFFCRNM:M=RFL05F_FD8
2;
MOF#M0N0EROFCHO_8IH0:ERR0HMCsoCRR:=5mAmph q'#bF5FLFD2_8R8*R_FOEH_OCI0H8E+2RRm5Amqp hF'b#F5LFID_2RR*IE_OFCHO_8IH0;E2
MOF#M0N0EROFCHO_b8C0:ERR0HMCsoCRR:=5mAmph q'#bF5FLFD2_8R8*R_FOEH_OC80CbE+2RRm5Amqp hF'b#F5LFID_2RR*IE_OFCHO_b8C0;E2
MOF#M0N0HRI8_0EM_klODCD#RR:HCM0oRCs:5=RApmm 'qhb5F#LDFF_R82*H5I8-0E482/_FOEH_OCI0H8E+2RRm5Amqp hF'b#F5LFID_2RR*58IH04E-2_/IOHEFOIC_HE802RR+4O;
F0M#NRM080CbEk_MlC_ODRD#:MRH0CCos=R:Rm5Amqp hF'b#F5LF8D_25R*80CbE2-4/O8_EOFHCC_8b20ER5+RApmm 'qhb5F#LDFF_RI2*8R5CEb0-/42IE_OFCHO_b8C0RE2+;R4
b0$CkRF0k_L#04_$RbCHN#Rs$sNRC58b_0EM_klODCD#R-48MFI0jFR,HRI8_0EM_klODCD#R-48MFI0jFR2VRFR8#0_oDFH
O;#MHoNsDRF_k0L4k#RF:RkL0_k_#40C$b;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFVsF_8k50RHkMb0FR0RH0s-N#002C#
o#HMRNDI0Fk_#Lk4RR:F_k0L4k#_b0$C0;
$RbCF_k0L.k#_b0$C#RHRsNsN5$R80CbEk_MlC_OD-D#4FR8IFM0RRj,.H*I8_0EM_klODCD#R+48MFI0jFR2VRFR8#0_oDFH
O;#MHoNsDRF_k0L.k#RF:RkL0_k_#.0C$b;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFVsF_8k50RHkMb0FR0RH0s-N#002C#
o#HMRNDI0Fk_#Lk.RR:F_k0L.k#_b0$C0;
$RbCF_k0Lck#_b0$C#RHRsNsN5$R80CbEk_MlC_OD-D#4FR8IFM0RRj,cH*I8_0EM_klODCD#R+d8MFI0jFR2VRFR8#0_oDFH
O;#MHoNsDRF_k0Lck#RF:RkL0_k_#c0C$b;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFVsF_8k50RHkMb0FR0RH0s-N#002C#
o#HMRNDI0Fk_#LkcRR:F_k0Lck#_b0$C0;
$RbCF_k0LUk#_b0$C#RHRsNsN5$R80CbEk_MlC_OD-D#4FR8IFM0RRj,UH*I8_0EM_klODCD#R+(8MFI0jFR2VRFR8#0_oDFH
O;#MHoNsDRF_k0LUk#RF:RkL0_k_#U0C$b;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFVsF_8k50RHkMb0FR0RH0s-N#002C#
o#HMRNDI0Fk_#LkURR:F_k0LUk#_b0$C0;
$RbCbHNs0L$_k_#U0C$bRRH#NNss$8R5CEb0_lMk_DOCD4#-RI8FMR0FjI,RHE80_lMk_DOCD4#-RI8FMR0FjF2RV0R#8F_Do;HO
o#HMRNDssbNH_0$LUk#Rb:RN0sH$k_L#0U_$;bCRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFR8s_FRk05bHMk00RFsR0H0-#N#0C2H
#oDMNRNIbs$H0_#LkURR:bHNs0L$_k_#U0C$b;$
0bFCRkL0_kn#4_b0$C#RHRsNsN5$R80CbEk_MlC_OD-D#4FR8IFM0RRj,4In*HE80_lMk_DOCD4#+6FR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNRksF0k_L#R4n:kRF0k_L#_4n0C$b;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RV_Rs80FkRM5HbRk000FRs#H-0CN0##2
HNoMDFRIkL0_kn#4RF:RkL0_kn#4_b0$C0;
$RbCbHNs0L$_kn#4_b0$C#RHRsNsN5$R80CbEk_MlC_OD-D#4FR8IFM0RRj,.H*I8_0EM_klODCD#R+48MFI0jFR2VRFR8#0_oDFH
O;#MHoNsDRbHNs0L$_kn#4Rb:RN0sH$k_L#_4n0C$b;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFVsF_8k50RHkMb0FR0RH0s-N#002C#
o#HMRNDIsbNH_0$L4k#nRR:bHNs0L$_kn#4_b0$C0;
$RbCF_k0Ldk#.$_0bHCR#sRNsRN$5b8C0ME_kOl_C#DD-84RF0IMF,RjR*d.I0H8Ek_MlC_OD+D#d84RF0IMF2RjRRFV#_08DHFoO#;
HNoMDFRskL0_k.#dRF:RkL0_k.#d_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$FsVR_k8F0HR5M0bkRR0F0-sH#00NC
#2#MHoNIDRF_k0Ldk#.RR:F_k0Ldk#.$_0b
C;0C$bRsbNH_0$Ldk#.$_0bHCR#sRNsRN$5b8C0ME_kOl_C#DD-84RF0IMF,RjRIc*HE80_lMk_DOCDd#+RI8FMR0FjF2RV0R#8F_Do;HO
o#HMRNDssbNH_0$Ldk#.RR:bHNs0L$_k.#d_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFR8s_FRk05bHMk00RFsR0H0-#N#0C2H
#oDMNRNIbs$H0_#Lkd:.RRsbNH_0$Ldk#.$_0b
C;#MHoNsDRF_k0C:MRR8#0_oDFHPO_CFO0sC58b_0EM_klODCD#R-48MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-MRCNCLD#FRVssR0H0-#N#0C
o#HMRNDI0Fk_RCM:0R#8F_Do_HOP0COF8s5CEb0_lMk_DOCD4#-RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-C-RMDNLCV#RF0sRs#H-0CN0#H
#oDMNR0Is_RCM:0R#8F_Do_HOP0COF8s5CEb0_lMk_DOCD4#-RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-I-RsCH0RNCML#DCRsVFROCNEFRsIVRFRv)qRDOCD##
HNoMDMRH_osCR#:R0D8_FOoH_OPC05FsI0H8E6+dRI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RCk#8FR0RosCHC#0sQR7h#R
HNoMDFRsks0_C:oRR8#0_oDFHPO_CFO0sH5I8+0Ed86RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-#RkC08RFCRso0H#C7sRm
za#MHoNIDRF_k0sRCo:0R#8F_Do_HOP0COFIs5HE80+Rd68MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-k-R#RC80sFRC#oH0RCs7amz
o#HMRNDs0Fk_osC4RR:#_08DHFoOC_POs0F58IH04E-RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-k-R#RC80OFRE#FFCCRL0CICMQR7hMRN8kRF00bkRRFVAODF	qR)vH
#oDMNR8sN_osCR#:R0D8_FOoH_OPC05FsNs88I0H8ER-48MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--k8#CRR0FsHCo#s0CR7)q7#)
HNoMDNRI8C_soRR:#_08DHFoOC_POs0F58N8s8IH04E-RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RCk#8FR0RosCHC#0sqRW7
7)#MHoNDDRFsI_Ns88R#:R0D8_FOoH_OPC05Fs48dRF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-s-RNs88R0LH#MRHbRk00)FRqOvRC#DDRR5cL#H0RJsCkCHs8#2
HNoMDFRDIN_I8R8s:0R#8F_Do_HOP0COF4s5dFR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-NRI8R8sL#H0RbHMk00RFqR)vCRODRD#5LcRHR0#skCJH8sC2H
#oDMNR7)q70)_l:bRR8#0_oDFHPO_CFO0s85N8HsI8-0E4FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-#RkC08RFHRbbHCDM)CRq)77
o#HMRNDW7q7)l_0bRR:#_08DHFoOC_POs0F58N8s8IH04E-RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RCk#8FR0RbbHCMDHCqRW7
7)#MHoN7DRQ0h_l:bRR8#0_oDFHPO_CFO0sH5I8-0E4FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--k8#CRR0FbCHbDCHMRh7Q
o#HMRNDW0 _l:bRR8#0_oDFHRO;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RCk#8FR0RbbHCMDHC RW
R--CRM8LODF	NRsllRHblDCCNM00MHFRo#HM#ND
R--LHCoMCR#D0CORlsNRbHlDCClM00NHRFM#MHoN
D#VOkM0MHFR0oC_lMk_5nc80CbEH:RMo0CCRs2skC0sHMRMo0CCHsR#N
PsLHNDPCRN:DRR0HMCsoCRR:=jL;
CMoH
PRRN:DR=CR8b/0En
c;RVRHR855CEb0R8lFR2ncRc>RU02RE
CMRRRRPRND:P=RN+DRR
4;RMRC8VRH;R
RskC0sPMRN
D;CRM8o_C0M_kln
c;VOkM0MHFR0oC_VDC0CFPs._d5b8C0:ERR0HMCsoC2CRs0MksR0HMCsoCR
H#LHCoMR
RskC0s8M5CEb0R8lFR2nc;M
C8CRo0C_DVP0FCds_.V;
k0MOHRFMo_C0D0CVFsPC5b8C0:ERR0HMCsoC;NRlGRR:HCM0o2CsR0sCkRsMHCM0oRCsHP#
NNsHLRDCPRND:MRH0CCos=R:R
j;LHCoMR
RH5VR80CbERR-lRNG>j=R2ER0CRM
RPRRN:DR=CR8bR0E-NRlGR;
R#CDCR
RRNRPD=R:Rb8C0
E;RMRC8VRH;R
RskC0sPM5N;D2
8CMR0oC_VDC0CFPsV;
k0MOHRFMo_C0M_kld8.5CEb0RH:RMo0CCRs2skC0sHMRMo0CCHsR#N
PsLHNDPCRN:DRR0HMCsoCRR:=jL;
CMoH
HRRV8R5CEb0RR<=cNURM88RCEb0R4>Rn02RE
CMRRRRRDPNRR:=4R;
R8CMR;HV
sRRCs0kMNRPDC;
Mo8RCM0_kdl_.V;
k0MOHRFMo_C0M_kl48n5CEb0RH:RMo0CCRs2skC0sHMRMo0CCHsR#N
PsLHNDPCRN:DRR0HMCsoCRR:=jL;
CMoH
HRRV8R5CEb0RR<=4NnRM88RCEb0Rj>R2ER0CRM
RRRRPRND:4=R;R
RCRM8H
V;RCRs0MksRDPN;M
C8CRo0k_Mln_4;F
OMN#0MM0RkOl_C_DDn:cRR0HMCsoCRR:=o_C0M_kln8c5CEb02O;
F0M#NRM0D0CVFsPC_Rd.:MRH0CCos=R:R0oC_VDC0CFPs._d5b8C0;E2
MOF#M0N0kRMlC_ODdD_.RR:HCM0oRCs:o=RCM0_kdl_.C5DVP0FCds_.
2;O#FM00NMRVDC0CFPsn_4RH:RMo0CC:sR=CRo0C_DVP0FCDs5CFV0P_CsdR.,d;.2
MOF#M0N0kRMlC_OD4D_nRR:HCM0oRCs:o=RCM0_k4l_nC5DVP0FC4s_n
2;
b0$CkRF0k_L#$_0bnC_cH#R#sRNsRN$5lMk_DOCDc_nRI8FMR0FjI,RHE80-84RF0IMF2RjRRFV#_08DHFoO0;
$RbCF_k0L_k#0C$b_#d.RRH#NNss$MR5kOl_C_DDd8.RF0IMF,RjR8IH04E-RI8FMR0FjF2RV0R#8F_Do;HO
b0$CkRF0k_L#$_0b4C_nH#R#sRNsRN$5lMk_DOCDn_4RI8FMR0FjI,RHE80-84RF0IMF2RjRRFV#_08DHFoO#;
HNoMDFRskL0_kn#_c:#RR0Fk_#Lk_b0$Cc_n#R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFRk8F0HR5M0bkRR0F0-sH#00NC
#2#MHoNIDRF_k0L_k#nRc#:kRF0k_L#$_0bnC_cR#;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RVFR8k50RHkMb0FR0RH0s-N#002C#
o#HMRNDs0Fk_#Lk_#d.RF:RkL0_k0#_$_bCd;.#RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$F8VRFRk05bHMk00RFsR0H0-#N#0C2H
#oDMNRkIF0k_L#._d#RR:F_k0L_k#0C$b_#d.;H
#oDMNRksF0k_L#n_4#RR:F_k0L_k#0C$b_#4n;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFV80FkRM5HbRk000FRs#H-0CN0##2
HNoMDFRIkL0_k4#_n:#RR0Fk_#Lk_b0$Cn_4##;
HNoMDFRskC0_MR_#:0R#8F_Do_HOP0COFMs5kOl_C_DDn8cRF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RNCML#DCRsVFRH0s-N#00
C##MHoNIDRF_k0C#M_R#:R0D8_FOoH_OPC05FsM_klODCD_Rnc8MFI0jFR2#;
HNoMDFRskC0_M._dR#:R0D8_FOoH;H
#oDMNRkIF0M_C_Rd.:0R#8F_Do;HO
o#HMRNDs0Fk__CM4:nRR8#0_oDFH
O;#MHoNIDRF_k0C4M_nRR:#_08DHFoO#;
HNoMDsRI0M_C_:#RR8#0_oDFHPO_CFO0sk5MlC_ODnD_cFR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--I0sHCMRCNCLD#FRVsNRCOsERFFIRVqR)vCROD
D##MHoNIDRsC0_M._dR#:R0D8_FOoH;H
#oDMNR0Is__CM4:nRR8#0_oDFH
O;#MHoNHDRMC_soR_#:0R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-k-R#RC80sFRC#oH0RCs7RQh
o#HMRNDs0Fk_osC_:#RR8#0_oDFHPO_CFO0sH5I8-0E4FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RCk#8FR0RosCHC#0smR7z#a
HNoMDFRIks0_C#o_R#:R0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2R;RRH
#oDMNR8sN_osC_:#RR8#0_oDFHPO_CFO0s85N8HsI8-0E4FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-#RkC08RFCRso0H#CqsR7
7)#MHoNIDRNs8_C#o_R#:R0D8_FOoH_OPC05FsNs88I0H8ER-48MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--k8#CRR0FsHCo#s0CR7q7)H
#oDMNRIDF_8sN8#s_R#:R0D8_FOoH_OPC05Fs6FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-8RN8LsRHR0#HkMb0FR0Rv)qRDOCD5#RcHRL0s#RCHJks2C8
o#HMRNDD_FII8N8sR_#:0R#8F_Do_HOP0COF6s5RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-R8N8sHRL0H#RM0bkRR0F)RqvODCD#cR5R0LH#CRsJskHC
82-C-RM#8RCODC0NRsllRHblDCCNM00MHFRo#HM#ND
0N0skHL0\CR3lsN_VFV#\C0R#:R0MsHo
;
LHCoMR
Rz:cdRRHV58sN8ss_CRo2oCCMsCN0RR--oCCMsCN0RFLDOs	RNRl
R-RR-VRQR8N8s8IH0<ERRFOEH_OCI0H8E#RN#MHoR''jRR0Fk#MkCL8RH
0#RRRRzRjR:VRHR85N8HsI8R0E=2R4RMoCC0sNCR
SRDRRFsI_Ns88RR<="jjjjjjjjjjjjRj"&NRs8C_so25j;R
SRDRRFII_Ns88RR<="jjjjjjjjjjjjRj"&NRI8C_so25j;C
SMo8RCsMCNR0Cz
j;RRRRzR4R:VRHR85N8HsI8R0E=2R.RMoCC0sNCS
SD_FIs8N8s=R<Rj"jjjjjjjjjjRj"&NRs8C_soR548MFI0jFR2S;
RRRRD_FII8N8s=R<Rj"jjjjjjjjjjRj"&NRI8C_soR548MFI0jFR2S;
CRM8oCCMsCN0R;z4
RRRRRz.RH:RVNR58I8sHE80Rd=R2CRoMNCs0SC
SIDF_8sN8<sR=jR"jjjjjjjjjRj"&NRs8C_soR5.8MFI0jFR2S;
RRRRD_FII8N8s=R<Rj"jjjjjjjjjj&"RR8IN_osC58.RF0IMF2Rj;C
SMo8RCsMCNR0Cz
.;RRRRzRdR:VRHR85N8HsI8R0E=2RcRMoCC0sNCS
SD_FIs8N8s=R<Rj"jjjjjjjjj"RR&s_N8s5CodFR8IFM0R;j2
RSRRFRDIN_I8R8s<"=RjjjjjjjjjRj"&NRI8C_soR5d8MFI0jFR2S;
CRM8oCCMsCN0R;zd
RRRRRzcRH:RVNR58I8sHE80R6=R2CRoMNCs0SC
RRRRD_FIs8N8s=R<Rj"jjjjjj"jjRs&RNs8_Cco5RI8FMR0Fj
2;SRRRRIDF_8IN8<sR=jR"jjjjjjjj"RR&I_N8s5CocFR8IFM0R;j2
MSC8CRoMNCs0zCRcR;
RzRR6:RRRRHV58N8s8IH0=ERRRn2oCCMsCN0
RSRRFRDIN_s8R8s<"=Rjjjjjjjj"RR&s_N8s5Co6FR8IFM0R;j2
DSSFII_Ns88RR<="jjjjjjjj&"RR8IN_osC586RF0IMF2Rj;C
SMo8RCsMCNR0Cz
6;RRRRzRnR:VRHR85N8HsI8R0E=2R(RMoCC0sNCR
SRDRRFsI_Ns88RR<="jjjjjjj"RR&s_N8s5ConFR8IFM0R;j2
DSSFII_Ns88RR<="jjjjjjj"RR&I_N8s5ConFR8IFM0R;j2
MSC8CRoMNCs0zCRnR;
RzRR(:RRRRHV58N8s8IH0=ERRRU2oCCMsCN0
RSRRFRDIN_s8R8s<"=RjjjjjRj"&NRs8C_soR5(8MFI0jFR2S;
SIDF_8IN8<sR=jR"jjjjj&"RR8IN_osC58(RF0IMF2Rj;C
SMo8RCsMCNR0Cz
(;RRRRzRUR:VRHR85N8HsI8R0E=2RgRMoCC0sNCR
SRDRRFsI_Ns88RR<="jjjjRj"&NRs8C_soR5U8MFI0jFR2S;
SIDF_8IN8<sR=jR"jjjj"RR&I_N8s5CoUFR8IFM0R;j2
MSC8CRoMNCs0zCRUR;
RzRRg:RRRRHV58N8s8IH0=ERR24jRMoCC0sNCR
SRDRRFsI_Ns88RR<="jjjj&"RR8sN_osC58gRF0IMF2Rj;S
SD_FII8N8s=R<Rj"jjRj"&NRI8C_soR5g8MFI0jFR2S;
CRM8oCCMsCN0R;zg
RRRRjz4RRR:H5VRNs88I0H8ERR=4R42oCCMsCN0
RSRRFRDIN_s8R8s<"=Rj"jjRs&RNs8_C4o5jFR8IFM0R;j2
DSSFII_Ns88RR<="jjj"RR&I_N8s5Co48jRF0IMF2Rj;C
SMo8RCsMCNR0Cz;4j
RRRR4z4RRR:H5VRNs88I0H8ERR=4R.2oCCMsCN0
RSRRFRDIN_s8R8s<"=RjRj"&NRs8C_so454RI8FMR0Fj
2;SFSDIN_I8R8s<"=RjRj"&NRI8C_so454RI8FMR0Fj
2;S8CMRMoCC0sNC4Rz4R;
RzRR4R.R:VRHR85N8HsI8R0E=dR42CRoMNCs0SC
RRRRD_FIs8N8s=R<R''jRs&RNs8_C4o5.FR8IFM0R;j2
DSSFII_Ns88RR<='Rj'&NRI8C_so.54RI8FMR0Fj
2;S8CMRMoCC0sNC4Rz.R;
RzRR4RdR:VRHR85N8HsI8R0E>dR42CRoMNCs0SC
RRRRD_FIs8N8s=R<R8sN_osC5R4d8MFI0jFR2S;
RRRRD_FII8N8s=R<R8IN_osC5R4d8MFI0jFR2S;
CRM8oCCMsCN0Rdz4;R

R-RR-VRQRH58MC_sos2RC#oH0RCs7RQhkM#HopRBiR
RR4Rzc:RRRRHV5M8H_osC2CRoMNCs0RC
RRRRRbRRsCFO#5#RB,piRh7Q2CRLo
HMRRRRRRRRRRRRH5VRBRpi=4R''MRN8pRBiP'CC2M0RC0EMR
RRRRRRRRRRRRRRMRH_osCRR<=5j"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjRj"&QR7h
2;RRRRRRRRRRRRCRM8H
V;RRRRRRRRCRM8bOsFC;##
MSC8CRoMNCs0zCR4
c;RRRRzR46RH:RVMR5F80RHsM_CRo2oCCMsCN0
RRRRRRRRRRRR_HMsRCo<5=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj&"RRh7Q2S;
CRM8oCCMsCN0R6z4;R

R-RR-VRQR85sF_k0s2CoRosCHC#0s_R)7amzRHk#M)oR_pmBiR
RR4RznFs8kR0R:VRHR85sF_k0s2CoRMoCC0sNCR
RRRRRRsRbF#OC#)R5_pmBis,RF_k0s2CoRoLCHRM
RRRRRRRRRHRRV)R5_pmBiRR='R4'NRM8)B_mpCi'P0CM2ER0CRM
RRRRRRRRRRRRR)RR_z7ma=R<RksF0C_so
4;RRRRRRRRRRRRCRM8H
V;RRRRRRRRCRM8bOsFC;##
RRRRRRRR8CMRMoCC0sNC4RznFs8k
0;RRRRzs4(80FkRRR:H5VRMRF0sk8F0C_soo2RCsMCN
0CRRRRRRRRRRRR)m_7z<aR=FRsks0_C;o4
MSC8CRoMNCs0zCR48(sF;k0
z
S48nIFRk0RH:RVIR580Fk_osC2CRoMNCs0RC
RRRRRbRRsCFO#5#RWB_mpRi,I0Fk_osC2CRLo
HMRRRRRRRRRRRRH5VRWB_mp=iRR''4R8NMRmW_B'piCMPC002RE
CMRRRRRRRRRRRRRRRRWm_7z<aR=FRIks0_CIo5HE80-84RF0IMF2Rj;R
RRRRRRRRRRMRC8VRH;R
RRRRRRMRC8sRbF#OC#R;
RRRRRCRRMo8RCsMCNR0CzI4n80Fk;R
RR4Rz(FI8kR0R:VRHRF5M08RIF_k0s2CoRMoCC0sNCR
RRRRRRRRRR_RW7amzRR<=I0Fk_osC58IH04E-RI8FMR0Fj
2;S8CMRMoCC0sNC4Rz(FI8k
0;
RRRRR--Q5VRs8N8sC_sos2RC#oH0RCs)7q7)#RkHRMomiBp
RRRRnz4s:RRRRHV58sN8ss_CRo2oCCMsCN0
R--RRRRRbRRsCFO#5#RmiBp,qR)727)RoLCH-M
-RRRRRRRRRRRRRHV5pmBiRR='R4'NRM8miBp'CCPMR020MEC
R--RRRRRRRRRRRRRsRRNs8_C<oR=qR)757)Ns88I0H8ER-48MFI0jFR2-;
-RRRRRRRRRRRR8CMR;HV
R--RRRRRCRRMb8RsCFO#
#;-C-SMo8RCsMCNR0Czs4n;-
-RRRRzs4(RH:RVMR5Fs0RNs88_osC2CRoMNCs0RC
RRRRRRRRRsRRNs8_C<oR=qR)7;7)
MSC8CRoMNCs0zCR4;ns
-
S-VRQRN5I8_8ss2CoRosCHC#0sqRW7R7)kM#Ho_RWmiBp
RRRRnz4I:RRRRHV58IN8ss_CRo2oCCMsCN0
RRRRRRRRFbsO#C#Rp5BiW,Rq)772CRLo
HMRRRRRRRRRRRRH5VRBRpi=4R''MRN8pRBiP'CC2M0RC0EMR
RRRRRRRRRRRRRRNRI8C_so=R<R7Wq7N)58I8sHE80-84RF0IMF2Rj;R
RRRRRRRRRRMRC8VRH;R
RRRRRRMRC8sRbF#OC#S;
CRM8oCCMsCN0Rnz4IR;
RzRR4R(I:VRHRF5M0NRI8_8ss2CoRMoCC0sNCR
RRRRRRRRRRNRI8C_so=R<R7Wq7
);S8CMRMoCC0sNC4Rz(
I;
RRRRR-- sG0NFRDoRHOVRFs7DkNRsbF0NRO#SC
zosCRb:RsCFO#B#5pRi2LHCoMR
SRRHV5iBp'  ehNaRMB8Rp=iRR''42ER0CSM
R7RRQ0h_l<bR=QR7hS;
R)RRq)77_b0lRR<=)7q7)S;
RWRRq)77_b0lRR<=W7q7)S;
RWRR l_0b=R<R;W 
RSRCRM8H
V;S8CMRFbsO#C#;S

-Q-RVCR)Nq8R8C8s#=#RRHWs0qCR8C8s#R#,LN$b#7#RQ0hRFkRF00bkRRHVWH R#MRCNCLD8z
SlRkG:sRbF#OC# 5W_b0l,qR)7_7)0,lbR7Wq70)_lRb,7_Qh0,lbRksF0C_soS2
RCRLo
HMSRRRRRHV57Wq70)_l=bRR7)q70)_lNbRMW8R l_0bRR='24'RC0EMS
SRFRsks0_CRo4<7=RQ0h_l
b;SDSC#SC
SsRRF_k0s4CoRR<=s0Fk_osC58IH04E-RI8FMR0Fj
2;SMSC8VRH;C
SMb8RsCFO#
#;SRRRRR
RR-R-RMtCC0sNCER0CqR)vCRODRD#NRM8#CCDOD0RFOoHRsVFRv)qA_4n114_4z
S4:URRRHV5FOEH_OCI0H8ERR=4o2RCsMCN
0CRRRRSgz4RV:RFHsRRRHM5b8C0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CSR--Q5VRNs88I0H8ERR>4Rc2M8CCRR0FONsC0ICRsCH0RNCMLRDCNRM8Fbk0kC0RMDNLCCR#D0CORoDFHRO
RRRRRSRRzR.j:VRHR85N8HsI8R0E>cR42CRoMNCs0SC
-V-RHVGRFOsRNRDD4UdU(#,RCODC0VRFRH0s#00NCFRM0CRLHRMosHCo#s0CCS8
SsSSF_k0CHM52=R<R''4RCIEM)R5q)77_b0l58N8s8IH04E-RI8FMR0F4Rc2=2RHR#CDCjR''S;
SISSF_k0CHM52=R<R''4RCIEMIR5Ns8_CNo58I8sHE80-84RF0IMFcR42RR=HC2RDR#C';j'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RWRCIEMIR5Ns8_CNo58I8sHE80-84RF0IMFcR42RR=HC2RDR#C';j'
RRRRRRRRMSC8CRoMNCs0zCR.
j;SR--Q5VRNs88I0H8E=R<R24cRRMFI0sHCMRCNCLDRRFsFbk0kC0RMDNLCCR#D0CORoDFHMORCCC88S
RRRRRS4z.RH:RVNR58I8sHE80RR<=4Rc2oCCMsCN0
SSSSksF0M_C5RH2<'=R4
';SSSSI0Fk_5CMH<2R=4R''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=W
 ;RRRRRRRRS8CMRMoCC0sNC.Rz4S;
-t-RCsMCNR0C0REC)RqvODCD#MRN8sR0H0-#N#0C
RRRRRRRR.Sz.RR:VRFs[MRHRH5I8_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
RRRRRRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVAv)q_d4nU4cX7RR:DCNLD#RHR""W;R
RRRRRRRRRRRRRRCRLo
HMRRRRRRRRRRRRSqA)vn_4dXUc4:7RRv)qA_4n114_4R
SRRRRRRRRRbRRFRs0lRNb5q7Q5Rj2=H>RMC_so25[,7Rq7R)q=D>RFII_Ns885R4d8MFI0jFR27,RQ=AR>jR""q,R7A7)RR=>D_FIs8N8sd54RI8FMR0Fj
2,SSSS Rhq='>R4R',1q1)RR=>',j'RqW RR=>I_s0CHM52B,RpRiq=B>RpRi, RhA='>R4R',1A1)RR=>',j'RAW RR=>',j'RiBpA>R=RiBp,S
SSRRRRq7m5Rj2=I>RF_k0L4k#5[H,27,RmjA52>R=RksF0k_L#H45,2[2;R

RRRRRRRRRRRRRsRRF_k0s5Co[<2R=FRskL0_k5#4H2,[RCIEMsR5F_k0CHM52RR='24'R#CDCZR''S;
SISSF_k0s5Co[<2R=FRIkL0_k5#4H2,KRCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRSRRCRM8oCCMsCN0R.z.;R
RRSRRCRM8oCCMsCN0Rgz4;R
RRMRC8CRoMNCs0zCR4RU;R
RRRRRRRRR
R-RR-CRtMNCs00CRE)CRqOvRC#DDR8NMRD#CCRO0DHFoOFRVsqR)vnA4__1.1S.
zR.d:VRHRE5OFCHO_8IH0=ERRR.2oCCMsCN0
RRRR.SzcRR:VRFsHMRHRC58b_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
-S-RRQV58N8s8IH0>ERR24dRCMC8FR0RCOsNR0CI0sHCMRCNCLDR8NMR0FkbRk0CLMND#CRCODC0FRDo
HORRRRRRRRS6z.RH:RVNR58I8sHE80R4>Rdo2RCsMCN
0CSR--VRHGVRFsODNDRU4dUR(,#CCDOF0RVsR0HN#00MCRFL0RCoHMRosCHC#0s
C8RRRRRRRRRRRRRRRRs0Fk_5CMH<2R=4R''ERIC5MR)7q7)l_0b85N8HsI8-0E4FR8IFM0R24dRH=R2DRC#'CRj
';SSSSI0Fk_5CMH<2R=4R''ERIC5MRI_N8s5CoNs88I0H8ER-48MFI04FRd=2RRRH2CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R ERIC5MRI_N8s5CoNs88I0H8ER-48MFI04FRd=2RRRH2CCD#R''j;R
RRRRRRCRSMo8RCsMCNR0Cz;.6
-S-RRQV58N8s8IH0<ER=dR42FRMRHIs0CCRMDNLCsRFR0FkbRk0CLMND#CRCODC0FRDoRHOM8CCCR8
SRRRR.SznRR:H5VRNs88I0H8E=R<R24dRMoCC0sNCR
SRRRRRRRRRsRRF_k0CHM52=R<R''4;S
SSFSIkC0_M25HRR<=';4'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RW;R
RRRRRRCRSMo8RCsMCNR0Cz;.n
-S-RMtCC0sNCER0CqR)vCRODRD#NRM80-sH#00NCR#
RRRRRSRRzR.(:FRVsRR[H5MRI0H8Ek_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0RC
RRRRRRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)RAqUv_4Xg..:7RRLDNCHDR#WR""R;
RRRRRRRRRRRRRLRRCMoH
RRRRRRRRRRRR)SAqUv_4Xg..:7RRv)qA_4n11._.R
SRRRRRRRRRbRRFRs0lRNb5q7QRR=>HsM_C.o5*4[+RI8FMR0F.2*[,7Rq7R)q=D>RFII_Ns885R4.8MFI0jFR27,RQ=AR>jR"jR",q)77A>R=RIDF_8sN84s5.FR8IFM0R,j2
SSSRRRR Rhq='>R4R',1q1)RR=>',j'RqW RR=>I_s0CHM52B,RpRiq=B>RpRi, RhA='>R4R',1A1)RR=>',j'RAW RR=>',j'RiBpA>R=RiBp,S
SSRRRRq7m5R42=I>RF_k0L.k#5.H,*4[+27,Rmjq52>R=RkIF0k_L#H.5,[.*27,Rm4A52>R=RksF0k_L#H.5,[.*+,42RA7m5Rj2=s>RF_k0L.k#5RH,.2*[2R;
RRRRRRRRRRRRRsRRF_k0s5Co.2*[RR<=s0Fk_#Lk.,5H.2*[RCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRsRRF_k0s5Co.+*[4<2R=FRskL0_k5#.H*,.[2+4RCIEMsR5F_k0CHM52RR='24'R#CDCZR''S;
SISSF_k0s5Co.2*[RR<=I0Fk_#Lk.,5H.2*[RCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRIRRF_k0s5Co.+*[4<2R=FRIkL0_k5#.H*,.[2+4RCIEMIR5F_k0CHM52RR='24'R#CDCZR''
;
RRRRRRRRS8CMRMoCC0sNC.Rz(R;
RRRRS8CMRMoCC0sNC.RzcR;
RCRRMo8RCsMCNR0Cz;.dR
R
SRRRRR--tCCMsCN0RC0ERv)qRDOCDN#RM#8RCODC0FRDoRHOVRFs)Aqv41n_cc_1
.SzURR:H5VROHEFOIC_HE80Rc=R2CRoMNCs0RC
RSRRzR.g:FRVsRRHH5MR80CbEk_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0SC
-Q-RVNR58I8sHE80R4>R.M2RCRC80OFRs0CNCsRIHR0CCLMNDNCRMF8Rkk0b0MRCNCLDRD#CCRO0DHFoOR
RRRRRRzRSd:jRRRHV58N8s8IH0>ERR24.RMoCC0sNC-
S-HRVGFRVsNROD4DRd(UU,CR#D0CORRFV0#sH0CN0R0MFRHLCMsoRC#oH0CCs8R
RRRRRRRRRRRRRRFRskC0_M25HRR<='R4'IMECRq5)7_7)05lbNs88I0H8ER-48MFI04FR.=2RRRH2CCD#R''j;S
SSFSIkC0_M25HRR<='R4'IMECRN5I8C_so85N8HsI8-0E4FR8IFM0R24.RH-R2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0CHM52=R<RRW IMECRN5I8C_so85N8HsI8-0E4FR8IFM0R24.RH=R2DRC#'CRj
';RRRRRRRRS8CMRMoCC0sNCdRzjS;
-Q-RVNR58I8sHE80RR<=4R.2MIFRsCH0RNCMLRDCFFsRkk0b0MRCNCLDRD#CCRO0DHFoOCRMC88C
RRSRSRRzRd4:VRHR85N8HsI8R0E<4=R.o2RCsMCN
0CSSSSs0Fk_5CMH<2R=4R''S;
SISSF_k0CHM52=R<R''4;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R R;
RRRRRSRRCRM8oCCMsCN0R4zd;-
S-CRtMNCs00CRE)CRqOvRC#DDR8NMRH0s-N#00
C#RRRRRRRRS.zdRV:RF[sRRRHM58IH0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CRRRRRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FAVR)_qvcnjgXRc7:NRDLRCDH"#RW
";RRRRRRRRRRRRRRRRLHCoMR
RRRRRRRRRRARS)_qvcnjgXRc7:qR)vnA4__1c1Sc
RRRRRRRRRRRRb0FsRblNRQ57q>R=R_HMs5Coc+*[dFR8IFM0R[c*2q,R7q7)RR=>D_FII8N8s454RI8FMR0FjR2,7RQA=">Rjjjj"q,R7A7)RR=>D_FIs8N8s454RI8FMR0Fj
2,SSSS Rhq='>R4R',1q1)RR=>',j'RqW RR=>I_s0CHM52B,RpRiq=B>RpRi, RhA='>R4R',1A1)RR=>',j'RAW RR=>',j'RiBpA>R=RiBp,S
SSmS7q25dRR=>I0Fk_#Lkc,5HR[c*+,d2RS
SSmS7q25.RR=>I0Fk_#Lkc,5Hc+*[.R2,
SSSSq7m5R42=I>RF_k0Lck#5cH,*4[+2
,RSSSS75mqj=2R>FRIkL0_k5#cHc,R*,[2
SSSSA7m5Rd2=s>RF_k0Lck#5RH,c+*[dR2,
SSSSA7m5R.2=s>RF_k0Lck#5cH,*.[+2
,RSSSS75mA4=2R>FRskL0_k5#cH*,c[2+4,SR
S7SSmjA52>R=RksF0k_L#Hc5,*Rc[;22
SSSSksF0C_so*5c[<2R=FRskL0_k5#cH*,c[I2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRksF0C_so*5c[2+4RR<=s0Fk_#Lkc,5Hc+*[4I2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRksF0C_so*5c[2+.RR<=s0Fk_#Lkc,5Hc+*[.I2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRksF0C_so*5c[2+dRR<=s0Fk_#Lkc,5Hc+*[dI2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRkIF0C_so*5c[<2R=FRIkL0_k5#cH*,c[I2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRkIF0C_so*5c[2+4RR<=I0Fk_#Lkc,5Hc+*[4I2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRkIF0C_so*5c[2+.RR<=I0Fk_#Lkc,5Hc+*[.I2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRkIF0C_so*5c[2+dRR<=I0Fk_#Lkc,5Hc+*[dI2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
R
RRRRRRCRSMo8RCsMCNR0Cz;d.
RRRRCRSMo8RCsMCNR0Cz;.g
RRRR8CMRMoCC0sNC.RzU
;
SRRRRR--tCCMsCN0RC0ERv)qRDOCDN#RM#8RCODC0FRDoRHOVRFs)Aqv41n_gg_1
dSzdRR:H5VROHEFOIC_HE80Rg=R2CRoMNCs0RC
RSRRzRdc:FRVsRRHH5MR80CbEk_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0SC
-Q-RVNR58I8sHE80R4>R4M2RCRC80OFRs0CNCsRIHR0CCLMNDNCRMF8Rkk0b0MRCNCLDRD#CCRO0DHFoOR
RRRRRRzRSd:6RRRHV58N8s8IH0>ERR244RMoCC0sNC-
S-HRVGFRVsNROD4DRd(UU,CR#D0CORRFV0#sH0CN0R0MFRHLCMsoRC#oH0CCs8R
RRRRRRRRRRRRRRFRskC0_M25HRR<='R4'IMECRq5)7_7)05lbNs88I0H8ER-48MFI04FR4=2RRRH2CCD#R''j;S
SSFSIkC0_M25HRR<='R4'IMECRN5I8C_so85N8HsI8-0E4FR8IFM0R244RH=R2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0CHM52=R<RRW IMECRN5I8C_so85N8HsI8-0E4FR8IFM0R244RH=R2DRC#'CRj
';RRRRRRRRS8CMRMoCC0sNCdRz6S;
-Q-RVNR58I8sHE80RR<=4R42MIFRsCH0RNCMLRDCFFsRkk0b0MRCNCLDRD#CCRO0DHFoOCRMC88C
RRSRSRRzRdn:VRHR85N8HsI8R0E<4=R4o2RCsMCN
0CSRRRRRRRRRRRRksF0M_C5RH2<'=R4
';SSSSI0Fk_5CMH<2R=4R''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=W
 ;RRRRRRRRS8CMRMoCC0sNCdRznS;
-t-RCsMCNR0C0REC)RqvODCD#MRN8sR0H0-#N#0C
RRRRRRRRdSz(RR:VRFs[MRHRH5I8_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
RRRRRRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVAv)q_c.jU7XURD:RNDLCRRH#";W"
RRRRRRRRRRRRRRRRoLCHRM
RRRRRRRRRSRRAv)q_c.jU7XUR):Rq4vAng_1_
1gRRRRRRRRRRRRRRRRRFRbsl0RN5bR7RQq=H>RMC_so*5g[R+(8MFI0gFR*,[2R7q7)=qR>FRDIN_I858s48jRF0IMF2Rj,QR7A>R=Rj"jjjjjj,j"R7q7)=AR>FRDIN_s858s48jRF0IMF2Rj,R
RRRRRRRRRRRRRRRRRRRRRRRRRRhR q>R=R''4,1R1)=qR>jR''W,R =qR>sRI0M_C5,H2RiBpq>R=RiBp,hR A>R=R''4,1R1)=AR>jR''W,R =AR>jR''B,RpRiA=B>RpRi,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRq7m5R(2=I>RF_k0LUk#5UH,*([+2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mqn=2R>FRIkL0_k5#UH*,U[2+n,RR
RRRRRRRRRRRRRRRRRRRRRRRRR7RRm6q52>R=RkIF0k_L#HU5,[U*+,62RR
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7q25cRR=>I0Fk_#LkU,5HU+*[cR2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRq7m5Rd2=I>RF_k0LUk#5UH,*d[+2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mq.=2R>FRIkL0_k5#UH*,U[2+.,RR
RRRRRRRRRRRRRRRRRRRRRRRRR7RRm4q52>R=RkIF0k_L#HU5,[U*+,42RR
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7q25jRR=>I0Fk_#LkU,5HU2*[,RR
RRRRRRRRRRRRRRRRRRRRRRRRR7RRm(A52>R=RksF0k_L#HU5,[U*+,(2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7A25nRR=>s0Fk_#LkU,5HU+*[nR2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRA7m5R62=s>RF_k0LUk#5UH,*6[+2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mAc=2R>FRskL0_k5#UH*,U[2+c,RR
RRRRRRRRRRRRRRRRRRRRRRRRR7RRmdA52>R=RksF0k_L#HU5,[U*+,d2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7A25.RR=>s0Fk_#LkU,5HU+*[.R2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRA7m5R42=s>RF_k0LUk#5UH,*4[+2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mAj=2R>FRskL0_k5#UH*,U[R2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRu7Qq25jRR=>HsM_Cgo5*U[+27,RQRuA=">Rj
",RRRRRRRRRRRRRRRRRRRRRRRRRRRR7qmu5Rj2=I>RbHNs0L$_k5#UH2,[,mR7ujA52>R=RNsbs$H0_#LkU,5H[;22
RRRRRRRRRRRRRRRRksF0C_so*5g[<2R=FRskL0_k5#UH*,U[I2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRksF0C_so*5g[2+4RR<=s0Fk_#LkU,5HU+*[4I2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRksF0C_so*5g[2+.RR<=s0Fk_#LkU,5HU+*[.I2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRksF0C_so*5g[2+dRR<=s0Fk_#LkU,5HU+*[dI2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRksF0C_so*5g[2+cRR<=s0Fk_#LkU,5HU+*[cI2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRksF0C_so*5g[2+6RR<=s0Fk_#LkU,5HU+*[6I2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRksF0C_so*5g[2+nRR<=s0Fk_#LkU,5HU+*[nI2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRksF0C_so*5g[2+(RR<=s0Fk_#LkU,5HU+*[(I2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRksF0C_so*5g[2+URR<=ssbNH_0$LUk#5[H,2ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRI0Fk_osC5[g*2=R<RkIF0k_L#HU5,[U*2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRI0Fk_osC5[g*+R42<I=RF_k0LUk#5UH,*4[+2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRI0Fk_osC5[g*+R.2<I=RF_k0LUk#5UH,*.[+2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRI0Fk_osC5[g*+Rd2<I=RF_k0LUk#5UH,*d[+2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRI0Fk_osC5[g*+Rc2<I=RF_k0LUk#5UH,*c[+2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRI0Fk_osC5[g*+R62<I=RF_k0LUk#5UH,*6[+2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRI0Fk_osC5[g*+Rn2<I=RF_k0LUk#5UH,*n[+2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRI0Fk_osC5[g*+R(2<I=RF_k0LUk#5UH,*([+2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRI0Fk_osC5[g*+RU2<I=RbHNs0L$_k5#UH2,[RCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRSRRCRM8oCCMsCN0R(zd;R
RRSRRCRM8oCCMsCN0Rczd;R
RRMRC8CRoMNCs0zCRd
d;
RSRR-R-RMtCC0sNCER0CqR)vCRODRD#NRM8#CCDOD0RFOoHRsVFRv)qA_4n1_4U1
4USUzdRH:RVOR5EOFHCH_I8R0E=UR42CRoMNCs0RC
RSRRzRdg:FRVsRRHH5MR80CbEk_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0SC
-Q-RVNR58I8sHE80R4>RjM2RCRC80OFRs0CNCsRIHR0CCLMNDNCRMF8Rkk0b0MRCNCLDRD#CCRO0DHFoOR
RRRRRRzRSc:jRRRHV58N8s8IH0>ERR24jRMoCC0sNC-
S-HRVGFRVsNROD4DRd(UU,CR#D0CORRFV0#sH0CN0R0MFRHLCMsoRC#oH0CCs8R
RRRRRRRRRRRRRRFRskC0_M25HRR<='R4'IMECRq5)7_7)05lbNs88I0H8ER-48MFI04FRj=2RRRH2CCD#R''j;S
SSFSIkC0_M25HRR<='R4'IMECRN5I8C_so85N8HsI8-0E4FR8IFM0R24jRH=RRC2RDR#C';j'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RWRCIEMIR5Ns8_CNo58I8sHE80-84RF0IMFjR42RR=HC2RDR#C';j'
RRRRRRRRMSC8CRoMNCs0zCRc
j;SR--Q5VRNs88I0H8E=R<R24jRRMFI0sHCMRCNCLDRRFsFbk0kC0RMDNLCCR#D0CORoDFHMORCCC88S
RRRRRS4zcRH:RVNR58I8sHE80RR<=4Rj2oCCMsCN0
RSRRRRRRRRRRFRskC0_M25HRR<=';4'
SSSSkIF0M_C5RH2<'=R4
';RRRRRRRRRRRRRRRRI_s0CHM52=R<R;W 
RRRRRRRRMSC8CRoMNCs0zCRc
4;SR--tCCMsCN0RC0ERv)qRDOCDN#RM08Rs#H-0CN0#R
RRRRRRzRSc:.RRsVFRH[RMIR5HE80_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNCR
RRRRRRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqA)vj_4.4cXn:7RRLDNCHDR#WR""R;
RRRRRRRRRRRRRLRRCMoH
RRRRRRRRRRRR)SAq4v_jX.c4Rn7:qR)vnA4_U14_U14
RRRRRRRRRRRRRRRRbRRFRs0lRNb5q7QRR=>HsM_C4o5U+*[486RF0IMFUR4*,[2R7q7)=qR>FRDIN_I858sgFR8IFM0R,j2RA7QRR=>"jjjjjjjjjjjjjjjjR",q)77A>R=RIDF_8sN8gs5RI8FMR0Fj
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRR Rhq='>R4R',1q1)RR=>',j'RqW RR=>I_s0CHM52B,RpRiq=B>RpRi, RhA='>R4R',1A1)RR=>',j'RAW RR=>',j'RiBpA>R=RiBp,RR
RRRRRRRRRRRRRRRRRRRRRRRRR7RRm4q56=2R>FRIkL0_kn#454H,n+*[4,62RR
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7qc542>R=RkIF0k_L#54nHn,4*4[+cR2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRq7m524dRR=>I0Fk_#Lk4Hn5,*4n[d+42
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mq4R.2=I>RF_k0L4k#n,5H4[n*+24.,RR
RRRRRRRRRRRRRRRRRRRRRRRRR7RRm4q54=2R>FRIkL0_kn#454H,n+*[4,42RR
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7qj542>R=RkIF0k_L#54nHn,4*4[+jR2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRq7m5Rg2=I>RF_k0L4k#n,5H4[n*+,g2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7q25URR=>I0Fk_#Lk4Hn5,*4n[2+U,RR
RRRRRRRRRRRRRRRRRRRRRRRRR7RRm(q52>R=RkIF0k_L#54nHn,4*([+2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mqn=2R>FRIkL0_kn#454H,n+*[nR2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRq7m5R62=I>RF_k0L4k#n,5H4[n*+,62RR
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7q25cRR=>I0Fk_#Lk4Hn5,*4n[2+c,RR
RRRRRRRRRRRRRRRRRRRRRRRRR7RRmdq52>R=RkIF0k_L#54nHn,4*d[+2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mq.=2R>FRIkL0_kn#454H,n+*[.R2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRq7m5R42=I>RF_k0L4k#n,5H4[n*+,42RR
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7q25jRR=>I0Fk_#Lk4Hn5,*4n[R2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRA7m5246RR=>s0Fk_#Lk4Hn5,*4n[6+42
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mA4Rc2=s>RF_k0L4k#n,5H4[n*+24c,RR
RRRRRRRRRRRRRRRRRRRRRRRRR7RRm4A5d=2R>FRskL0_kn#454H,n+*[4,d2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7A.542>R=RksF0k_L#54nHn,4*4[+.R2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRA7m5244RR=>s0Fk_#Lk4Hn5,*4n[4+42
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mA4Rj2=s>RF_k0L4k#n,5H4[n*+24j,RR
RRRRRRRRRRRRRRRRRRRRRRRRR7RRmgA52>R=RksF0k_L#54nHn,4*g[+2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mAU=2R>FRskL0_kn#454H,n+*[UR2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRA7m5R(2=s>RF_k0L4k#n,5H4[n*+,(2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7A25nRR=>s0Fk_#Lk4Hn5,*4n[2+n,RR
RRRRRRRRRRRRRRRRRRRRRRRRR7RRm6A52>R=RksF0k_L#54nHn,4*6[+2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mAc=2R>FRskL0_kn#454H,n+*[cR2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRA7m5Rd2=s>RF_k0L4k#n,5H4[n*+,d2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7A25.RR=>s0Fk_#Lk4Hn5,*4n[2+.,RR
RRRRRRRRRRRRRRRRRRRRRRRRR7RRm4A52>R=RksF0k_L#54nHn,4*4[+2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mAj=2R>FRskL0_kn#454H,n2*[,RR
RRRRRRRRRRRRRRRRRRRRRRRRR7RRQRuq=H>RMC_soU54*4[+(FR8IFM0R*4U[n+427,RQRuA=">Rj,j"
RRRRRRRRRRRRRRRRRRRRRRRRRRRRu7mq254RR=>IsbNH_0$L4k#n,5H.+*[4R2,7qmu5Rj2=I>RbHNs0L$_kn#45.H,*,[2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRu7mA254RR=>ssbNH_0$L4k#n,5H.+*[4R2,7Amu5Rj2=s>RbHNs0L$_kn#45.H,*2[2;R
RRRRRRRRRRRRRRFRsks0_C4o5U2*[RR<=s0Fk_#Lk4Hn5,*4n[I2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRksF0C_soU54*4[+2=R<RksF0k_L#54nHn,4*4[+2ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRs0Fk_osC5*4U[2+.RR<=s0Fk_#Lk4Hn5,*4n[2+.RCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRsRRF_k0s5Co4[U*+Rd2<s=RF_k0L4k#n,5H4[n*+Rd2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRsks0_C4o5U+*[c<2R=FRskL0_kn#454H,n+*[cI2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRksF0C_soU54*6[+2=R<RksF0k_L#54nHn,4*6[+2ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRs0Fk_osC5*4U[2+nRR<=s0Fk_#Lk4Hn5,*4n[2+nRCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRsRRF_k0s5Co4[U*+R(2<s=RF_k0L4k#n,5H4[n*+R(2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRsks0_C4o5U+*[U<2R=FRskL0_kn#454H,n+*[UI2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRksF0C_soU54*g[+2=R<RksF0k_L#54nHn,4*g[+2ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRs0Fk_osC5*4U[j+42=R<RksF0k_L#54nHn,4*4[+jI2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRksF0C_soU54*4[+4<2R=FRskL0_kn#454H,n+*[4R42IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRsks0_C4o5U+*[4R.2<s=RF_k0L4k#n,5H4[n*+24.RCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRsRRF_k0s5Co4[U*+24dRR<=s0Fk_#Lk4Hn5,*4n[d+42ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRs0Fk_osC5*4U[c+42=R<RksF0k_L#54nHn,4*4[+cI2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRksF0C_soU54*4[+6<2R=FRskL0_kn#454H,n+*[4R62IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRsks0_C4o5U+*[4Rn2<s=RbHNs0L$_kn#45.H,*R[2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRsks0_C4o5U+*[4R(2<s=RbHNs0L$_kn#45.H,*4[+2ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';
RRRRRRRRRRRRRRRRkIF0C_soU54*R[2<I=RF_k0L4k#n,5H4[n*2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRI0Fk_osC5*4U[2+4RR<=I0Fk_#Lk4Hn5,*4n[2+4RCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRIRRF_k0s5Co4[U*+R.2<I=RF_k0L4k#n,5H4[n*+R.2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRIks0_C4o5U+*[d<2R=FRIkL0_kn#454H,n+*[dI2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRkIF0C_soU54*c[+2=R<RkIF0k_L#54nHn,4*c[+2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRI0Fk_osC5*4U[2+6RR<=I0Fk_#Lk4Hn5,*4n[2+6RCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRIRRF_k0s5Co4[U*+Rn2<I=RF_k0L4k#n,5H4[n*+Rn2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRIks0_C4o5U+*[(<2R=FRIkL0_kn#454H,n+*[(I2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRkIF0C_soU54*U[+2=R<RkIF0k_L#54nHn,4*U[+2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRI0Fk_osC5*4U[2+gRR<=I0Fk_#Lk4Hn5,*4n[2+gRCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRIRRF_k0s5Co4[U*+24jRR<=I0Fk_#Lk4Hn5,*4n[j+42ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRI0Fk_osC5*4U[4+42=R<RkIF0k_L#54nHn,4*4[+4I2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRkIF0C_soU54*4[+.<2R=FRIkL0_kn#454H,n+*[4R.2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRIks0_C4o5U+*[4Rd2<I=RF_k0L4k#n,5H4[n*+24dRCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRIRRF_k0s5Co4[U*+24cRR<=I0Fk_#Lk4Hn5,*4n[c+42ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRI0Fk_osC5*4U[6+42=R<RkIF0k_L#54nHn,4*4[+6I2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRkIF0C_soU54*4[+n<2R=bRIN0sH$k_L#54nH*,.[I2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRkIF0C_soU54*4[+(<2R=bRIN0sH$k_L#54nH*,.[2+4RCIEMIR5F_k0CHM52RR='24'R#CDCZR''
;
RRRRRRRRS8CMRMoCC0sNCcRz.R;
RRRRS8CMRMoCC0sNCdRzgR;
RCRRMo8RCsMCNR0Cz;dU
R
SR-RR-CRtMNCs00CRE)CRqOvRC#DDR8NMRD#CCRO0DHFoOFRVsqR)vnA4_n1d_n1d
dSzU:NRRRHV5FOEH_OCI0H8ERR=dRn2oCCMsCN0
RSRRdRzg:NRRsVFRHHRM8R5CEb0_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNC-
S-VRQR85N8HsI8R0E>2RgRCMC8FR0RCOsNR0CI0sHCMRCNCLDR8NMR0FkbRk0CLMND#CRCODC0FRDo
HOSzSScRjN:VRHR85N8HsI8R0E>2RgRMoCC0sNC-
S-HRVGFRVsNROD4DRd(UU,CR#D0CORRFV0#sH0CN0R0MFRHLCMsoRC#oH0CCs8S
SSFSskC0_M25HRR<='R4'IMECRq5)7_7)05lbNs88I0H8ER-48MFI0gFR2RR=HC2RDR#C';j'
SSSSkIF0M_C5RH2<'=R4I'RERCM58IN_osC58N8s8IH04E-RI8FMR0Fg=2RR2HRR#CDCjR''S;
SISSsC0_M25HRR<=WI RERCM58IN_osC58N8s8IH04E-RI8FMR0Fg=2RRRH2CCD#R''j;S
SS8CMRMoCC0sNCcRzj
N;SR--Q5VRNs88I0H8E=R<RRg2MIFRsCH0RNCMLRDCFFsRkk0b0MRCNCLDRD#CCRO0DHFoOCRMC88C
SSSzNc4RH:RVNR58I8sHE80RR<=go2RCsMCN
0CSSSSs0Fk_5CMH<2R=4R''S;
SISSF_k0CHM52=R<R''4;S
SSsSI0M_C5RH2<W=R S;
SMSC8CRoMNCs0zCRc;4N
-S-RMtCC0sNCER0CqR)vCRODRD#NRM80-sH#00NCS#
ScSz.:NRRsVFRH[RMIR5HE80_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNCR
RRRRRRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqA)v4_6..Xd7RR:DCNLD#RHR""W;R
RRRRRRRRRRRRRRCRLo
HMRRRRRRRRRRRRRRRRR)RAq6v_4d.X.:7RRv)qA_4n1_dn1
dnRRRRRRRRRRRRRRRRRRRRb0FsRblNRQ57q>R=R_HMs5Cod[n*+Rd48MFI0dFRn2*[,7Rq7R)q=D>RFII_Ns8858URF0IMF2Rj,QR7A>R=Rj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjj,j"R7q7)=AR>FRDIN_s858sUFR8IFM0R,j2
RRRRRRRRRRRRRRRRRRRRRRRRRRRR RRh=qR>4R''1,R1R)q='>RjR',WR q=I>RsC0_M25H,pRBi=qR>pRBi ,Rh=AR>4R''1,R1R)A='>RjR',WR A='>RjR',BApiRR=>B,pi
RRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRmdq54=2R>FRIkL0_k.#d5dH,.+*[d,42RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mqdRj2=I>RF_k0Ldk#.,5Hd[.*+2dj,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mq.Rg2=I>RF_k0Ldk#.,5Hd[.*+2.g,RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRq7m52.URR=>I0Fk_#LkdH.5,*d.[U+.2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7q(5.2>R=RkIF0k_L#5d.H.,d*.[+(
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7qn5.2>R=RkIF0k_L#5d.H.,d*.[+nR2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRm.q56=2R>FRIkL0_k.#d5dH,.+*[.,62RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mq.Rc2=I>RF_k0Ldk#.,5Hd[.*+2.c,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mq.Rd2=I>RF_k0Ldk#.,5Hd[.*+2.d,RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRq7m52..RR=>I0Fk_#LkdH.5,*d.[.+.2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7q45.2>R=RkIF0k_L#5d.H.,d*.[+4
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7qj5.2>R=RkIF0k_L#5d.H.,d*.[+jR2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRm4q5g=2R>FRIkL0_k.#d5dH,.+*[4,g2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mq4RU2=I>RF_k0Ldk#.,5Hd[.*+24U,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mq4R(2=I>RF_k0Ldk#.,5Hd[.*+24(,RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRq7m524nRR=>I0Fk_#LkdH.5,*d.[n+42
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7q6542>R=RkIF0k_L#5d.H.,d*4[+6
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7qc542>R=RkIF0k_L#5d.H.,d*4[+cR2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRm4q5d=2R>FRIkL0_k.#d5dH,.+*[4,d2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mq4R.2=I>RF_k0Ldk#.,5Hd[.*+24.,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mq4R42=I>RF_k0Ldk#.,5Hd[.*+244,RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRq7m524jRR=>I0Fk_#LkdH.5,*d.[j+42
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7q25gRR=>I0Fk_#LkdH.5,*d.[2+g,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mqU=2R>FRIkL0_k.#d5dH,.+*[UR2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRm(q52>R=RkIF0k_L#5d.H.,d*([+2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7q25nRR=>I0Fk_#LkdH.5,*d.[2+n,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mq6=2R>FRIkL0_k.#d5dH,.+*[6R2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRmcq52>R=RkIF0k_L#5d.H.,d*c[+2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7q25dRR=>I0Fk_#LkdH.5,*d.[2+d,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mq.=2R>FRIkL0_k.#d5dH,.+*[.R2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRm4q52>R=RkIF0k_L#5d.H.,d*4[+2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7q25jRR=>I0Fk_#LkdH.5,*d.[
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7A45d2>R=RksF0k_L#5d.H.,d*d[+4R2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRmdA5j=2R>FRskL0_k.#d5dH,.+*[d,j2
RRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRm.A5g=2R>FRskL0_k.#d5dH,.+*[.,g2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mA.RU2=s>RF_k0Ldk#.,5Hd[.*+2.U,RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRA7m52.(RR=>s0Fk_#LkdH.5,*d.[(+.2R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRA7m52.nRR=>s0Fk_#LkdH.5,*d.[n+.2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7A65.2>R=RksF0k_L#5d.H.,d*.[+6R2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRm.A5c=2R>FRskL0_k.#d5dH,.+*[.,c2
RRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRm.A5d=2R>FRskL0_k.#d5dH,.+*[.,d2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mA.R.2=s>RF_k0Ldk#.,5Hd[.*+2..,RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRA7m52.4RR=>s0Fk_#LkdH.5,*d.[4+.2R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRA7m52.jRR=>s0Fk_#LkdH.5,*d.[j+.2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7Ag542>R=RksF0k_L#5d.H.,d*4[+gR2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRm4A5U=2R>FRskL0_k.#d5dH,.+*[4,U2
RRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRm4A5(=2R>FRskL0_k.#d5dH,.+*[4,(2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mA4Rn2=s>RF_k0Ldk#.,5Hd[.*+24n,RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRA7m5246RR=>s0Fk_#LkdH.5,*d.[6+42R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRA7m524cRR=>s0Fk_#LkdH.5,*d.[c+42
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7Ad542>R=RksF0k_L#5d.H.,d*4[+dR2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRm4A5.=2R>FRskL0_k.#d5dH,.+*[4,.2
RRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRm4A54=2R>FRskL0_k.#d5dH,.+*[4,42RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mA4Rj2=s>RF_k0Ldk#.,5Hd[.*+24j,RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRA7m5Rg2=s>RF_k0Ldk#.,5Hd[.*+,g2
RRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRmUA52>R=RksF0k_L#5d.H.,d*U[+2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7A25(RR=>s0Fk_#LkdH.5,*d.[2+(,RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRA7m5Rn2=s>RF_k0Ldk#.,5Hd[.*+,n2
RRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRm6A52>R=RksF0k_L#5d.H.,d*6[+2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7A25cRR=>s0Fk_#LkdH.5,*d.[2+c,RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRA7m5Rd2=s>RF_k0Ldk#.,5Hd[.*+,d2
RRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRm.A52>R=RksF0k_L#5d.H.,d*.[+2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7A254RR=>s0Fk_#LkdH.5,*d.[2+4,RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRA7m5Rj2=s>RF_k0Ldk#.,5Hd[.*2R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRu7Qq>R=R_HMs5Cod[n*+Rd68MFI0dFRn+*[d,.2Ru7QA>R=Rj"jj,j"
RRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRm5uqd=2R>bRIN0sH$k_L#5d.H*,c[2+d,mR7u.q52>R=RNIbs$H0_#LkdH.5,[c*+,.2
RRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRm5uq4=2R>bRIN0sH$k_L#5d.H*,c[2+4,mR7ujq52>R=RNIbs$H0_#LkdH.5,[c*2R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRu7mA25dRR=>ssbNH_0$Ldk#.,5Hc+*[dR2,7Amu5R.2=s>RbHNs0L$_k.#d5cH,*.[+2R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRu7mA254RR=>ssbNH_0$Ldk#.,5Hc+*[4R2,7Amu5Rj2=s>RbHNs0L$_k.#d5cH,*2[2;R
RRRRRRRRRRRRRRRRRs0Fk_osC5*dn[<2R=FRskL0_k.#d5dH,.2*[RCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRksF0C_son5d*4[+2=R<RksF0k_L#5d.H.,d*4[+2ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRsks0_Cdo5n+*[.<2R=FRskL0_k.#d5dH,.+*[.I2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRsRRF_k0s5Cod[n*+Rd2<s=RF_k0Ldk#.,5Hd[.*+Rd2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRs0Fk_osC5*dn[2+cRR<=s0Fk_#LkdH.5,*d.[2+cRCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRksF0C_son5d*6[+2=R<RksF0k_L#5d.H.,d*6[+2ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRsks0_Cdo5n+*[n<2R=FRskL0_k.#d5dH,.+*[nI2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRsRRF_k0s5Cod[n*+R(2<s=RF_k0Ldk#.,5Hd[.*+R(2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRs0Fk_osC5*dn[2+URR<=s0Fk_#LkdH.5,*d.[2+URCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRksF0C_son5d*g[+2=R<RksF0k_L#5d.H.,d*g[+2ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRsks0_Cdo5n+*[4Rj2<s=RF_k0Ldk#.,5Hd[.*+24jRCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRksF0C_son5d*4[+4<2R=FRskL0_k.#d5dH,.+*[4R42IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRs0Fk_osC5*dn[.+42=R<RksF0k_L#5d.H.,d*4[+.I2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRsRRF_k0s5Cod[n*+24dRR<=s0Fk_#LkdH.5,*d.[d+42ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRsks0_Cdo5n+*[4Rc2<s=RF_k0Ldk#.,5Hd[.*+24cRCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRksF0C_son5d*4[+6<2R=FRskL0_k.#d5dH,.+*[4R62IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRs0Fk_osC5*dn[n+42=R<RksF0k_L#5d.H.,d*4[+nI2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRsRRF_k0s5Cod[n*+24(RR<=s0Fk_#LkdH.5,*d.[(+42ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRsks0_Cdo5n+*[4RU2<s=RF_k0Ldk#.,5Hd[.*+24URCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRksF0C_son5d*4[+g<2R=FRskL0_k.#d5dH,.+*[4Rg2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRs0Fk_osC5*dn[j+.2=R<RksF0k_L#5d.H.,d*.[+jI2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRsRRF_k0s5Cod[n*+2.4RR<=s0Fk_#LkdH.5,*d.[4+.2ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRsks0_Cdo5n+*[.R.2<s=RF_k0Ldk#.,5Hd[.*+2..RCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRksF0C_son5d*.[+d<2R=FRskL0_k.#d5dH,.+*[.Rd2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRs0Fk_osC5*dn[c+.2=R<RksF0k_L#5d.H.,d*.[+cI2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRsRRF_k0s5Cod[n*+2.6RR<=s0Fk_#LkdH.5,*d.[6+.2ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRsks0_Cdo5n+*[.Rn2<s=RF_k0Ldk#.,5Hd[.*+2.nRCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRksF0C_son5d*.[+(<2R=FRskL0_k.#d5dH,.+*[.R(2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRs0Fk_osC5*dn[U+.2=R<RksF0k_L#5d.H.,d*.[+UI2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRsRRF_k0s5Cod[n*+2.gRR<=s0Fk_#LkdH.5,*d.[g+.2ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRsks0_Cdo5n+*[dRj2<s=RF_k0Ldk#.,5Hd[.*+2djRCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRksF0C_son5d*d[+4<2R=FRskL0_k.#d5dH,.+*[dR42IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRs0Fk_osC5*dn[.+d2=R<RNsbs$H0_#LkdH.5,[c*2ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRsks0_Cdo5n+*[dRd2<s=RbHNs0L$_k.#d5cH,*4[+2ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRsks0_Cdo5n+*[dRc2<s=RbHNs0L$_k.#d5cH,*.[+2ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRsks0_Cdo5n+*[dR62<s=RbHNs0L$_k.#d5cH,*d[+2ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRR
RRRRRRRRRRRRRRRRRkIF0C_son5d*R[2<I=RF_k0Ldk#.,5Hd[.*2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRIks0_Cdo5n+*[4<2R=FRIkL0_k.#d5dH,.+*[4I2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRIRRF_k0s5Cod[n*+R.2<I=RF_k0Ldk#.,5Hd[.*+R.2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRI0Fk_osC5*dn[2+dRR<=I0Fk_#LkdH.5,*d.[2+dRCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRkIF0C_son5d*c[+2=R<RkIF0k_L#5d.H.,d*c[+2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRIks0_Cdo5n+*[6<2R=FRIkL0_k.#d5dH,.+*[6I2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRIRRF_k0s5Cod[n*+Rn2<I=RF_k0Ldk#.,5Hd[.*+Rn2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRI0Fk_osC5*dn[2+(RR<=I0Fk_#LkdH.5,*d.[2+(RCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRkIF0C_son5d*U[+2=R<RkIF0k_L#5d.H.,d*U[+2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRIks0_Cdo5n+*[g<2R=FRIkL0_k.#d5dH,.+*[gI2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRIRRF_k0s5Cod[n*+24jRR<=I0Fk_#LkdH.5,*d.[j+42ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRIks0_Cdo5n+*[4R42<I=RF_k0Ldk#.,5Hd[.*+244RCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRkIF0C_son5d*4[+.<2R=FRIkL0_k.#d5dH,.+*[4R.2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRI0Fk_osC5*dn[d+42=R<RkIF0k_L#5d.H.,d*4[+dI2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRIRRF_k0s5Cod[n*+24cRR<=I0Fk_#LkdH.5,*d.[c+42ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRIks0_Cdo5n+*[4R62<I=RF_k0Ldk#.,5Hd[.*+246RCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRkIF0C_son5d*4[+n<2R=FRIkL0_k.#d5dH,.+*[4Rn2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRI0Fk_osC5*dn[(+42=R<RkIF0k_L#5d.H.,d*4[+(I2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRIRRF_k0s5Cod[n*+24URR<=I0Fk_#LkdH.5,*d.[U+42ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRIks0_Cdo5n+*[4Rg2<I=RF_k0Ldk#.,5Hd[.*+24gRCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRkIF0C_son5d*.[+j<2R=FRIkL0_k.#d5dH,.+*[.Rj2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRI0Fk_osC5*dn[4+.2=R<RkIF0k_L#5d.H.,d*.[+4I2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRIRRF_k0s5Cod[n*+2..RR<=I0Fk_#LkdH.5,*d.[.+.2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRIks0_Cdo5n+*[.Rd2<I=RF_k0Ldk#.,5Hd[.*+2.dRCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRkIF0C_son5d*.[+c<2R=FRIkL0_k.#d5dH,.+*[.Rc2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRI0Fk_osC5*dn[6+.2=R<RkIF0k_L#5d.H.,d*.[+6I2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRIRRF_k0s5Cod[n*+2.nRR<=I0Fk_#LkdH.5,*d.[n+.2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRIks0_Cdo5n+*[.R(2<I=RF_k0Ldk#.,5Hd[.*+2.(RCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRkIF0C_son5d*.[+U<2R=FRIkL0_k.#d5dH,.+*[.RU2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRI0Fk_osC5*dn[g+.2=R<RkIF0k_L#5d.H.,d*.[+gI2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRIRRF_k0s5Cod[n*+2djRR<=I0Fk_#LkdH.5,*d.[j+d2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRIks0_Cdo5n+*[dR42<I=RF_k0Ldk#.,5Hd[.*+2d4RCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRkIF0C_son5d*d[+.<2R=bRIN0sH$k_L#5d.H*,c[I2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRIRRF_k0s5Cod[n*+2ddRR<=IsbNH_0$Ldk#.,5Hc+*[4I2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRIRRF_k0s5Cod[n*+2dcRR<=IsbNH_0$Ldk#.,5Hc+*[.I2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRIRRF_k0s5Cod[n*+2d6RR<=IsbNH_0$Ldk#.,5Hc+*[dI2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
S
SS8CMRMoCC0sNCcRz.
N;SMSC8CRoMNCs0zCRd;gN
MSC8CRoMNCs0zCRd;UN
CRRMo8RCsMCNR0Cz;cd
R
RzRcc:VRHRF5M0NRs8_8ss2CoRMoCC0sNC-R-RMoCC0sNCCR#D0CORlsN
RRRRR--QNVR8I8sHE80R6<RR#N#HRoM'Rj'0kFRMCk#8HRL0R#
RzRRj:RRRRHV58N8s8IH0=ERRR42oCCMsCN0
RRRRRRRRIDF_8sN8#s_RR<="jjjjRj"&NRs8C_so5_#j
2;RRRRRRRRD_FII8N8sR_#<"=Rjjjjj&"RR8IN_osC_j#52R;
RCRRMo8RCsMCNR0Cz
j;RRRRzR4R:VRHR85N8HsI8R0E=2R.RMoCC0sNCR
RRRRRRFRDIN_s8_8s#=R<Rj"jjRj"&NRs8C_so5_#4FR8IFM0R;j2
RRRRRRRRIDF_8IN8#s_RR<="jjjj&"RR8IN_osC_4#5RI8FMR0Fj
2;RRRRCRM8oCCMsCN0R;z4
RRRRRz.RH:RVNR58I8sHE80Rd=R2CRoMNCs0RC
RRRRRDRRFsI_Ns88_<#R=jR"jRj"&NRs8C_so5_#.FR8IFM0R;j2
RRRRRRRRIDF_8IN8#s_RR<="jjj"RR&I_N8s_Co#R5.8MFI0jFR2R;
RCRRMo8RCsMCNR0Cz
.;RRRRzRdR:VRHR85N8HsI8R0E=2RcRMoCC0sNCR
RRRRRRFRDIN_s8_8s#=R<Rj"j"RR&s_N8s_Co#R5d8MFI0jFR2R;
RRRRRDRRFII_Ns88_<#R=jR"j&"RR8IN_osC_d#5RI8FMR0Fj
2;RRRRCRM8oCCMsCN0R;zd
cSzSH:RVNR58I8sHE80R6=R2CRoMNCs0SC
SIDF_8sN8#s_RR<='Rj'&NRs8C_so5_#cFR8IFM0R;j2
DSSFII_Ns88_<#R=jR''RR&I_N8s_Co#R5c8MFI0jFR2S;
CRM8oCCMsCN0R;zc
RRRRRz6RH:RVNR58I8sHE80R6>R2CRoMNCs0RC
RRRRRDRRFsI_Ns88_<#R=NRs8C_so5_#6FR8IFM0R;j2
RRRRRRRRIDF_8IN8#s_RR<=I_N8s_Co#R568MFI0jFR2R;
RCRRMo8RCsMCNR0Cz
6;
RRRRR--Q5VR8_HMs2CoRosCHC#0sQR7h#RkHRMoB
piRRRRzRnR:VRHRH58MC_soo2RCsMCN
0CRRRRRRRRbOsFCR##5iBp,QR7hL2RCMoH
RRRRRRRRRRRRRHV5iBpR'=R4N'RMB8RpCi'P0CM2ER0CRM
RRRRRRRRRRRRRHRRMC_soR_#<7=RQ
h;RRRRRRRRRRRRCRM8H
V;RRRRRRRRCRM8bOsFC;##
RRRR8CMRMoCC0sNCnRz;R
RR(RzRRR:H5VRMRF08_HMs2CoRMoCC0sNCR
RRRRRRRRRRMRH_osC_<#R=QR7hR;
RCRRMo8RCsMCNR0Cz
(;
RRRRR--Q5VRsk8F0C_sos2RC#oH0RCs7amzRHk#MmoRB
piRRRRzRUsRH:RVsR580Fk_osC2CRoMNCs0RC
RRRRRbRRsCFO#5#R)B_mpRi,s0Fk_osC_R#2LHCoMR
RRRRRRRRRRVRHR_5)miBpR'=R4N'RM)8R_pmBiP'CC2M0RC0EMR
RRRRRRRRRRRRRR_R)7amzRR<=s0Fk_osC_
#;RRRRRRRRRRRRCRM8H
V;RRRRRRRRCRM8bOsFC;##
RRRR8CMRMoCC0sNCURzsR;
RzRRgRsR:VRHRF5M08RsF_k0s2CoRMoCC0sNCR
RRRRRRRRRR_R)7amzRR<=s0Fk_osC_
#;RRRRCRM8oCCMsCN0Rszg;S

zRUIRH:RVIR580Fk_osC2CRoMNCs0RC
RRRRRbRRsCFO#5#RWB_mpRi,I0Fk_osC_R#2LHCoMR
RRRRRRRRRRVRHR_5WmiBpR'=R4N'RMW8R_pmBiP'CC2M0RC0EMR
RRRRRRRRRRRRRR_RW7amzRR<=I0Fk_osC_
#;RRRRRRRRRRRRCRM8H
V;RRRRRRRRCRM8bOsFC;##
RRRR8CMRMoCC0sNCURzIR;
RzRRgRIR:VRHRF5M08RIF_k0s2CoRMoCC0sNCR
RRRRRRRRRR_RW7amzRR<=I0Fk_osC_
#;RRRRCRM8oCCMsCN0RIzg;R

R-RR-VRQRN5s8_8ss2CoRosCHC#0s7Rq7k)R#oHMRiBp
RRRRjz4RRR:H5VRs8N8sC_soo2RCsMCN
0CRRRRRRRRbOsFCR##5m)_B,piR7)q7R)2LHCoMR
RRRRRRRRRRVRHR_5)miBpR'=R4N'RM)8R_pmBiP'CC2M0RC0EMR
RRRRRRRRRRRRRRNRs8C_soR_#<)=Rq)7758N8s8IH04E-RI8FMR0Fj
2;RRRRRRRRRRRRCRM8H
V;RRRRRRRRCRM8bOsFC;##
RRRR8CMRMoCC0sNC4RzjR;
RzRR4:4RRRHV50MFR8sN8ss_CRo2oCCMsCN0
RRRRRRRRRRRR8sN_osC_<#R=qR)7;7)
RRRR8CMRMoCC0sNC4Rz4
;
RRRR-Q-RVIR5Ns88_osC2CRso0H#CqsR7R7)kM#HopRBiR
RR4Rz.:RRRRHV58IN8ss_CRo2oCCMsCN0
RRRRRRRRFbsO#C#Rp5BiW,Rq)772CRLo
HMRRRRRRRRRRRRH5VRBRpi=4R''MRN8pRBiP'CC2M0RC0EMR
RRRRRRRRRRRRRRNRI8C_soR_#<W=Rq)7758N8s8IH04E-RI8FMR0Fj
2;RRRRRRRRRRRRCRM8H
V;RRRRRRRRCRM8bOsFC;##
RRRR8CMRMoCC0sNC4Rz.R;
RzRR4:dRRRHV50MFR8IN8ss_CRo2oCCMsCN0
RRRRRRRRRRRR8IN_osC_<#R=qRW7;7)
RRRR8CMRMoCC0sNC4RzdR;
RRRRR
RRRRRR-t-RCsMCNR0C0REC)RqvODCD#MRN8CR#D0CORoDFHRO
RzRR4:cRRsVFRHHRMMR5kOl_C_DDn-cRRR428MFI0jFRRMoCC0sNCR
RR-R-RRQV58N8s8IH0>ERRR62M8CCRR0FONsC0ICRsCH0RNCMLRDCNRM8Fbk0kC0RMDNLCCR#D0CORoDFHRO
RRRRRzRR4:6RRRHV58N8s8IH0>ERRRn2oCCMsCN0
RRRRRRRRRRRRRRRRksF0M_C_H#52=R<R''4RCIEMsR5Ns8_C#o_58N8s8IH04E-RI8FMR0Fn=2RRRH2CCD#R''j;S
SSFSIkC0_M5_#H<2R=4R''ERIC5MRI_N8s_Co#85N8HsI8-0E4FR8IFM0RRn2=2RHR#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_M5_#H<2R= RWRCIEMIR5Ns8_C#o_58N8s8IH04E-RI8FMR0Fn=2RRRH2CCD#R''j;R
RRRRRRMRC8CRoMNCs0zCR4
6;RRRR-Q-RVNR58I8sHE80RR<=6M2RFsRIHR0CCLMNDFCRskRF00bkRNCMLRDC#CCDOD0RFOoHRCMC8
C8RRRRRRRRzR4n:VRHR85N8HsI8R0E<n=R2CRoMNCs0RC
RRRRRRRRRRRRRsRRF_k0C#M_5RH2<'=R4
';SSSSI0Fk__CM#25HRR<=';4'
RRRRRRRRRRRRRRRR0Is__CM#25HRR<=W
 ;RRRRRRRRCRM8oCCMsCN0Rnz4;R
RR-R-RMtCC0sNCER0CqR)vCRODRD#NRM80-sH#00NCR#
RRRRRzRR4:(RRsVFRH[RMIR5HE80R4-R2FR8IFM0RojRCsMCN
0CRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FzVR)nqvcRR:DCNLD#RHR7"1a&"RR0HMCsoC'NHloIC5HE802RR&"R7"&MRH0CCosl'HN5oCHc*n2RR&"RW"&MRH0CCosl'HN5oC[&2RR"" RH&RMo0CCHs'lCNo50oC_8CM_b8C05E5H2+4*,ncRb8C02E2R"&RX&"RR0HMCsoC'NHlo[C5+;42
RRRRRRRRRRRRoLCHRM
RRRRRRRRRzRR)nqvcRR:Xv)qn4cX7RR
RRRRRRRRRRRRRbRRFRs0lRNb5=7R>MRH_osC_[#52q,Rj>R=RIDF_8IN8#s_5,j2RRq4=D>RFII_Ns88_4#52q,R.>R=RIDF_8IN8#s_5,.2
RRRRRRRRRRRRRRRRRRRRRRRRqRRd>R=RIDF_8IN8#s_5,d2RRqc=D>RFII_Ns88_c#52q,R6>R=RIDF_8IN8#s_5,62RS
SSSSSRuR7)Rqj=D>RFsI_Ns88_j#527,Ru4)qRR=>D_FIs8N8s5_#4R2,7qu).>R=RIDF_8sN8#s_5,.2
SSSSRSSR)7uq=dR>FRDIN_s8_8s#25d,uR7)Rqc=D>RFsI_Ns88_c#527,Ru6)qRR=>D_FIs8N8s5_#6R2,
SSSSRSSRRW =I>RsC0_M5_#HR2,WiBpRR=>B,piRm7uRR=>s0Fk_#Lk_#nc5[H,21,Ru=mR>FRIkL0_kn#_cH#5,2[2;R
RRRRRRRRRRRRRRFRsks0_C#o_5R[2<s=RF_k0L_k#n5c#H2,[RCIEMsR5F_k0C#M_5RH2=4R''C2RDR#C';Z'
SSSSkIF0C_so5_#[<2R=FRIkL0_kn#_cH#5,R[2IMECRF5IkC0_M5_#H=2RR''42DRC#'CRZ
';RRRRRRRRCRM8oCCMsCN0R(z4;R
RRCRRMo8RCsMCNR0Cz;4cRRRRRRRRRRRR
RRRR
RRRRRR-t-RCsMCNR0CN.RdRsIF8CR8C)bRqOvRCRDDHNVRbFbsbNsH0RCRRRRRRRRRRRRRRR
RR4RzURR:H5VRM_klODCD_Rd.=2R4RMoCC0sNCR
RR-R-RRQV58N8s8IH0>ERRR(2M8CCRR0FONsC0ICRsCH0RNCMLRDCNRM8Fbk0kC0RMDNLCCR#D0CORoDFHRO
RRRRRzRR4RgN:VRHR85N8HsI8R0E>2RnRMoCC0sNCR
RRRRRRRRRRRRRRFRskC0_M._dRR<='R4'IMECRs55Ns8_C#o_58N8s8IH04E-RI8FMR0Fn=2RRlMk_DOCDc_n2MRN8sR5Ns8_C#o_5R62=jR''R22CCD#R''j;S
SSFSIkC0_M._dRR<='R4'IMECRI55Ns8_C#o_58N8s8IH04E-RI8FMR0Fn=2RRlMk_DOCDc_n2MRN8IR5Ns8_C#o_5R62=jR''R22CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C_Rd.<W=R ERIC5MR58IN_osC_N#58I8sHE80-84RF0IMF2RnRM=RkOl_C_DDnRc2NRM858IN_osC_6#52RR='2j'2DRC#'CRj
';RRRRRRRRCRM8oCCMsCN0Rgz4NR;
RRRRRzRR4RgL:VRHR85N8HsI8R0E=RRnNRM8M_klODCD_Rnc=2RjRMoCC0sNCR
RRRRRRRRRRRRRRFRskC0_M._dRR<='R4'IMECRs55Ns8_C#o_5R62=jR''R22CCD#R''j;S
SSFSIkC0_M._dRR<='R4'IMECRI55Ns8_C#o_5R62=jR''R22CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C_Rd.<W=R ERIC5MR58IN_osC_6#52RR='2j'2DRC#'CRj
';RRRRRRRRCRM8oCCMsCN0Rgz4LR;RR-R-RRQV58N8s8IH0<ER=2R6RRMFI0sHCMRCNCLDRRFsFbk0kC0RMDNLCCR#D0CORoDFHMORCCC88R
RRRRRR.RzjRR:H5VRNs88I0H8E=R<RR62oCCMsCN0
RRRRRRRRRRRRRRRRksF0M_C_Rd.<'=R4
';SSSSI0Fk__CMd<.R=4R''R;
RRRRRRRRRRRRRIRRsC0_M._dRR<=W
 ;RRRRRRRRCRM8oCCMsCN0Rjz.;R
RR-R-RMtCC0sNCER0CqR)vCRODNDRM08Rs#H-0CN0
RRRRRRRR4z.RV:RF[sRRRHM58IH0-ERRR428MFI0jFRRMoCC0sNCR
RRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqz)vRd.:NRDLRCDH"#R1"7aRH&RMo0CCHs'lCNo58IH0RE2&7R""RR&HCM0o'CsHolNCk5MlC_ODnD_cc*n2RR&"RW"&MRH0CCosl'HN5oC[&2RR"" RH&RMo0CCHs'lCNo50oC_8CM_b8C0ME5kOl_C_DDnnc*cRR+dR.,80CbER22&XR""RR&HCM0o'CsHolNC+5[4
2;RRRRRRRRRRRRLHCoMR
RRRRRRRRRR)Rzq.vdRX:R)dqv.7X4RR
RRRRRRRRRRRRRRFRbsl0RN5bR7>R=R_HMs_Co#25[,jRqRR=>D_FII8N8s5_#jR2,q=4R>FRDIN_I8_8s#254,.RqRR=>D_FII8N8s5_#.
2,RRRRRRRRRRRRRRRRRRRRRRRRRdRqRR=>D_FII8N8s5_#dR2,q=cR>FRDIN_I8_8s#25c,SR
SSSSS7RRuj)qRR=>D_FIs8N8s5_#jR2,7qu)4>R=RIDF_8sN8#s_5,42R)7uq=.R>FRDIN_s8_8s#25.,S
SSSSSRuR7)Rqd=D>RFsI_Ns88_d#527,Ruc)qRR=>D_FIs8N8s5_#cR2,
SSSSRSSRRW =I>RsC0_M._d,BRWp=iR>pRBi7,Ru=mR>FRskL0_kd#_.M#5kOl_C_DDd[.,21,Ru=mR>FRIkL0_kd#_.M#5kOl_C_DDd[.,2
2;RRRRRRRRRRRRRRRRs0Fk_osC_[#52=R<RksF0k_L#._d#k5MlC_ODdD_.2,[RCIEMsR5F_k0CdM_.RR='24'R#CDCZR''S;
SISSF_k0s_Co#25[RR<=I0Fk_#Lk_#d.5lMk_DOCD._d,R[2IMECRF5IkC0_M._dR'=R4R'2CCD#R''Z;R
RRRRRRCRRMo8RCsMCNR0Cz;.4
RRRRMRC8CRoMNCs0zCR4RU;RRRRRRRRRR

R-RR-CRtMNCs0NCRRR4nI8FsRC8CbqR)vCRODHDRVbRNbbsFs0HNCRRRRRRRRRRRRRRR
RRRR.z.RH:RVMR5kOl_C_DD4=nRRR42oCCMsCN0
RRRRR--Q5VRNs88I0H8ERR>6M2RCRC80OFRs0CNCsRIHR0CCLMNDNCRMF8Rkk0b0MRCNCLDRD#CCRO0DHFoOR
RRRRRR.Rzd:NRRRHV58N8s8IH0>ERRNnRMM8RkOl_C_DDd=.RRR42oCCMsCN0
RRRRRRRRRRRRRRRRksF0M_C_R4n<'=R4I'RERCM5N5s8C_so5_#Ns88I0H8ER-48MFI0nFR2RR=M_klODCD_2ncR8NMRN5s8C_so5_#6=2RR''42MRN8sR5Ns8_C#o_5Rc2=jR''R22CCD#R''j;S
SSFSIkC0_Mn_4RR<='R4'IMECRI55Ns8_C#o_58N8s8IH04E-RI8FMR0Fn=2RRlMk_DOCDc_n2MRN8IR5Ns8_C#o_5R62=4R''N2RM58RI_N8s_Co#25cR'=Rj2'2R#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_Mn_4RR<=WI RERCM5N5I8C_so5_#Ns88I0H8ER-48MFI0nFR2RR=M_klODCD_2ncR8NMRN5I8C_so5_#6=2RR''42MRN8IR5Ns8_C#o_5Rc2=jR''R22CCD#R''j;R
RRRRRRMRC8CRoMNCs0zCR.;dN
RRRRRRRRdz.LRR:H5VRNs88I0H8ERR>nMRN8kRMlC_ODdD_.=R/RR42oCCMsCN0
RRRRRRRRRRRRRRRRksF0M_C_R4n<'=R4I'RERCM5N5s8C_so5_#Ns88I0H8ER-48MFI0nFR2RR=M_klODCD_2ncR8NMRN5s8C_so5_#6=2RR''j2MRN8sR5Ns8_C#o_5Rc2=jR''R22CCD#R''j;S
SSFSIkC0_Mn_4RR<='R4'IMECRI55Ns8_C#o_58N8s8IH04E-RI8FMR0Fn=2RRlMk_DOCDc_n2MRN8IR5Ns8_C#o_5R62=jR''N2RM58RI_N8s_Co#25cR'=Rj2'2R#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_Mn_4RR<=WI RERCM5N5I8C_so5_#Ns88I0H8ER-48MFI0nFR2RR=M_klODCD_2ncR8NMRN5I8C_so5_#6=2RR''j2MRN8IR5Ns8_C#o_5Rc2=jR''R22CCD#R''j;R
RRRRRRMRC8CRoMNCs0zCR.;dL
RRRRRRRRdz.ORR:H5VRNs88I0H8ERR=nMRN8kRMlC_ODdD_.RR=4o2RCsMCN
0CRRRRRRRRRRRRRRRRs0Fk__CM4<nR=4R''ERIC5MR58sN_osC_6#52RR='24'R8NMRN5s8C_so5_#c=2RR''j2C2RDR#C';j'
SSSSkIF0M_C_R4n<'=R4I'RERCM5N5I8C_so5_#6=2RR''42MRN8IR5Ns8_C#o_5Rc2=jR''R22CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C_R4n<W=R ERIC5MR58IN_osC_6#52RR='24'R8NMRN5I8C_so5_#c=2RR''j2C2RDR#C';j'
RRRRRRRR8CMRMoCC0sNC.Rzd
O;RRRRRRRRz8.dRH:RVNR58I8sHE80R6=RR8NMRlMk_DOCD._dRR/=4o2RCsMCN
0CRRRRRRRRRRRRRRRRs0Fk__CM4<nR=4R''ERIC5MR58sN_osC_N#58I8sHE80-84RF0IMF2RcRM=RkOl_C_DDd2.2R#CDCjR''S;
SISSF_k0C4M_n=R<R''4RCIEM5R5I_N8s_Co#85N8HsI8-0E4FR8IFM0RRc2=kRMlC_ODdD_.R22CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C_R4n<W=R ERIC5MR58IN_osC_N#58I8sHE80-84RF0IMF2RcRM=RkOl_C_DDd2.2R#CDCjR''R;
RRRRRCRRMo8RCsMCNR0Cz8.d;RRRRR--Q5VRNs88I0H8E=R<RR62MIFRsCH0RNCMLRDCFFsRkk0b0MRCNCLDRD#CCRO0DHFoOCRMC88C
RRRRRRRRcz.RH:RVNR58I8sHE80RR<=co2RCsMCN
0CRRRRRRRRRRRRRRRRs0Fk__CM4<nR=4R''S;
SISSF_k0C4M_n=R<R''4;R
RRRRRRRRRRRRRRsRI0M_C_R4n<W=R R;
RRRRRCRRMo8RCsMCNR0Cz;.c
RRRRR--tCCMsCN0RC0ERv)qRDOCDMRN8sR0H0-#N
0CRRRRRRRRzR.6:FRVsRR[H5MRI0H8ERR-482RF0IMFRRjoCCMsCN0
RRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVzv)q4:nRRLDNCHDR#1R"7Ra"&MRH0CCosl'HN5oCI0H8E&2RR""7RH&RMo0CCHs'lCNo5lMk_DOCDc_n*Rnc+kRMlC_ODdD_..*d2RR&"RW"&MRH0CCosl'HN5oC[&2RR"" RH&RMo0CCHs'lCNo50oC_8CM_b8C0ME5kOl_C_DDnnc*cRR+M_klODCD_*d.d+.RR,4nRb8C02E2R"&RX&"RR0HMCsoC'NHlo[C5+;42
RRRRRRRRRRRRoLCHRM
RRRRRRRRRzRR)4qvnRR:)4qvn7X4RR
RRRRRRRRRRRRRRFRbsl0RN5bR7>R=R_HMs_Co#25[,jRqRR=>D_FII8N8s5_#jR2,q=4R>FRDIN_I8_8s#254,.RqRR=>D_FII8N8s5_#.
2,RRRRRRRRRRRRRRRRRRRRRRRRRdRqRR=>D_FII8N8s5_#dR2,7qu)j>R=RIDF_8sN8#s_5,j2R)7uq=4R>FRDIN_s8_8s#254,uR7)Rq.=D>RFsI_Ns88_.#52S,
SSSSS7RRud)qRR=>D_FIs8N8s5_#dR2,W= R>sRI0M_C_,4nRpWBi>R=RiBp,uR7m>R=RksF0k_L#n_4#k5MlC_OD4D_n2,[,uR1m>R=RkIF0k_L#n_4#k5MlC_OD4D_n2,[2R;
RRRRRRRRRRRRRsRRF_k0s_Co#25[RR<=s0Fk_#Lk_#4n5lMk_DOCDn_4,R[2IMECRF5skC0_Mn_4R'=R4R'2CCD#R''Z;S
SSFSIks0_C#o_5R[2<I=RF_k0L_k#45n#M_klODCD_,4n[I2RERCM5kIF0M_C_R4n=4R''C2RDR#C';Z'
RRRRRRRR8CMRMoCC0sNC.Rz6R;
RCRRMo8RCsMCNR0Cz;..RRRR
CRRMo8RCsMCNR0Cz;cc
8CMRONsECH0Os0kCDRLF_O	s;Nl
-
----------------------F-M__sIOOEC	------------------------N

sHOE00COkRsCMsF_IE_OCRO	F)VRq)v_W)u_R
H#ObFlFMMC0)RXq.vdXR47RFRbs50R
RRRRRRRRm7uR:RRR0FkR8#0_FkDo;HORRRRRRRR
RRRRRRRRm1uR:RRR0FkR8#0_FkDo;HO
R
RRRRRRjRqRRRR:MRHR8#0_FkDo;HO
RRRRRRRRRq4R:RRRRHM#_08koDFH
O;RRRRRRRRqR.RRRR:H#MR0k8_DHFoOR;
RRRRRqRRdRRRRH:RM0R#8D_kFOoH;R
RRRRRRcRqRRRR:MRHR8#0_FkDo;HO
RRRRRRRRR7RR:RRRRHM#_08koDFH
O;RRRRRRRR7qu)jRR:H#MR0k8_DHFoOR;
RRRRR7RRu4)qRH:RM0R#8D_kFOoH;R
RRRRRRuR7)Rq.:MRHR8#0_FkDo;HO
RRRRRRRR)7uq:dRRRHM#_08koDFH
O;RRRRRRRR7qu)cRR:H#MR0k8_DHFoOR;
RRRRRWRRBRpiRH:RM0R#8D_kFOoH;RRRRRRRRR
RRRRRR RWRRRR:MRHR8#0_FkDo
HORRRRR2RR;
RRCRM8ObFlFMMC0O;
FFlbM0CMRqX)vXnc4R7RRsbF0
R5RRRRRRRR7RumRRR:FRk0#_08koDFHRO;RRRRR
RRRRRRRRRR1RumRRR:FRk0#_08koDFH
O;
RRRRRRRRRqjR:RRRRHM#_08koDFH
O;RRRRRRRRqR4RRRR:H#MR0k8_DHFoOR;
RRRRRqRR.RRRRH:RM0R#8D_kFOoH;R
RRRRRRdRqRRRR:MRHR8#0_FkDo;HO
RRRRRRRRRqcR:RRRRHM#_08koDFH
O;RRRRRRRRqR6RRRR:H#MR0k8_DHFoOR;
RRRRR7RRRRRRRH:RM0R#8D_kFOoH;R
RRRRRRuR7)Rqj:MRHR8#0_FkDo;HO
RRRRRRRR)7uq:4RRRHM#_08koDFH
O;RRRRRRRR7qu).RR:H#MR0k8_DHFoOR;
RRRRR7RRud)qRH:RM0R#8D_kFOoH;R
RRRRRRuR7)Rqc:MRHR8#0_FkDo;HO
RRRRRRRR)7uq:6RRRHM#_08koDFH
O;RRRRRRRRWiBpRRR:H#MR0k8_DHFoOR;RRRRRRRR
RRRRRWRR RRRRH:RM0R#8D_kFOoH
RRRRRRR2R;R
8CMRlOFbCFMM
0;VOkM0MHFRMVkOM_HHL05RL:RFCFDNRM2skC0s#MR0MsHo#RH
oLCHRM
RRHV5RL20MEC
RRRR0sCk5sM";"2
CRRD
#CRRRRskC0s"M5BDFk8FRM0lRHblDCCRM0AODF	qR)vQ3R#ER0CCRsNN8R8C8s#s#RC#oH0CCs8#RkHRMo0REC#CNlRFODON	R#ER0CqR)v2?";R
RCRM8H
V;CRM8VOkM_HHM0V;
k0MOHRFMo_C0C_M880CbEH5#x:CRR0HMCsoCR8;RCEb0RH:RMo0CCRs2skC0sHMRMo0CCHsR#N
PsLHNDlCRH#M_HRxC:MRH0CCos=R:R
j;LHCoMR
Rl_HM#CHxRR:=80CbER;
RRHV5x#HCRR<80CbE02RE
CMRRRRl_HM#CHxRR:=#CHx;R
RCRM8H
V;RCRs0MksRMlH_x#HCC;
Mo8RCC0_M88_CEb0;0
N0LsHkR0CoCCMsFN0sC_sb0FsR#:R0MsHoN;
0H0sLCk0RMoCC0sNFss_CsbF0VRFR_MFsOI_E	CORN:RsHOE00COkRsCHV#Rk_MOH0MH58sN8ss_C;o2
R--LHCoMDRLFRO	sRNlHDlbCMlC0HN0F#MRHNoMD0#
$RbCH_M0NNss$#RHRsNsN5$RjFR0RR62FHVRMo0CC
s;O#FM00NMR8IH0NE_s$sNRH:RMN0_s$sNRR:=5R4,.c,R,,RgR,4UR2dn;F
OMN#0M80RCEb0_sNsN:$RR0HM_sNsN:$R=4R5ncdU,4RUgR.,cnjg,jR.cRU,4cj.,4R6.
2;O#FM00NMRP8Hd:.RR0HMCsoCRR:=58IH04E-2n/d;F
OMN#0M80RHnP4RH:RMo0CC:sR=IR5HE80-/424
U;O#FM00NMRP8HURR:HCM0oRCs:5=RI0H8E2-4/
g;O#FM00NMRP8HcRR:HCM0oRCs:5=RI0H8E2-4/
c;O#FM00NMRP8H.RR:HCM0oRCs:5=RI0H8E2-4/
.;O#FM00NMRP8H4RR:HCM0oRCs:5=RI0H8E2-4/
4;
MOF#M0N0FRLFRD4:FRLFNDCM=R:RH58P>4RR;j2
MOF#M0N0FRLFRD.:FRLFNDCM=R:RH58P>.RR;j2
MOF#M0N0FRLFRDc:FRLFNDCM=R:RH58P>cRR;j2
MOF#M0N0FRLFRDU:FRLFNDCM=R:RH58P>URR;j2
MOF#M0N0FRLFnD4RL:RFCFDN:MR=8R5HnP4Rj>R2O;
F0M#NRM0LDFFd:.RRFLFDMCNRR:=5P8Hd>.RR;j2
F
OMN#0M80RHnP4dRUc:MRH0CCos=R:RC58b-0E442/ncdU;F
OMN#0M80RH4PUg:.RR0HMCsoCRR:=5b8C04E-24/Ug
.;O#FM00NMRP8HcnjgRH:RMo0CC:sR=8R5CEb0-/42cnjg;F
OMN#0M80RHjP.c:URR0HMCsoCRR:=5b8C04E-2j/.c
U;O#FM00NMRP8H4cj.RH:RMo0CC:sR=8R5CEb0-/424cj.;F
OMN#0M80RH4P6.RR:HCM0oRCs:5=R80CbE2-4/.64;O

F0M#NRM0LDFF6R4.:FRLFNDCM=R:RH58P.64Rj>R2O;
F0M#NRM0LDFF4cj.RL:RFCFDN:MR=8R5HjP4.>cRR;j2
MOF#M0N0FRLFjD.c:URRFLFDMCNRR:=5P8H.UjcRj>R2O;
F0M#NRM0LDFFcnjgRL:RFCFDN:MR=8R5HjPcg>nRR;j2
MOF#M0N0FRLF4DUg:.RRFLFDMCNRR:=5P8HU.4gRj>R2O;
F0M#NRM0LDFF4UndcRR:LDFFCRNM:5=R84HPncdURj>R2
;
O#FM00NMRl#k_8IH0:ERR0HMCsoCRR:=Apmm 'qhb5F#LDFF4+2RRmAmph q'#bF5FLFDR.2+mRAmqp hF'b#F5LF2DcRA+Rm mpqbh'FL#5FUFD2RR+Apmm 'qhb5F#LDFF4;n2
MOF#M0N0kR#lC_8bR0E:MRH0CCos=R:R-6RRm5Amqp hF'b#F5LF4D6.+2RRmAmph q'#bF5FLFD.4jc+2RRmAmph q'#bF5FLFDc.jU+2RRmAmph q'#bF5FLFDgcjn+2RRmAmph q'#bF5FLFDgU4.;22
F
OMN#0MI0R_FOEH_OCI0H8ERR:HCM0oRCs:I=RHE80_sNsN#$5kIl_HE802O;
F0M#NRM0IE_OFCHO_b8C0:ERR0HMCsoCRR:=80CbEs_Ns5N$#_klI0H8E
2;O#FM00NMRO8_EOFHCH_I8R0E:MRH0CCos=R:R8IH0NE_s$sN5l#k_b8C0;E2
MOF#M0N0_R8OHEFO8C_CEb0RH:RMo0CC:sR=CR8b_0ENNss$k5#lC_8b20E;O

F0M#NRM0IH_I8_0EM_klODCD#RR:HCM0oRCs:5=RI0H8E2-4/OI_EOFHCH_I8R0E+;R4
MOF#M0N0_RI80CbEk_MlC_ODRD#:MRH0CCos=R:RC58b-0E4I2/_FOEH_OC80CbERR+4
;
O#FM00NMRI8_HE80_lMk_DOCD:#RR0HMCsoCRR:=58IH04E-2_/8OHEFOIC_HE80R4+R;F
OMN#0M80R_b8C0ME_kOl_C#DDRH:RMo0CC:sR=8R5CEb0-/428E_OFCHO_b8C0+ERR
4;
MOF#M0N0_RI#CHxRH:RMo0CC:sR=_RII0H8Ek_MlC_ODRD#*_RI80CbEk_MlC_OD;D#
MOF#M0N0_R8#CHxRH:RMo0CC:sR=_R8I0H8Ek_MlC_ODRD#*_R880CbEk_MlC_OD;D#
F
OMN#0ML0RF_FD8RR:LDFFCRNM:5=R8H_#x-CRR#I_HRxC<j=R2O;
F0M#NRM0LDFF_:IRRFLFDMCNRR:=M5F0LDFF_;82
F
OMN#0MO0REOFHCH_I8R0E:MRH0CCos=R:Rm5Amqp hF'b#F5LF8D_2RR*8E_OFCHO_8IH0RE2+AR5m mpqbh'FL#5F_FDI*2RROI_EOFHCH_I820E;F
OMN#0MO0REOFHCC_8bR0E:MRH0CCos=R:Rm5Amqp hF'b#F5LF8D_2RR*8E_OFCHO_b8C0RE2+AR5m mpqbh'FL#5F_FDI*2RROI_EOFHCC_8b20E;F
OMN#0MI0RHE80_lMk_DOCD:#RR0HMCsoCRR:=5mAmph q'#bF5FLFD2_8RI*5HE80-/428E_OFCHO_8IH0RE2+AR5m mpqbh'FL#5F_FDI*2RRH5I8-0E4I2/_FOEH_OCI0H8E+2RR
4;O#FM00NMRb8C0ME_kOl_C#DDRH:RMo0CC:sR=AR5m mpqbh'FL#5F_FD8*2R5b8C04E-2_/8OHEFO8C_CEb02RR+5mAmph q'#bF5FLFD2_IR5*R80CbE2-4/OI_EOFHCC_8b20ER4+R;$
0bFCRkL0_k_#40C$bRRH#NNss$8R5CEb0_lMk_DOCD4#-RI8FMR0FjI,RHE80_lMk_DOCD4#-RI8FMR0FjF2RV0R#8F_Do;HO
o#HMRNDs0Fk_#Lk4RR:F_k0L4k#_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFR8s_FRk05bHMk00RFsR0H0-#N#0C2H
#oDMNRkIF0k_L#:4RR0Fk_#Lk4$_0b
C;0C$bR0Fk_#Lk.$_0bHCR#sRNsRN$5b8C0ME_kOl_C#DD-84RF0IMF,RjRI.*HE80_lMk_DOCD4#+RI8FMR0FjF2RV0R#8F_Do;HO
o#HMRNDs0Fk_#Lk.RR:F_k0L.k#_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFR8s_FRk05bHMk00RFsR0H0-#N#0C2H
#oDMNRkIF0k_L#:.RR0Fk_#Lk.$_0b
C;0C$bR0Fk_#Lkc$_0bHCR#sRNsRN$5b8C0ME_kOl_C#DD-84RF0IMF,RjRIc*HE80_lMk_DOCDd#+RI8FMR0FjF2RV0R#8F_Do;HO
o#HMRNDs0Fk_#LkcRR:F_k0Lck#_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFR8s_FRk05bHMk00RFsR0H0-#N#0C2H
#oDMNRkIF0k_L#:cRR0Fk_#Lkc$_0b
C;0C$bR0Fk_#LkU$_0bHCR#sRNsRN$5b8C0ME_kOl_C#DD-84RF0IMF,RjRIU*HE80_lMk_DOCD(#+RI8FMR0FjF2RV0R#8F_Do;HO
o#HMRNDs0Fk_#LkURR:F_k0LUk#_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFR8s_FRk05bHMk00RFsR0H0-#N#0C2H
#oDMNRkIF0k_L#:URR0Fk_#LkU$_0b
C;0C$bRsbNH_0$LUk#_b0$C#RHRsNsN5$R80CbEk_MlC_OD-D#4FR8IFM0RRj,I0H8Ek_MlC_OD-D#4FR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNRNsbs$H0_#LkURR:bHNs0L$_k_#U0C$b;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RV_Rs80FkRM5HbRk000FRs#H-0CN0##2
HNoMDbRIN0sH$k_L#:URRsbNH_0$LUk#_b0$C0;
$RbCF_k0L4k#n$_0bHCR#sRNsRN$5b8C0ME_kOl_C#DD-84RF0IMF,RjR*4nI0H8Ek_MlC_OD+D#486RF0IMF2RjRRFV#_08DHFoO#;
HNoMDFRskL0_kn#4RF:RkL0_kn#4_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFR8s_FRk05bHMk00RFsR0H0-#N#0C2H
#oDMNRkIF0k_L#R4n:kRF0k_L#_4n0C$b;$
0bbCRN0sH$k_L#_4n0C$bRRH#NNss$8R5CEb0_lMk_DOCD4#-RI8FMR0Fj.,R*8IH0ME_kOl_C#DD+84RF0IMF2RjRRFV#_08DHFoO#;
HNoMDbRsN0sH$k_L#R4n:NRbs$H0_#Lk40n_$;bCRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$FsVR_k8F0HR5M0bkRR0F0-sH#00NC
#2#MHoNIDRbHNs0L$_kn#4Rb:RN0sH$k_L#_4n0C$b;$
0bFCRkL0_k.#d_b0$C#RHRsNsN5$R80CbEk_MlC_OD-D#4FR8IFM0RRj,dI.*HE80_lMk_DOCDd#+4FR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNRksF0k_L#Rd.:kRF0k_L#_d.0C$b;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFVsF_8k50RHkMb0FR0RH0s-N#002C#
o#HMRNDI0Fk_#Lkd:.RR0Fk_#Lkd0._$;bC
b0$CNRbs$H0_#Lkd0._$RbCHN#Rs$sNRC58b_0EM_klODCD#R-48MFI0jFR,*RcI0H8Ek_MlC_OD+D#dFR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNRNsbs$H0_#Lkd:.RRsbNH_0$Ldk#.$_0bRC;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RV_Rs80FkRM5HbRk000FRs#H-0CN0##2
HNoMDbRIN0sH$k_L#Rd.:NRbs$H0_#Lkd0._$;bC
o#HMRNDs0Fk_RCM:0R#8F_Do_HOP0COF8s5CEb0_lMk_DOCD4#-RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-C-RMDNLCV#RF0sRs#H-0CN0#H
#oDMNRkIF0M_CR#:R0D8_FOoH_OPC05Fs80CbEk_MlC_OD-D#4FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--CLMNDRC#VRFs0-sH#00NC##
HNoMDsRI0M_CR#:R0D8_FOoH_OPC05Fs80CbEk_MlC_OD-D#4FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--I0sHCMRCNCLD#FRVsNRCOsERFFIRVqR)vCROD
D##MHoNHDRMC_soRR:#_08DHFoOC_POs0F58IH0dE+6FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-#RkC08RFCRso0H#C7sRQ
hR#MHoNsDRF_k0sRCo:0R#8F_Do_HOP0COFIs5HE80+Rd68MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-k-R#RC80sFRC#oH0RCs7amz
o#HMRNDI0Fk_osCR#:R0D8_FOoH_OPC05FsI0H8E6+dRI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--k8#CRR0FsHCo#s0CRz7maH
#oDMNRksF0C_so:4RR8#0_oDFHPO_CFO0sH5I8-0E4FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--k8#CRR0FOFEF#LCRCC0IC7MRQNhRMF8Rkk0b0VRFRFADO)	Rq#v
HNoMDNRs8C_soRR:#_08DHFoOC_POs0F58N8s8IH04E-RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RCk#8FR0RosCHC#0sqR)7
7)#MHoNIDRNs8_C:oRR8#0_oDFHPO_CFO0s85N8HsI8-0E4FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-#RkC08RFCRso0H#CWsRq)77
o#HMRNDD_FIs8N8sRR:#_08DHFoOC_POs0F5R4d8MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--s8N8sHRL0H#RM0bkRR0F)RqvODCD#cR5R0LH#CRsJskHC
82#MHoNDDRFII_Ns88R#:R0D8_FOoH_OPC05Fs48dRF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-I-RNs88R0LH#MRHbRk00)FRqOvRC#DDRR5cL#H0RJsCkCHs8#2
HNoMDqR)7_7)0Rlb:0R#8F_Do_HOP0COFNs58I8sHE80-84RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-k-R#RC80bFRHDbCHRMC)7q7)H
#oDMNR7Wq70)_l:bRR8#0_oDFHPO_CFO0s85N8HsI8-0E4FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-#RkC08RFHRbbHCDMWCRq)77
o#HMRND7_Qh0Rlb:0R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RCk#8FR0RbbHCMDHCQR7hH
#oDMNR_W 0Rlb:0R#8F_Do;HORRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-#RkC08RFHRbbHCDMWCR H
#oDMNRNs_8_8ssRCo:0R#8F_Do_HOP0COFNs58I8sHE80-84RF0IMF2Rj;-
-R8CMRFLDOs	RNHlRlCbDl0CMNF0HMHR#oDMN#-
-RoLCH#MRCODC0NRsllRHblDCCNM00MHFRo#HM#ND
MVkOF0HMCRo0k_Mlc_n5b8C0RE:HCM0o2CsR0sCkRsMHCM0oRCsHP#
NNsHLRDCPRND:MRH0CCos=R:R
j;LHCoMR
RPRND:8=RCEb0/;nc
HRRV5R580CbEFRl8cRn2RR>cRU20MEC
RRRRDPNRR:=PRND+;R4
CRRMH8RVR;
R0sCkRsMP;ND
8CMR0oC_lMk_;nc
MVkOF0HMCRo0C_DVP0FCds_.C58bR0E:MRH0CCoss2RCs0kMMRH0CCos#RH
oLCHRM
R0sCk5sM80CbEFRl8cRn2C;
Mo8RCD0_CFV0P_Csd
.;VOkM0MHFR0oC_VDC0CFPsC58bR0E:MRH0CCosl;RN:GRR0HMCsoC2CRs0MksR0HMCsoCR
H#PHNsNCLDRDPNRH:RMo0CC:sR=;Rj
oLCHRM
RRHV5b8C0-ERRGlNRR>=j02RE
CMRRRRPRND:8=RCEb0Rl-RN
G;RDRC#RC
RPRRN:DR=CR8b;0E
CRRMH8RVR;
R0sCk5sMP2ND;M
C8CRo0C_DVP0FC
s;VOkM0MHFR0oC_lMk_5d.80CbERR:HCM0o2CsR0sCkRsMHCM0oRCsHP#
NNsHLRDCPRND:MRH0CCos=R:R
j;LHCoMR
RH5VR80CbE=R<RRcUNRM880CbERR>4Rn20MEC
RRRRNRPD=R:R
4;RMRC8VRH;R
RskC0sPMRN
D;CRM8o_C0M_kld
.;VOkM0MHFR0oC_lMk_54n80CbERR:HCM0o2CsR0sCkRsMHCM0oRCsHP#
NNsHLRDCPRND:MRH0CCos=R:R
j;LHCoMR
RH5VR80CbE=R<RR4nNRM880CbERR>j02RE
CMRRRRRDPNRR:=4R;
R8CMR;HV
sRRCs0kMNRPDC;
Mo8RCM0_k4l_nO;
F0M#NRM0M_klODCD_Rnc:MRH0CCos=R:R0oC_lMk_5nc80CbE
2;O#FM00NMRVDC0CFPs._dRH:RMo0CC:sR=CRo0C_DVP0FCds_.C58b20E;F
OMN#0MM0RkOl_C_DDd:.RR0HMCsoCRR:=o_C0M_kldD.5CFV0P_Csd;.2
MOF#M0N0CRDVP0FC4s_nRR:HCM0oRCs:o=RCD0_CFV0P5CsD0CVFsPC_,d.R2d.;F
OMN#0MM0RkOl_C_DD4:nRR0HMCsoCRR:=o_C0M_kl4Dn5CFV0P_Cs4;n2
$
0bFCRkL0_k0#_$_bCnRc#HN#Rs$sNRk5MlC_ODnD_cFR8IFM0RRj,I0H8ER-48MFI0jFR2VRFR8#0_oDFH
O;0C$bR0Fk_#Lk_b0$C._d##RHRsNsN5$RM_klODCD_Rd.8MFI0jFR,HRI8-0E4FR8IFM0RRj2F#VR0D8_FOoH;$
0bFCRkL0_k0#_$_bC4Rn#HN#Rs$sNRk5MlC_OD4D_nFR8IFM0RRj,I0H8ER-48MFI0jFR2VRFR8#0_oDFH
O;#MHoNsDRF_k0L_k#nRc#:kRF0k_L#$_0bnC_cR#;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RVFR8k50RHkMb0FR0RH0s-N#002C#
o#HMRNDI0Fk_#Lk_#ncRF:RkL0_k0#_$_bCn;c#RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$F8VRFRk05bHMk00RFsR0H0-#N#0C2H
#oDMNRksF0k_L#._d#RR:F_k0L_k#0C$b_#d.;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFV80FkRM5HbRk000FRs#H-0CN0##2
HNoMDFRIkL0_kd#_.:#RR0Fk_#Lk_b0$C._d##;
HNoMDFRskL0_k4#_n:#RR0Fk_#Lk_b0$Cn_4#R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFRk8F0HR5M0bkRR0F0-sH#00NC
#2#MHoNIDRF_k0L_k#4Rn#:kRF0k_L#$_0b4C_n
#;#MHoNsDRF_k0C#M_R#:R0D8_FOoH_OPC05FsM_klODCD_Rnc8MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-MRCNCLD#FRVssR0H0-#N#0C
o#HMRNDI0Fk__CM#RR:#_08DHFoOC_POs0F5lMk_DOCDc_nRI8FMR0Fj
2;#MHoNsDRF_k0CdM_.RR:#_08DHFoO#;
HNoMDFRIkC0_M._dR#:R0D8_FOoH;H
#oDMNRksF0M_C_R4n:0R#8F_Do;HO
o#HMRNDI0Fk__CM4:nRR8#0_oDFH
O;#MHoNIDRsC0_MR_#:0R#8F_Do_HOP0COFMs5kOl_C_DDn8cRF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RHIs0CCRMDNLCV#RFCsRNROEsRFIF)VRqOvRC#DD
o#HMRNDI_s0CdM_.RR:#_08DHFoO#;
HNoMDsRI0M_C_R4n:0R#8F_Do;HO
o#HMRNDHsM_C#o_R#:R0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--k8#CRR0FsHCo#s0CRh7QRH
#oDMNRksF0C_soR_#:0R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-#RkC08RFCRso0H#C7sRm
za#MHoNIDRF_k0s_Co#RR:#_08DHFoOC_POs0F58IH04E-RI8FMR0FjR2;R#R
HNoMDNRs8C_soR_#:0R#8F_Do_HOP0COFNs58I8sHE80-84RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-k-R#RC80sFRC#oH0RCsq)77
o#HMRNDI_N8s_Co#RR:#_08DHFoOC_POs0F58N8s8IH04E-RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RCk#8FR0RosCHC#0s7Rq7#)
HNoMDFRDIN_s8_8s#RR:#_08DHFoOC_POs0F586RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-N-R8R8sL#H0RbHMk00RFqR)vCRODRD#5LcRHR0#skCJH8sC2H
#oDMNRIDF_8IN8#s_R#:R0D8_FOoH_OPC05Fs6FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-8RN8LsRHR0#HkMb0FR0Rv)qRDOCD5#RcHRL0s#RCHJks2C8
R--CRM8#CCDOs0RNHlRlCbDl0CMNF0HMHR#oDMN#0
N0LsHkR0C\N3slV_FV0#C\RR:#H0sM
o;
oLCHRM
Rdzc:VRHRN5s8_8ss2CoRMoCC0sNC-R-RMoCC0sNCDRLFRO	s
NlRRRR-Q-RV8RN8HsI8R0E<EROFCHO_8IH0NER#o#HMjR''FR0RkkM#RC8L#H0
RRRRRzjRH:RVNR58I8sHE80R4=R2CRoMNCs0SC
RRRRD_FIs8N8s=R<Rj"jjjjjjjjjj"jjRs&RNs8_Cjo52S;
RRRRD_FII8N8s=R<Rj"jjjjjjjjjj"jjRI&RNs8_Cjo52S;
CRM8oCCMsCN0R;zj
RRRRRz4RH:RVNR58I8sHE80R.=R2CRoMNCs0SC
SIDF_8sN8<sR=jR"jjjjjjjjj"jjRs&RNs8_C4o5RI8FMR0Fj
2;SRRRRIDF_8IN8<sR=jR"jjjjjjjjj"jjRI&RNs8_C4o5RI8FMR0Fj
2;S8CMRMoCC0sNC4Rz;R
RR.RzRRR:H5VRNs88I0H8ERR=do2RCsMCN
0CSFSDIN_s8R8s<"=Rjjjjjjjjj"jjRs&RNs8_C.o5RI8FMR0Fj
2;SRRRRIDF_8IN8<sR=jR"jjjjjjjjjRj"&NRI8C_soR5.8MFI0jFR2S;
CRM8oCCMsCN0R;z.
RRRRRzdRH:RVNR58I8sHE80Rc=R2CRoMNCs0SC
SIDF_8sN8<sR=jR"jjjjjjjjj&"RR8sN_osC58dRF0IMF2Rj;R
SRDRRFII_Ns88RR<="jjjjjjjj"jjRI&RNs8_Cdo5RI8FMR0Fj
2;S8CMRMoCC0sNCdRz;R
RRcRzRRR:H5VRNs88I0H8ERR=6o2RCsMCN
0CSRRRRIDF_8sN8<sR=jR"jjjjjjjj"RR&s_N8s5CocFR8IFM0R;j2
RSRRFRDIN_I8R8s<"=Rjjjjjjjjj&"RR8IN_osC58cRF0IMF2Rj;C
SMo8RCsMCNR0Cz
c;RRRRzR6R:VRHR85N8HsI8R0E=2RnRMoCC0sNCR
SRDRRFsI_Ns88RR<="jjjjjjjj&"RR8sN_osC586RF0IMF2Rj;S
SD_FII8N8s=R<Rj"jjjjjjRj"&NRI8C_soR568MFI0jFR2S;
CRM8oCCMsCN0R;z6
RRRRRznRH:RVNR58I8sHE80R(=R2CRoMNCs0SC
RRRRD_FIs8N8s=R<Rj"jjjjjj&"RR8sN_osC58nRF0IMF2Rj;S
SD_FII8N8s=R<Rj"jjjjjj&"RR8IN_osC58nRF0IMF2Rj;C
SMo8RCsMCNR0Cz
n;RRRRzR(R:VRHR85N8HsI8R0E=2RURMoCC0sNCR
SRDRRFsI_Ns88RR<="jjjj"jjRs&RNs8_C(o5RI8FMR0Fj
2;SFSDIN_I8R8s<"=RjjjjjRj"&NRI8C_soR5(8MFI0jFR2S;
CRM8oCCMsCN0R;z(
RRRRRzURH:RVNR58I8sHE80Rg=R2CRoMNCs0SC
RRRRD_FIs8N8s=R<Rj"jj"jjRs&RNs8_CUo5RI8FMR0Fj
2;SFSDIN_I8R8s<"=Rjjjjj&"RR8IN_osC58URF0IMF2Rj;C
SMo8RCsMCNR0Cz
U;RRRRzRgR:VRHR85N8HsI8R0E=jR42CRoMNCs0SC
RRRRD_FIs8N8s=R<Rj"jjRj"&NRs8C_soR5g8MFI0jFR2S;
SIDF_8IN8<sR=jR"j"jjRI&RNs8_Cgo5RI8FMR0Fj
2;S8CMRMoCC0sNCgRz;R
RR4Rzj:RRRRHV58N8s8IH0=ERR244RMoCC0sNCR
SRDRRFsI_Ns88RR<="jjj"RR&s_N8s5Co48jRF0IMF2Rj;S
SD_FII8N8s=R<Rj"jj&"RR8IN_osC5R4j8MFI0jFR2S;
CRM8oCCMsCN0Rjz4;R
RR4Rz4:RRRRHV58N8s8IH0=ERR24.RMoCC0sNCR
SRDRRFsI_Ns88RR<=""jjRs&RNs8_C4o54FR8IFM0R;j2
DSSFII_Ns88RR<=""jjRI&RNs8_C4o54FR8IFM0R;j2
MSC8CRoMNCs0zCR4
4;RRRRzR4.RH:RVNR58I8sHE80R4=Rdo2RCsMCN
0CSRRRRIDF_8sN8<sR=jR''RR&s_N8s5Co48.RF0IMF2Rj;S
SD_FII8N8s=R<R''jRI&RNs8_C4o5.FR8IFM0R;j2
MSC8CRoMNCs0zCR4
.;RRRRzR4dRH:RVNR58I8sHE80R4>Rdo2RCsMCN
0CSRRRRIDF_8sN8<sR=NRs8C_sod54RI8FMR0Fj
2;SRRRRIDF_8IN8<sR=NRI8C_sod54RI8FMR0Fj
2;S8CMRMoCC0sNC4Rzd
;
RRRR-Q-RV8R5HsM_CRo2sHCo#s0CRh7QRHk#MBoRpRi
RzRR4RcR:VRHRH58MC_soo2RCsMCN
0CRRRRRRRRbOsFCR##5iBp,QR7hL2RCMoH
RRRRRRRRRRRRRHV5iBpR'=R4N'RMB8RpCi'P0CM2ER0CRM
RRRRRRRRRRRRRHRRMC_so=R<Rj5"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jjR7&RQ;h2
RRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMRFbsO#C#;C
SMo8RCsMCNR0Cz;4c
RRRR6z4RRR:H5VRMRF08_HMs2CoRMoCC0sNCR
RRRRRRRRRRMRH_osCRR<=5j"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjRj"&QR7h
2;S8CMRMoCC0sNC4Rz6
;
RRRR-Q-RVsR580Fk_osC2CRso0H#C)sR_z7ma#RkHRMo)B_mpRi
RzRR48nsFRk0RH:RVsR580Fk_osC2CRoMNCs0RC
RRRRRbRRsCFO#5#R)B_mpRi,s0Fk_osC4L2RCMoH
RRRRRRRRRRRRRHV5m)_BRpi=4R''MRN8_R)miBp'CCPMR020MEC
RRRRRRRRRRRRRRRR7)_mRza<s=RF_k0s4Co;R
RRRRRRRRRRMRC8VRH;R
RRRRRRMRC8sRbF#OC#R;
RRRRRCRRMo8RCsMCNR0Czs4n80Fk;R
RR4Rz(Fs8kR0R:VRHRF5M08RsF_k0s2CoRMoCC0sNCR
RRRRRRRRRR_R)7amzRR<=s0Fk_osC4S;
CRM8oCCMsCN0R(z4sk8F0
;
Snz4Ik8F0:RRRRHV5FI8ks0_CRo2oCCMsCN0
RRRRRRRRFbsO#C#R_5WmiBp,FRIks0_CRo2LHCoMR
RRRRRRRRRRVRHR_5WmiBpR'=R4N'RMW8R_pmBiP'CC2M0RC0EMR
RRRRRRRRRRRRRR_RW7amzRR<=I0Fk_osC58IH04E-RI8FMR0Fj
2;RRRRRRRRRRRRCRM8H
V;RRRRRRRRCRM8bOsFC;##
RRRRRRRR8CMRMoCC0sNC4RznFI8k
0;RRRRzI4(80FkRRR:H5VRMRF0Ik8F0C_soo2RCsMCN
0CRRRRRRRRRRRRWm_7z<aR=FRIks0_CIo5HE80-84RF0IMF2Rj;C
SMo8RCsMCNR0CzI4(80Fk;R

R-RR-VRQRN5s8_8ss2CoRosCHC#0sqR)7R7)kM#HoBRmpRi
RzRR4RnsRH:RVsR5Ns88_osC2CRoMNCs0-C
-RRRRRRRRFbsO#C#RB5mpRi,)7q7)L2RCMoH
R--RRRRRRRRRHRRVmR5BRpi=4R''MRN8BRmpCi'P0CM2ER0C-M
-RRRRRRRRRRRRRRRR8sN_osCRR<=)7q7)85N8HsI8-0E4FR8IFM0R;j2
R--RRRRRRRRRCRRMH8RV-;
-RRRRRRRR8CMRFbsO#C#;-
-S8CMRMoCC0sNC4Rzn
s;-R-RR4Rz(:sRRRHV50MFR8sN8ss_CRo2oCCMsCN0
RRRRRRRRRRRR8sN_osCRR<=)7q7)S;
CRM8oCCMsCN0Rnz4s
;
SR--Q5VRI8N8sC_sos2RC#oH0RCsW7q7)#RkHRMoWB_mpRi
RzRR4RnIRH:RVIR5Ns88_osC2CRoMNCs0RC
RRRRRbRRsCFO#5#RB,piR7Wq7R)2LHCoMR
RRRRRRRRRRVRHRp5BiRR='R4'NRM8B'piCMPC002RE
CMRRRRRRRRRRRRRRRRI_N8sRCo<W=Rq)7758N8s8IH04E-RI8FMR0Fj
2;RRRRRRRRRRRRCRM8H
V;RRRRRRRRCRM8bOsFC;##
MSC8CRoMNCs0zCR4;nI
RRRR(z4IRR:H5VRMRF0I8N8sC_soo2RCsMCN
0CRRRRRRRRRRRRI_N8sRCo<W=Rq)77;C
SMo8RCsMCNR0CzI4(;R

R-RR-GR 0RsNDHFoOFRVskR7NbDRFRs0OCN#
-S-MRF0M8CCCV8RFMsRFI_s_COEOS	
-s-zC:oRRFbsO#C#5iBp2CRLo
HM-R-SRRHV5iBp'  ehNaRMB8Rp=iRR''42ER0C-M
-RSRRh7Q_b0lRR<=7;Qh
S--R)RRq)77_b0lRR<=)7q7)-;
-RSRR7Wq70)_l<bR=qRW7;7)
S--RWRR l_0b=R<R;W 
S--RMRC8VRH;-
-S8CMRFbsO#C#;S

-Q-RVCR)Nq8R8C8s#=#RRHWs0qCR8C8s#R#,LN$b#7#RQ0hRFkRF00bkRRHVWH R#MRCNCLD8z
SlRkG:sRbF#OC# 5W_b0l,qR)7_7)0,lbR7Wq70)_lRb,7_Qh0,lbRksF0C_soS2
RCRLo
HM-R-SRHRRVWR5q)77_b0lR)=Rq)77_b0lR8NMR_W 0Rlb=4R''02RE
CM-S-SRFRsks0_CRo4<7=RQ0h_l
b;-S-SCCD#
RSSRksF0C_so<4R=FRsks0_CIo5HE80-84RF0IMF2Rj;-
-SMSC8VRH;C
SMb8RsCFO#
#;SRRRRR
RR-R-RMtCC0sNCER0CqR)vCRODRD#NRM8#CCDOD0RFOoHRsVFRv)qA_4n114_4z
S4:URRRHV5FOEH_OCI0H8ERR=4o2RCsMCN
0CSSRRRzRRO:E	RRHV58N8s8IH0>ERR24cRMoCC0sNCR
RRRRRRORkD:	RRFbsO#C#5iBp2R
RRRRRRLRRCMoH
RRRRRRRRHRRVBR5pCi'P0CMR8NMRiBpR'=R4R'20MEC
RRRRRRRRRRRRNs_8_8ss5CoNs88I0H8ER-48MFI04FRc<2R=qR)757)Ns88I0H8ER-48MFI04FRc
2;RRRRRRRRRMRC8VRH;R
RRRRRRMRC8sRbF#OC#ORkD
	;SCRRMo8RCsMCNR0Cz	OE;R
RRzRS4:gRRsVFRHHRM8R5CEb0_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNC-
S-VRQR85N8HsI8R0E>cR42CRMC08RFsROCCN0RHIs0CCRMDNLCMRN8kRF00bkRNCMLRDC#CCDOD0RFOoH
RRRRRRRR.SzjRR:H5VRNs88I0H8ERR>4Rc2oCCMsCN0
-S-RGVHRsVFRDONDdR4U,U(RD#CCRO0F0VRs0H#NR0CMRF0LMCHoCRso0H#C8sC
SSSSksF0M_C5RH2<'=R4I'RERCM5Ns_8_8ss5CoNs88I0H8ER-48MFI04FRc=2RRRH2CCD#R''j;S
SSFSIkC0_M25HRR<='R4'IMECRN5I8C_so85N8HsI8-0E4FR8IFM0R24cRH=R2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0CHM52=R<RRW IMECRN5I8C_so85N8HsI8-0E4FR8IFM0R24cRH=R2DRC#'CRj
';RRRRRRRRS8CMRMoCC0sNC.RzjS;
-Q-RVNR58I8sHE80RR<=4Rc2MIFRsCH0RNCMLRDCFFsRkk0b0MRCNCLDRD#CCRO0DHFoOCRMC88C
RRSRSRRzR.4:VRHR85N8HsI8R0E<4=Rco2RCsMCN
0CSSSSs0Fk_5CMH<2R=4R''S;
SISSF_k0CHM52=R<R''4;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R R;
RRRRRSRRCRM8oCCMsCN0R4z.;-
S-CRtMNCs00CRE)CRqOvRC#DDR8NMRH0s-N#00
C#RRRRRRRRS.z.RV:RF[sRRRHM58IH0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CRRRRRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FAVR)_qv4Undc7X4RD:RNDLCRRH#";W"
RRRRRRRRRRRRRRRRoLCHRM
RRRRRRRRRSRRAv)q_d4nU4cX7RR:)Aqv41n_44_1
RSRRRRRRRRRRFRbsl0RN5bR75Qqj=2R>MRH_osC5,[2R7q7)=qR>FRDIN_I858s48dRF0IMF2Rj,QR7A>R=R""j,7Rq7R)A=D>RFsI_Ns885R4d8MFI0jFR2S,
S SSh=qR>4R''1,R1R)q='>RjR',WR q=I>RsC0_M25H,pRBi=qR>pRBi ,Rh=AR>4R''1,R1R)A='>RjR',WR A='>RjR',BApiRR=>B,pi
SSSRRRR75mqj=2R>FRIkL0_k5#4H2,[,mR7A25jRR=>s0Fk_#Lk4,5H[;22
R
RRRRRRRRRRRRRRFRsks0_C[o52=R<RksF0k_L#H45,R[2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;S
SSFSIks0_C[o52=R<RkIF0k_L#H45,RK2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRCRSMo8RCsMCNR0Cz;..
RRRRCRSMo8RCsMCNR0Cz;4g
RRRR8CMRMoCC0sNC4RzUR;RRRR
RRRRRR
RR-R-RMtCC0sNCER0CqR)vCRODRD#NRM8#CCDOD0RFOoHRsVFRv)qA_4n11._.z
S.:dRRRHV5FOEH_OCI0H8ERR=.o2RCsMCN
0CSzRRORE	:VRHR85N8HsI8R0E>dR42CRoMNCs0RC
RRRRRkRRORD	:sRbF#OC#p5BiR2
RRRRRRRRLHCoMR
RRRRRRRRRH5VRB'piCMPC0MRN8pRBiRR='24'RC0EMR
RRRRRRRRRR_RsNs88_osC58N8s8IH04E-RI8FMR0F4Rd2<)=Rq)7758N8s8IH04E-RI8FMR0F4;d2
RRRRRRRRCRRMH8RVR;
RRRRRCRRMb8RsCFO#k#RO;D	
RSRCRM8oCCMsCN0REzO	R;
RSRRzR.c:FRVsRRHH5MR80CbEk_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0SC
-Q-RVNR58I8sHE80R4>RdM2RCRC80OFRs0CNCsRIHR0CCLMNDNCRMF8Rkk0b0MRCNCLDRD#CCRO0DHFoOR
RRRRRRzRS.:6RRRHV58N8s8IH0>ERR24dRMoCC0sNC-
S-HRVGFRVsNROD4DRd(UU,CR#D0CORRFV0#sH0CN0R0MFRHLCMsoRC#oH0CCs8R
RRRRRRRRRRRRRRFRskC0_M25HRR<='R4'IMECR_5sNs88_osC58N8s8IH04E-RI8FMR0F4Rd2=2RHR#CDCjR''S;
SISSF_k0CHM52=R<R''4RCIEMIR5Ns8_CNo58I8sHE80-84RF0IMFdR42RR=HC2RDR#C';j'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RWRCIEMIR5Ns8_CNo58I8sHE80-84RF0IMFdR42RR=HC2RDR#C';j'
RRRRRRRRMSC8CRoMNCs0zCR.
6;SR--Q5VRNs88I0H8E=R<R24dRRMFI0sHCMRCNCLDRRFsFbk0kC0RMDNLCCR#D0CORoDFHMORCCC88S
RRRRRSnz.RH:RVNR58I8sHE80RR<=4Rd2oCCMsCN0
RSRRRRRRRRRRFRskC0_M25HRR<=';4'
SSSSkIF0M_C5RH2<'=R4
';RRRRRRRRRRRRRRRRI_s0CHM52=R<R;W 
RRRRRRRRMSC8CRoMNCs0zCR.
n;SR--tCCMsCN0RC0ERv)qRDOCDN#RM08Rs#H-0CN0#R
RRRRRRzRS.:(RRsVFRH[RMIR5HE80_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNCR
RRRRRRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqA)v4_Ug..X7RR:DCNLD#RHR""W;R
RRRRRRRRRRRRRRCRLo
HMRRRRRRRRRRRRSqA)v4_Ug..X7RR:)Aqv41n_.._1
RSRRRRRRRRRRFRbsl0RN5bR7RQq=H>RMC_so*5.[R+48MFI0.FR*,[2R7q7)=qR>FRDIN_I858s48.RF0IMF2Rj,QR7A>R=Rj"j"q,R7A7)RR=>D_FIs8N8s.54RI8FMR0Fj
2,SRSSR RRh=qR>4R''1,R1R)q='>RjR',WR q=I>RsC0_M25H,pRBi=qR>pRBi ,Rh=AR>4R''1,R1R)A='>RjR',WR A='>RjR',BApiRR=>B,pi
SSSRRRR75mq4=2R>FRIkL0_k5#.H*,.[2+4,mR7q25jRR=>I0Fk_#Lk.,5H.2*[,mR7A254RR=>s0Fk_#Lk.,5H.+*[4R2,75mAj=2R>FRskL0_k5#.H.,R*2[2;R
RRRRRRRRRRRRRRFRsks0_C.o5*R[2<s=RF_k0L.k#5.H,*R[2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRsks0_C.o5*4[+2=R<RksF0k_L#H.5,[.*+R42IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;S
SSFSIks0_C.o5*R[2<I=RF_k0L.k#5.H,*R[2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRIks0_C.o5*4[+2=R<RkIF0k_L#H.5,[.*+R42IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R

RRRRRSRRCRM8oCCMsCN0R(z.;R
RRSRRCRM8oCCMsCN0Rcz.;R
RRMRC8CRoMNCs0zCR.Rd;RS

RRRR-t-RCsMCNR0C0REC)RqvODCD#MRN8CR#D0CORoDFHVORF)sRq4vAnc_1_
1cSUz.RH:RVOR5EOFHCH_I8R0E=2RcRMoCC0sNCz
SO:E	RRHV58N8s8IH0>ERR24.RMoCC0sNCRR
RRRRRkRRORD	:sRbF#OC#p5BiR2
RRRRRRRRLHCoMR
RRRRRRRRRH5VRB'piCMPC0MRN8pRBiRR='24'RC0EMR
RRRRRRRRRR_RsNs88_osC58N8s8IH04E-RI8FMR0F4R.2<)=Rq)7758N8s8IH04E-RI8FMR0F4;.2
RRRRRRRRCRRMH8RVR;
RRRRRCRRMb8RsCFO#k#RO;D	
RSRCRM8oCCMsCN0REzO	R;
RSRRzR.g:FRVsRRHH5MR80CbEk_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0SC
-Q-RVNR58I8sHE80R4>R.M2RCRC80OFRs0CNCsRIHR0CCLMNDNCRMF8Rkk0b0MRCNCLDRD#CCRO0DHFoOR
RRRRRRzRSd:jRRRHV58N8s8IH0>ERR24.RMoCC0sNC-
S-HRVGFRVsNROD4DRd(UU,CR#D0CORRFV0#sH0CN0R0MFRHLCMsoRC#oH0CCs8R
RRRRRRRRRRRRRRFRskC0_M25HRR<='R4'IMECR_5sNs88_osC58N8s8IH04E-RI8FMR0F4R.2=2RHR#CDCjR''S;
SISSF_k0CHM52=R<R''4RCIEMIR5Ns8_CNo58I8sHE80-84RF0IMF.R42RR-HC2RDR#C';j'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RWRCIEMIR5Ns8_CNo58I8sHE80-84RF0IMF.R42RR=HC2RDR#C';j'
RRRRRRRRMSC8CRoMNCs0zCRd
j;SR--Q5VRNs88I0H8E=R<R24.RRMFI0sHCMRCNCLDRRFsFbk0kC0RMDNLCCR#D0CORoDFHMORCCC88S
RRRRRS4zdRH:RVNR58I8sHE80RR<=4R.2oCCMsCN0
SSSSksF0M_C5RH2<'=R4
';SSSSI0Fk_5CMH<2R=4R''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=W
 ;RRRRRRRRS8CMRMoCC0sNCdRz4S;
-t-RCsMCNR0C0REC)RqvODCD#MRN8sR0H0-#N#0C
RRRRRRRRdSz.RR:VRFs[MRHRH5I8_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
RRRRRRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVAv)q_gcjn7XcRD:RNDLCRRH#";W"
RRRRRRRRRRRRRRRRoLCHRM
RRRRRRRRRSRRAv)q_gcjn7XcR):Rq4vAnc_1_
1cSRRRRRRRRRRRRsbF0NRlb7R5Q=qR>MRH_osC5[c*+8dRF0IMF*Rc[R2,q)77q>R=RIDF_8IN84s54FR8IFM0R,j2RA7QRR=>"jjjjR",q)77A>R=RIDF_8sN84s54FR8IFM0R,j2
SSSSq hRR=>',4'R)11q>R=R''j, RWq>R=R0Is_5CMHR2,BqpiRR=>B,piRA hRR=>',4'R)11A>R=R''j, RWA>R=R''j,pRBi=AR>pRBiS,
S7SSmdq52>R=RkIF0k_L#Hc5,*Rc[2+d,SR
S7SSm.q52>R=RkIF0k_L#Hc5,[c*+,.2RS
SSmS7q254RR=>I0Fk_#Lkc,5Hc+*[4R2,
SSSSq7m5Rj2=I>RF_k0Lck#5RH,c2*[,S
SSmS7A25dRR=>s0Fk_#Lkc,5HR[c*+,d2RS
SSmS7A25.RR=>s0Fk_#Lkc,5Hc+*[.R2,
SSSSA7m5R42=s>RF_k0Lck#5cH,*4[+2
,RSSSS75mAj=2R>FRskL0_k5#cHc,R*2[2;S
SSFSsks0_Cco5*R[2<s=RF_k0Lck#5cH,*R[2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRsks0_Cco5*4[+2=R<RksF0k_L#Hc5,[c*+R42IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRsks0_Cco5*.[+2=R<RksF0k_L#Hc5,[c*+R.2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRsks0_Cco5*d[+2=R<RksF0k_L#Hc5,[c*+Rd2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRIks0_Cco5*R[2<I=RF_k0Lck#5cH,*R[2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRIks0_Cco5*4[+2=R<RkIF0k_L#Hc5,[c*+R42IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRIks0_Cco5*.[+2=R<RkIF0k_L#Hc5,[c*+R.2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRIks0_Cco5*d[+2=R<RkIF0k_L#Hc5,[c*+Rd2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R

RRRRRSRRCRM8oCCMsCN0R.zd;R
RRSRRCRM8oCCMsCN0Rgz.;R
RRMRC8CRoMNCs0zCR.
U;
RSRR-R-RMtCC0sNCER0CqR)vCRODRD#NRM8#CCDOD0RFOoHRsVFRv)qA_4n11g_gz
Sd:dRRRHV5FOEH_OCI0H8ERR=go2RCsMCN
0CSEzO	RR:H5VRNs88I0H8ERR>4R42oCCMsCN0
RRRRRRRRDkO	RR:bOsFC5##B2pi
RRRRRRRRCRLo
HMRRRRRRRRRVRHRp5BiP'CCRM0NRM8BRpi=4R''02RE
CMRRRRRRRRRRRRs8_N8ss_CNo58I8sHE80-84RF0IMF4R42=R<R7)q7N)58I8sHE80-84RF0IMF4R42R;
RRRRRRRRR8CMR;HV
RRRRRRRR8CMRFbsO#C#RDkO	S;
RMRC8CRoMNCs0zCRO;E	
RRRRdSzcRR:VRFsHMRHRC58b_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
-S-RRQV58N8s8IH0>ERR244RCMC8FR0RCOsNR0CI0sHCMRCNCLDR8NMR0FkbRk0CLMND#CRCODC0FRDo
HORRRRRRRRS6zdRH:RVNR58I8sHE80R4>R4o2RCsMCN
0CSR--VRHGVRFsODNDRU4dUR(,#CCDOF0RVsR0HN#00MCRFL0RCoHMRosCHC#0s
C8RRRRRRRRRRRRRRRRs0Fk_5CMH<2R=4R''ERIC5MRs8_N8ss_CNo58I8sHE80-84RF0IMF4R42RR=HC2RDR#C';j'
SSSSkIF0M_C5RH2<'=R4I'RERCM58IN_osC58N8s8IH04E-RI8FMR0F4R42=2RHR#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=WI RERCM58IN_osC58N8s8IH04E-RI8FMR0F4R42=2RHR#CDCjR''R;
RRRRRSRRCRM8oCCMsCN0R6zd;-
S-VRQR85N8HsI8R0E<4=R4M2RFsRIHR0CCLMNDFCRskRF00bkRNCMLRDC#CCDOD0RFOoHRCMC8
C8RRSRRzRSd:nRRRHV58N8s8IH0<ER=4R42CRoMNCs0SC
RRRRRRRRRRRRs0Fk_5CMH<2R=4R''S;
SISSF_k0CHM52=R<R''4;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R R;
RRRRRSRRCRM8oCCMsCN0Rnzd;-
S-CRtMNCs00CRE)CRqOvRC#DDR8NMRH0s-N#00
C#RRRRRRRRS(zdRV:RF[sRRRHM58IH0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CRRRRRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FAVR)_qv.UjcXRU7:NRDLRCDH"#RW
";RRRRRRRRRRRRRRRRLHCoMR
RRRRRRRRRRARS)_qv.UjcXRU7:qR)vnA4__1g1Rg
RRRRRRRRRRRRRRRRRsbF0NRlb7R5Q=qR>MRH_osC5[g*+8(RF0IMF*Rg[R2,q)77q>R=RIDF_8IN84s5jFR8IFM0R,j2RA7QRR=>"jjjjjjjjR",q)77A>R=RIDF_8sN84s5jFR8IFM0R,j2
SSSSq hRR=>',4'R)11q>R=R''j, RWq>R=R0Is_5CMHR2,BqpiRR=>B,piRA hRR=>',4'R)11A>R=R''j, RWA>R=R''j,pRBi=AR>pRBi
,RSSSS75mq(=2R>FRIkL0_k5#UH*,U[2+(,SR
S7SSmnq52>R=RkIF0k_L#HU5,[U*+,n2RS
SSmS7q256RR=>I0Fk_#LkU,5HU+*[6R2,
SSSSq7m5Rc2=I>RF_k0LUk#5UH,*c[+2
,RSSSS75mqd=2R>FRIkL0_k5#UH*,U[2+d,SR
S7SSm.q52>R=RkIF0k_L#HU5,[U*+,.2RS
SSmS7q254RR=>I0Fk_#LkU,5HU+*[4R2,
SSSSq7m5Rj2=I>RF_k0LUk#5UH,*,[2RS
SSmS7A25(RR=>s0Fk_#LkU,5HU+*[(R2,
SSSSA7m5Rn2=s>RF_k0LUk#5UH,*n[+2
,RSSSS75mA6=2R>FRskL0_k5#UH*,U[2+6,SR
S7SSmcA52>R=RksF0k_L#HU5,[U*+,c2RS
SSmS7A25dRR=>s0Fk_#LkU,5HU+*[dR2,
SSSSA7m5R.2=s>RF_k0LUk#5UH,*.[+2
,RSSSS75mA4=2R>FRskL0_k5#UH*,U[2+4,SR
S7SSmjA52>R=RksF0k_L#HU5,[U*2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRR7qQu5Rj2=H>RMC_so*5g[2+U,QR7u=AR>jR""R,
RRRRRRRRRRRRRRRRRRRRRRRRR7RRm5uqj=2R>bRIN0sH$k_L#HU5,,[2Ru7mA25jRR=>ssbNH_0$LUk#5[H,2
2;RRRRRRRRRRRRRRRRs0Fk_osC5[g*2=R<RksF0k_L#HU5,[U*2ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRs0Fk_osC5[g*+R42<s=RF_k0LUk#5UH,*4[+2ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRs0Fk_osC5[g*+R.2<s=RF_k0LUk#5UH,*.[+2ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRs0Fk_osC5[g*+Rd2<s=RF_k0LUk#5UH,*d[+2ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRs0Fk_osC5[g*+Rc2<s=RF_k0LUk#5UH,*c[+2ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRs0Fk_osC5[g*+R62<s=RF_k0LUk#5UH,*6[+2ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRs0Fk_osC5[g*+Rn2<s=RF_k0LUk#5UH,*n[+2ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRs0Fk_osC5[g*+R(2<s=RF_k0LUk#5UH,*([+2ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRs0Fk_osC5[g*+RU2<s=RbHNs0L$_k5#UH2,[RCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRIRRF_k0s5Cog2*[RR<=I0Fk_#LkU,5HU2*[RCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRIRRF_k0s5Cog+*[4<2R=FRIkL0_k5#UH*,U[2+4RCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRIRRF_k0s5Cog+*[.<2R=FRIkL0_k5#UH*,U[2+.RCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRIRRF_k0s5Cog+*[d<2R=FRIkL0_k5#UH*,U[2+dRCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRIRRF_k0s5Cog+*[c<2R=FRIkL0_k5#UH*,U[2+cRCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRIRRF_k0s5Cog+*[6<2R=FRIkL0_k5#UH*,U[2+6RCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRIRRF_k0s5Cog+*[n<2R=FRIkL0_k5#UH*,U[2+nRCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRIRRF_k0s5Cog+*[(<2R=FRIkL0_k5#UH*,U[2+(RCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRIRRF_k0s5Cog+*[U<2R=bRIN0sH$k_L#HU5,R[2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRCRSMo8RCsMCNR0Cz;d(
RRRRCRSMo8RCsMCNR0Cz;dc
RRRR8CMRMoCC0sNCdRzd
;
SRRRRR--tCCMsCN0RC0ERv)qRDOCDN#RM#8RCODC0FRDoRHOVRFs)Aqv41n_41U_4SU
zRdU:VRHRE5OFCHO_8IH0=ERR24URMoCC0sNCz
SORE	:VRHR85N8HsI8R0E>jR42CRoMNCs0RC
RRRRRkRRORD	:sRbF#OC#p5BiR2
RRRRRRRRLHCoMR
RRRRRRRRRH5VRB'piCMPC0MRN8pRBiRR='24'RC0EMR
RRRRRRRRRR_RsNs88_osC58N8s8IH04E-RI8FMR0F4Rj2<)=Rq)7758N8s8IH04E-RI8FMR0F4;j2
RRRRRRRRCRRMH8RVR;
RRRRRCRRMb8RsCFO#k#RO;D	
RSRR8CMRMoCC0sNCORzE
	;RRRRSgzdRV:RFHsRRRHM5b8C0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CSR--Q5VRNs88I0H8ERR>4Rj2M8CCRR0FONsC0ICRsCH0RNCMLRDCNRM8Fbk0kC0RMDNLCCR#D0CORoDFHRO
RRRRRSRRzRcj:VRHR85N8HsI8R0E>jR42CRoMNCs0SC
-V-RHVGRFOsRNRDD4UdU(#,RCODC0VRFRH0s#00NCFRM0CRLHRMosHCo#s0CCR8
RRRRRRRRRRRRRsRRF_k0CHM52=R<R''4RCIEMsR5_8N8sC_so85N8HsI8-0E4FR8IFM0R24jRH=R2DRC#'CRj
';SSSSI0Fk_5CMH<2R=4R''ERIC5MRI_N8s5CoNs88I0H8ER-48MFI04FRj=2RR2HRR#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=WI RERCM58IN_osC58N8s8IH04E-RI8FMR0F4Rj2=2RHR#CDCjR''R;
RRRRRSRRCRM8oCCMsCN0Rjzc;-
S-VRQR85N8HsI8R0E<4=RjM2RFsRIHR0CCLMNDFCRskRF00bkRNCMLRDC#CCDOD0RFOoHRCMC8
C8RRSRRzRSc:4RRRHV58N8s8IH0<ER=jR42CRoMNCs0SC
RRRRRRRRRRRRs0Fk_5CMH<2R=4R''S;
SISSF_k0CHM52=R<R''4;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R R;
RRRRRSRRCRM8oCCMsCN0R4zc;-
S-CRtMNCs00CRE)CRqOvRC#DDR8NMRH0s-N#00
C#RRRRRRRRS.zcRV:RF[sRRRHM58IH0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CRRRRRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FAVR)_qv4cj.X74nRD:RNDLCRRH#";W"
RRRRRRRRRRRRRRRRoLCHRM
RRRRRRRRRSRRAv)q_.4jcnX47RR:)Aqv41n_41U_4RU
RRRRRRRRRRRRRRRRRsbF0NRlb7R5Q=qR>MRH_osC5*4U[6+4RI8FMR0F4[U*2q,R7q7)RR=>D_FII8N8sR5g8MFI0jFR27,RQ=AR>jR"jjjjjjjjjjjjj"jj,7Rq7R)A=D>RFsI_Ns8858gRF0IMF2Rj,S
SShS q>R=R''4,1R1)=qR>jR''W,R =qR>sRI0M_C5,H2RiBpq>R=RiBp,hR A>R=R''4,1R1)=AR>jR''W,R =AR>jR''B,RpRiA=B>RpRi,
SSSSq7m5246RR=>I0Fk_#Lk4Hn5,*4n[6+42
,RSSSS75mq4Rc2=I>RF_k0L4k#n,5H4[n*+24c,SR
S7SSm4q5d=2R>FRIkL0_kn#454H,n+*[4,d2RS
SSmS7q.542>R=RkIF0k_L#54nHn,4*4[+.R2,
SSSSq7m5244RR=>I0Fk_#Lk4Hn5,*4n[4+42
,RSSSS75mq4Rj2=I>RF_k0L4k#n,5H4[n*+24j,SR
S7SSmgq52>R=RkIF0k_L#54nHn,4*g[+2
,RSSSS75mqU=2R>FRIkL0_kn#454H,n+*[UR2,
SSSSq7m5R(2=I>RF_k0L4k#n,5H4[n*+,(2RS
SSmS7q25nRR=>I0Fk_#Lk4Hn5,*4n[2+n,SR
S7SSm6q52>R=RkIF0k_L#54nHn,4*6[+2
,RSSSS75mqc=2R>FRIkL0_kn#454H,n+*[cR2,
SSSSq7m5Rd2=I>RF_k0L4k#n,5H4[n*+,d2RS
SSmS7q25.RR=>I0Fk_#Lk4Hn5,*4n[2+.,SR
S7SSm4q52>R=RkIF0k_L#54nHn,4*4[+2
,RSSSS75mqj=2R>FRIkL0_kn#454H,n2*[,SR
S7SSm4A56=2R>FRskL0_kn#454H,n+*[4,62RS
SSmS7Ac542>R=RksF0k_L#54nHn,4*4[+cR2,
SSSSA7m524dRR=>s0Fk_#Lk4Hn5,*4n[d+42
,RSSSS75mA4R.2=s>RF_k0L4k#n,5H4[n*+24.,SR
S7SSm4A54=2R>FRskL0_kn#454H,n+*[4,42RS
SSmS7Aj542>R=RksF0k_L#54nHn,4*4[+jR2,
SSSSA7m5Rg2=s>RF_k0L4k#n,5H4[n*+,g2RS
SSmS7A25URR=>s0Fk_#Lk4Hn5,*4n[2+U,SR
S7SSm(A52>R=RksF0k_L#54nHn,4*([+2
,RSSSS75mAn=2R>FRskL0_kn#454H,n+*[nR2,
SSSSA7m5R62=s>RF_k0L4k#n,5H4[n*+,62RS
SSmS7A25cRR=>s0Fk_#Lk4Hn5,*4n[2+c,SR
S7SSmdA52>R=RksF0k_L#54nHn,4*d[+2
,RSSSS75mA.=2R>FRskL0_kn#454H,n+*[.R2,
SSSSA7m5R42=s>RF_k0L4k#n,5H4[n*+,42RS
SSmS7A25jRR=>s0Fk_#Lk4Hn5,*4n[R2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRu7Qq>R=R_HMs5Co4[U*+R4(8MFI04FRU+*[4,n2Ru7QA>R=Rj"j"R,
RRRRRRRRRRRRRRRRRRRRRRRRR7RRm5uq4=2R>bRIN0sH$k_L#54nH*,.[2+4,mR7ujq52>R=RNIbs$H0_#Lk4Hn5,[.*2R,
RRRRRRRRRRRRRRRRRRRRRRRRR7RRm5uA4=2R>bRsN0sH$k_L#54nH*,.[2+4,mR7ujA52>R=RNsbs$H0_#Lk4Hn5,[.*2
2;RRRRRRRRRRRRRRRRs0Fk_osC5*4U[<2R=FRskL0_kn#454H,n2*[RCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRsRRF_k0s5Co4[U*+R42<s=RF_k0L4k#n,5H4[n*+R42IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRsks0_C4o5U+*[.<2R=FRskL0_kn#454H,n+*[.I2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRksF0C_soU54*d[+2=R<RksF0k_L#54nHn,4*d[+2ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRs0Fk_osC5*4U[2+cRR<=s0Fk_#Lk4Hn5,*4n[2+cRCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRsRRF_k0s5Co4[U*+R62<s=RF_k0L4k#n,5H4[n*+R62IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRsks0_C4o5U+*[n<2R=FRskL0_kn#454H,n+*[nI2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRksF0C_soU54*([+2=R<RksF0k_L#54nHn,4*([+2ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRs0Fk_osC5*4U[2+URR<=s0Fk_#Lk4Hn5,*4n[2+URCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRsRRF_k0s5Co4[U*+Rg2<s=RF_k0L4k#n,5H4[n*+Rg2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRsks0_C4o5U+*[4Rj2<s=RF_k0L4k#n,5H4[n*+24jRCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRsRRF_k0s5Co4[U*+244RR<=s0Fk_#Lk4Hn5,*4n[4+42ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRs0Fk_osC5*4U[.+42=R<RksF0k_L#54nHn,4*4[+.I2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRksF0C_soU54*4[+d<2R=FRskL0_kn#454H,n+*[4Rd2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRsks0_C4o5U+*[4Rc2<s=RF_k0L4k#n,5H4[n*+24cRCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRsRRF_k0s5Co4[U*+246RR<=s0Fk_#Lk4Hn5,*4n[6+42ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRs0Fk_osC5*4U[n+42=R<RNsbs$H0_#Lk4Hn5,[.*2ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRs0Fk_osC5*4U[(+42=R<RNsbs$H0_#Lk4Hn5,[.*+R42IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R

RRRRRRRRRRRRRIRRF_k0s5Co4[U*2=R<RkIF0k_L#54nHn,4*R[2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRIks0_C4o5U+*[4<2R=FRIkL0_kn#454H,n+*[4I2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRkIF0C_soU54*.[+2=R<RkIF0k_L#54nHn,4*.[+2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRI0Fk_osC5*4U[2+dRR<=I0Fk_#Lk4Hn5,*4n[2+dRCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRIRRF_k0s5Co4[U*+Rc2<I=RF_k0L4k#n,5H4[n*+Rc2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRIks0_C4o5U+*[6<2R=FRIkL0_kn#454H,n+*[6I2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRkIF0C_soU54*n[+2=R<RkIF0k_L#54nHn,4*n[+2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRI0Fk_osC5*4U[2+(RR<=I0Fk_#Lk4Hn5,*4n[2+(RCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRIRRF_k0s5Co4[U*+RU2<I=RF_k0L4k#n,5H4[n*+RU2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRIks0_C4o5U+*[g<2R=FRIkL0_kn#454H,n+*[gI2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRkIF0C_soU54*4[+j<2R=FRIkL0_kn#454H,n+*[4Rj2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRIks0_C4o5U+*[4R42<I=RF_k0L4k#n,5H4[n*+244RCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRIRRF_k0s5Co4[U*+24.RR<=I0Fk_#Lk4Hn5,*4n[.+42ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRI0Fk_osC5*4U[d+42=R<RkIF0k_L#54nHn,4*4[+dI2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRkIF0C_soU54*4[+c<2R=FRIkL0_kn#454H,n+*[4Rc2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRIks0_C4o5U+*[4R62<I=RF_k0L4k#n,5H4[n*+246RCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRIRRF_k0s5Co4[U*+24nRR<=IsbNH_0$L4k#n,5H.2*[RCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRIRRF_k0s5Co4[U*+24(RR<=IsbNH_0$L4k#n,5H.+*[4I2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
R
RRRRRRCRSMo8RCsMCNR0Cz;c.
RRRRCRSMo8RCsMCNR0Cz;dg
RRRR8CMRMoCC0sNCdRzU
;
SRRRRR--tCCMsCN0RC0ERv)qRDOCDN#RM#8RCODC0FRDoRHOVRFs)Aqv41n_d1n_dSn
zNdURH:RVOR5EOFHCH_I8R0E=nRd2CRoMNCs0SC
z	OERH:RVNR58I8sHE80Rg>R2CRoMNCs0SC
RRRRk	ODRb:RsCFO#B#5p
i2SLSRCMoH
RSSRRHV5iBp'CCPMN0RMB8Rp=iRR''42ER0CSM
SRRRRNs_8_8ss5CoNs88I0H8ER-48MFI0gFR2=R<R7)q7N)58I8sHE80-84RF0IMF2Rg;S
SRMRC8VRH;S
SCRM8bOsFCR##k	OD;R
SRMRC8CRoMNCs0zCRO;E	
RSRRdRzg:NRRsVFRHHRM8R5CEb0_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNC-
S-VRQR85N8HsI8R0E>2RgRCMC8FR0RCOsNR0CI0sHCMRCNCLDR8NMR0FkbRk0CLMND#CRCODC0FRDo
HOSzSScRjN:VRHR85N8HsI8R0E>2RgRMoCC0sNC-
S-HRVGFRVsNROD4DRd(UU,CR#D0CORRFV0#sH0CN0R0MFRHLCMsoRC#oH0CCs8S
SSFSskC0_M25HRR<='R4'IMECR_5sNs88_osC58N8s8IH04E-RI8FMR0Fg=2RRRH2CCD#R''j;S
SSFSIkC0_M25HRR<='R4'IMECRN5I8C_so85N8HsI8-0E4FR8IFM0RRg2=RRH2DRC#'CRj
';SSSSI_s0CHM52=R<RRW IMECRN5I8C_so85N8HsI8-0E4FR8IFM0RRg2=2RHR#CDCjR''S;
SMSC8CRoMNCs0zCRc;jN
-S-RRQV58N8s8IH0<ER=2RgRRMFI0sHCMRCNCLDRRFsFbk0kC0RMDNLCCR#D0CORoDFHMORCCC88S
SS4zcNRR:H5VRNs88I0H8E=R<RRg2oCCMsCN0
SSSSksF0M_C5RH2<'=R4
';SSSSI0Fk_5CMH<2R=4R''S;
SISSsC0_M25HRR<=W
 ;SCSSMo8RCsMCNR0CzNc4;-
S-CRtMNCs00CRE)CRqOvRC#DDR8NMRH0s-N#00
C#SzSScR.N:FRVsRR[H5MRI0H8Ek_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0RC
RRRRRRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)RAq6v_4d.X.:7RRLDNCHDR#WR""R;
RRRRRRRRRRRRRLRRCMoH
SSSSqA)v4_6..Xd7RR:)Aqv41n_d1n_dRn
RRRRRRRRRRRRRRRRRbRRFRs0lRNb5q7QRR=>HsM_Cdo5n+*[d84RF0IMFnRd*,[2R7q7)=qR>FRDIN_I858sUFR8IFM0R,j2RA7QRR=>"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjR",q)77A>R=RIDF_8sN8Us5RI8FMR0Fj
2,SSSS Rhq='>R4R',1q1)RR=>',j'RqW RR=>I_s0CHM52B,RpRiq=B>RpRi, RhA='>R4R',1A1)RR=>',j'RAW RR=>',j'RiBpA>R=RiBp,S
SSmS7q45d2>R=RkIF0k_L#5d.H.,d*d[+4R2,
SSSSq7m52djRR=>I0Fk_#LkdH.5,*d.[j+d2S,
S7SSm.q5g=2R>FRIkL0_k.#d5dH,.+*[.,g2RS
SSmS7qU5.2>R=RkIF0k_L#5d.H.,d*.[+UR2,
SSSSq7m52.(RR=>I0Fk_#LkdH.5,*d.[(+.2S,
S7SSm.q5n=2R>FRIkL0_k.#d5dH,.+*[.,n2RS
SSmS7q65.2>R=RkIF0k_L#5d.H.,d*.[+6R2,
SSSSq7m52.cRR=>I0Fk_#LkdH.5,*d.[c+.2S,
S7SSm.q5d=2R>FRIkL0_k.#d5dH,.+*[.,d2RS
SSmS7q.5.2>R=RkIF0k_L#5d.H.,d*.[+.R2,
SSSSq7m52.4RR=>I0Fk_#LkdH.5,*d.[4+.2S,
S7SSm.q5j=2R>FRIkL0_k.#d5dH,.+*[.,j2RS
SSmS7qg542>R=RkIF0k_L#5d.H.,d*4[+gR2,
SSSSq7m524URR=>I0Fk_#LkdH.5,*d.[U+42S,
S7SSm4q5(=2R>FRIkL0_k.#d5dH,.+*[4,(2RS
SSmS7qn542>R=RkIF0k_L#5d.H.,d*4[+nR2,
SSSSq7m5246RR=>I0Fk_#LkdH.5,*d.[6+42S,
S7SSm4q5c=2R>FRIkL0_k.#d5dH,.+*[4,c2RS
SSmS7qd542>R=RkIF0k_L#5d.H.,d*4[+dR2,
SSSSq7m524.RR=>I0Fk_#LkdH.5,*d.[.+42S,
S7SSm4q54=2R>FRIkL0_k.#d5dH,.+*[4,42RS
SSmS7qj542>R=RkIF0k_L#5d.H.,d*4[+jR2,
SSSSq7m5Rg2=I>RF_k0Ldk#.,5Hd[.*+,g2
SSSSq7m5RU2=I>RF_k0Ldk#.,5Hd[.*+,U2RS
SSmS7q25(RR=>I0Fk_#LkdH.5,*d.[2+(,SR
S7SSmnq52>R=RkIF0k_L#5d.H.,d*n[+2S,
S7SSm6q52>R=RkIF0k_L#5d.H.,d*6[+2
,RSSSS75mqc=2R>FRIkL0_k.#d5dH,.+*[cR2,
SSSSq7m5Rd2=I>RF_k0Ldk#.,5Hd[.*+,d2
SSSSq7m5R.2=I>RF_k0Ldk#.,5Hd[.*+,.2RS
SSmS7q254RR=>I0Fk_#LkdH.5,*d.[2+4,SR
S7SSmjq52>R=RkIF0k_L#5d.H.,d*,[2
SSSSA7m52d4RR=>s0Fk_#LkdH.5,*d.[4+d2
,RSSSS75mAdRj2=s>RF_k0Ldk#.,5Hd[.*+2dj,S
SSmS7Ag5.2>R=RksF0k_L#5d.H.,d*.[+gR2,
SSSSA7m52.URR=>s0Fk_#LkdH.5,*d.[U+.2
,RSSSS75mA.R(2=s>RF_k0Ldk#.,5Hd[.*+2.(,S
SSmS7An5.2>R=RksF0k_L#5d.H.,d*.[+nR2,
SSSSA7m52.6RR=>s0Fk_#LkdH.5,*d.[6+.2
,RSSSS75mA.Rc2=s>RF_k0Ldk#.,5Hd[.*+2.c,S
SSmS7Ad5.2>R=RksF0k_L#5d.H.,d*.[+dR2,
SSSSA7m52..RR=>s0Fk_#LkdH.5,*d.[.+.2
,RSSSS75mA.R42=s>RF_k0Ldk#.,5Hd[.*+2.4,S
SSmS7Aj5.2>R=RksF0k_L#5d.H.,d*.[+jR2,
SSSSA7m524gRR=>s0Fk_#LkdH.5,*d.[g+42
,RSSSS75mA4RU2=s>RF_k0Ldk#.,5Hd[.*+24U,S
SSmS7A(542>R=RksF0k_L#5d.H.,d*4[+(R2,
SSSSA7m524nRR=>s0Fk_#LkdH.5,*d.[n+42
,RSSSS75mA4R62=s>RF_k0Ldk#.,5Hd[.*+246,S
SSmS7Ac542>R=RksF0k_L#5d.H.,d*4[+cR2,
SSSSA7m524dRR=>s0Fk_#LkdH.5,*d.[d+42
,RSSSS75mA4R.2=s>RF_k0Ldk#.,5Hd[.*+24.,S
SSmS7A4542>R=RksF0k_L#5d.H.,d*4[+4R2,
SSSSA7m524jRR=>s0Fk_#LkdH.5,*d.[j+42
,RSSSS75mAg=2R>FRskL0_k.#d5dH,.+*[g
2,SSSS75mAU=2R>FRskL0_k.#d5dH,.+*[UR2,
SSSSA7m5R(2=s>RF_k0Ldk#.,5Hd[.*+,(2RS
SSmS7A25nRR=>s0Fk_#LkdH.5,*d.[2+n,S
SSmS7A256RR=>s0Fk_#LkdH.5,*d.[2+6,SR
S7SSmcA52>R=RksF0k_L#5d.H.,d*c[+2
,RSSSS75mAd=2R>FRskL0_k.#d5dH,.+*[d
2,SSSS75mA.=2R>FRskL0_k.#d5dH,.+*[.R2,
SSSSA7m5R42=s>RF_k0Ldk#.,5Hd[.*+,42RS
SSmS7A25jRR=>s0Fk_#LkdH.5,*d.[
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRQR7u=qR>MRH_osC5*dn[6+dRI8FMR0Fd[n*+2d.,QR7u=AR>jR"j"jj,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR7qmu5Rd2=I>RbHNs0L$_k.#d5cH,*d[+27,Rm5uq.=2R>bRIN0sH$k_L#5d.H*,c[2+.,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR7qmu5R42=I>RbHNs0L$_k.#d5cH,*4[+27,Rm5uqj=2R>bRIN0sH$k_L#5d.H*,c[
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7udA52>R=RNsbs$H0_#LkdH.5,[c*+,d2Ru7mA25.RR=>ssbNH_0$Ldk#.,5Hc+*[.
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7u4A52>R=RNsbs$H0_#LkdH.5,[c*+,42Ru7mA25jRR=>ssbNH_0$Ldk#.,5Hc2*[2R;
RRRRRRRRRRRRRRRRRksF0C_son5d*R[2<s=RF_k0Ldk#.,5Hd[.*2ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRsks0_Cdo5n+*[4<2R=FRskL0_k.#d5dH,.+*[4I2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRsRRF_k0s5Cod[n*+R.2<s=RF_k0Ldk#.,5Hd[.*+R.2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRs0Fk_osC5*dn[2+dRR<=s0Fk_#LkdH.5,*d.[2+dRCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRksF0C_son5d*c[+2=R<RksF0k_L#5d.H.,d*c[+2ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRsks0_Cdo5n+*[6<2R=FRskL0_k.#d5dH,.+*[6I2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRsRRF_k0s5Cod[n*+Rn2<s=RF_k0Ldk#.,5Hd[.*+Rn2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRs0Fk_osC5*dn[2+(RR<=s0Fk_#LkdH.5,*d.[2+(RCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRksF0C_son5d*U[+2=R<RksF0k_L#5d.H.,d*U[+2ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRsks0_Cdo5n+*[g<2R=FRskL0_k.#d5dH,.+*[gI2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRsRRF_k0s5Cod[n*+24jRR<=s0Fk_#LkdH.5,*d.[j+42ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRsks0_Cdo5n+*[4R42<s=RF_k0Ldk#.,5Hd[.*+244RCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRksF0C_son5d*4[+.<2R=FRskL0_k.#d5dH,.+*[4R.2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRs0Fk_osC5*dn[d+42=R<RksF0k_L#5d.H.,d*4[+dI2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRsRRF_k0s5Cod[n*+24cRR<=s0Fk_#LkdH.5,*d.[c+42ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRsks0_Cdo5n+*[4R62<s=RF_k0Ldk#.,5Hd[.*+246RCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRksF0C_son5d*4[+n<2R=FRskL0_k.#d5dH,.+*[4Rn2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRs0Fk_osC5*dn[(+42=R<RksF0k_L#5d.H.,d*4[+(I2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRsRRF_k0s5Cod[n*+24URR<=s0Fk_#LkdH.5,*d.[U+42ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRsks0_Cdo5n+*[4Rg2<s=RF_k0Ldk#.,5Hd[.*+24gRCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRksF0C_son5d*.[+j<2R=FRskL0_k.#d5dH,.+*[.Rj2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRs0Fk_osC5*dn[4+.2=R<RksF0k_L#5d.H.,d*.[+4I2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRsRRF_k0s5Cod[n*+2..RR<=s0Fk_#LkdH.5,*d.[.+.2ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRsks0_Cdo5n+*[.Rd2<s=RF_k0Ldk#.,5Hd[.*+2.dRCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRksF0C_son5d*.[+c<2R=FRskL0_k.#d5dH,.+*[.Rc2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRs0Fk_osC5*dn[6+.2=R<RksF0k_L#5d.H.,d*.[+6I2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRsRRF_k0s5Cod[n*+2.nRR<=s0Fk_#LkdH.5,*d.[n+.2ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRsks0_Cdo5n+*[.R(2<s=RF_k0Ldk#.,5Hd[.*+2.(RCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRksF0C_son5d*.[+U<2R=FRskL0_k.#d5dH,.+*[.RU2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRs0Fk_osC5*dn[g+.2=R<RksF0k_L#5d.H.,d*.[+gI2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRsRRF_k0s5Cod[n*+2djRR<=s0Fk_#LkdH.5,*d.[j+d2ERIC5MRs0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRsks0_Cdo5n+*[dR42<s=RF_k0Ldk#.,5Hd[.*+2d4RCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRksF0C_son5d*d[+.<2R=bRsN0sH$k_L#5d.H*,c[I2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRsRRF_k0s5Cod[n*+2ddRR<=ssbNH_0$Ldk#.,5Hc+*[4I2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRsRRF_k0s5Cod[n*+2dcRR<=ssbNH_0$Ldk#.,5Hc+*[.I2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRsRRF_k0s5Cod[n*+2d6RR<=ssbNH_0$Ldk#.,5Hc+*[dI2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR
RRRRRRRRRRRRRRRRRRRFRIks0_Cdo5n2*[RR<=I0Fk_#LkdH.5,*d.[I2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRIRRF_k0s5Cod[n*+R42<I=RF_k0Ldk#.,5Hd[.*+R42IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRI0Fk_osC5*dn[2+.RR<=I0Fk_#LkdH.5,*d.[2+.RCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRkIF0C_son5d*d[+2=R<RkIF0k_L#5d.H.,d*d[+2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRIks0_Cdo5n+*[c<2R=FRIkL0_k.#d5dH,.+*[cI2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRIRRF_k0s5Cod[n*+R62<I=RF_k0Ldk#.,5Hd[.*+R62IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRI0Fk_osC5*dn[2+nRR<=I0Fk_#LkdH.5,*d.[2+nRCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRkIF0C_son5d*([+2=R<RkIF0k_L#5d.H.,d*([+2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRIks0_Cdo5n+*[U<2R=FRIkL0_k.#d5dH,.+*[UI2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRIRRF_k0s5Cod[n*+Rg2<I=RF_k0Ldk#.,5Hd[.*+Rg2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRI0Fk_osC5*dn[j+42=R<RkIF0k_L#5d.H.,d*4[+jI2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRIRRF_k0s5Cod[n*+244RR<=I0Fk_#LkdH.5,*d.[4+42ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRIks0_Cdo5n+*[4R.2<I=RF_k0Ldk#.,5Hd[.*+24.RCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRkIF0C_son5d*4[+d<2R=FRIkL0_k.#d5dH,.+*[4Rd2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRI0Fk_osC5*dn[c+42=R<RkIF0k_L#5d.H.,d*4[+cI2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRIRRF_k0s5Cod[n*+246RR<=I0Fk_#LkdH.5,*d.[6+42ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRIks0_Cdo5n+*[4Rn2<I=RF_k0Ldk#.,5Hd[.*+24nRCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRkIF0C_son5d*4[+(<2R=FRIkL0_k.#d5dH,.+*[4R(2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRI0Fk_osC5*dn[U+42=R<RkIF0k_L#5d.H.,d*4[+UI2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRIRRF_k0s5Cod[n*+24gRR<=I0Fk_#LkdH.5,*d.[g+42ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRIks0_Cdo5n+*[.Rj2<I=RF_k0Ldk#.,5Hd[.*+2.jRCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRkIF0C_son5d*.[+4<2R=FRIkL0_k.#d5dH,.+*[.R42IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRI0Fk_osC5*dn[.+.2=R<RkIF0k_L#5d.H.,d*.[+.I2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRIRRF_k0s5Cod[n*+2.dRR<=I0Fk_#LkdH.5,*d.[d+.2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRIks0_Cdo5n+*[.Rc2<I=RF_k0Ldk#.,5Hd[.*+2.cRCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRkIF0C_son5d*.[+6<2R=FRIkL0_k.#d5dH,.+*[.R62IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRI0Fk_osC5*dn[n+.2=R<RkIF0k_L#5d.H.,d*.[+nI2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRIRRF_k0s5Cod[n*+2.(RR<=I0Fk_#LkdH.5,*d.[(+.2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRIks0_Cdo5n+*[.RU2<I=RF_k0Ldk#.,5Hd[.*+2.URCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRkIF0C_son5d*.[+g<2R=FRIkL0_k.#d5dH,.+*[.Rg2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRI0Fk_osC5*dn[j+d2=R<RkIF0k_L#5d.H.,d*d[+jI2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRIRRF_k0s5Cod[n*+2d4RR<=I0Fk_#LkdH.5,*d.[4+d2ERIC5MRI0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRFRIks0_Cdo5n+*[dR.2<I=RbHNs0L$_k.#d5cH,*R[2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRI0Fk_osC5*dn[d+d2=R<RNIbs$H0_#LkdH.5,[c*+R42IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRI0Fk_osC5*dn[c+d2=R<RNIbs$H0_#LkdH.5,[c*+R.2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRI0Fk_osC5*dn[6+d2=R<RNIbs$H0_#LkdH.5,[c*+Rd2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;S

SMSC8CRoMNCs0zCRc;.N
CSSMo8RCsMCNR0CzNdg;C
SMo8RCsMCNR0CzNdU;R
RCRM8oCCMsCN0Rdzc;R

RczcRH:RVMR5Fs0RNs88_osC2CRoMNCs0-CR-CRoMNCs0#CRCODC0NRslR
RR-R-RRQVNs88I0H8ERR<6#RN#MHoR''jRR0Fk#MkCL8RH
0#RRRRzRjR:VRHR85N8HsI8R0E=2R4RMoCC0sNCR
RRRRRRFRDIN_s8_8s#=R<Rj"jj"jjRs&RNs8_C#o_5;j2
RRRRRRRRIDF_8IN8#s_RR<="jjjjRj"&NRI8C_so5_#j
2;RRRRCRM8oCCMsCN0R;zj
RRRRRz4RH:RVNR58I8sHE80R.=R2CRoMNCs0RC
RRRRRDRRFsI_Ns88_<#R=jR"j"jjRs&RNs8_C#o_584RF0IMF2Rj;R
RRRRRRFRDIN_I8_8s#=R<Rj"jjRj"&NRI8C_so5_#4FR8IFM0R;j2
RRRR8CMRMoCC0sNC4Rz;R
RR.RzRRR:H5VRNs88I0H8ERR=do2RCsMCN
0CRRRRRRRRD_FIs8N8sR_#<"=Rj"jjRs&RNs8_C#o_58.RF0IMF2Rj;R
RRRRRRFRDIN_I8_8s#=R<Rj"jj&"RR8IN_osC_.#5RI8FMR0Fj
2;RRRRCRM8oCCMsCN0R;z.
RRRRRzdRH:RVNR58I8sHE80Rc=R2CRoMNCs0RC
RRRRRDRRFsI_Ns88_<#R=jR"j&"RR8sN_osC_d#5RI8FMR0Fj
2;RRRRRRRRD_FII8N8sR_#<"=RjRj"&NRI8C_so5_#dFR8IFM0R;j2
RRRR8CMRMoCC0sNCdRz;z
ScRS:H5VRNs88I0H8ERR=6o2RCsMCN
0CSFSDIN_s8_8s#=R<R''jRs&RNs8_C#o_58cRF0IMF2Rj;S
SD_FII8N8sR_#<'=Rj&'RR8IN_osC_c#5RI8FMR0Fj
2;S8CMRMoCC0sNCcRz;R
RR6RzRRR:H5VRNs88I0H8ERR>6o2RCsMCN
0CRRRRRRRRD_FIs8N8sR_#<s=RNs8_C#o_586RF0IMF2Rj;R
RRRRRRFRDIN_I8_8s#=R<R8IN_osC_6#5RI8FMR0Fj
2;RRRRCRM8oCCMsCN0R;z6
R
RR-R-RRQV5M8H_osC2CRso0H#C7sRQkhR#oHMRiBp
RRRRRznRH:RV8R5HsM_CRo2oCCMsCN0
RRRRRRRRFbsO#C#Rp5Bi7,RQRh2LHCoMR
RRRRRRRRRRVRHRp5BiRR='R4'NRM8B'piCMPC002RE
CMRRRRRRRRRRRRRRRRHsM_C#o_RR<=7;Qh
RRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMRFbsO#C#;R
RRMRC8CRoMNCs0zCRnR;
RzRR(:RRRRHV50MFRM8H_osC2CRoMNCs0RC
RRRRRRRRRHRRMC_soR_#<7=RQ
h;RRRRCRM8oCCMsCN0R;z(
R
RR-R-RRQV5Fs8ks0_CRo2sHCo#s0CRz7ma#RkHRMomiBp
RRRRszURRR:H5VRsk8F0C_soo2RCsMCN
0CRRRRRRRRbOsFCR##5m)_B,piRksF0C_so2_#RoLCHRM
RRRRRRRRRHRRV)R5_pmBiRR='R4'NRM8)B_mpCi'P0CM2ER0CRM
RRRRRRRRRRRRR)RR_z7ma=R<RksF0C_so;_#
RRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMRFbsO#C#;R
RRMRC8CRoMNCs0zCRU
s;RRRRzRgsRH:RVMR5Fs0R80Fk_osC2CRoMNCs0RC
RRRRRRRRR)RR_z7ma=R<RksF0C_so;_#
RRRR8CMRMoCC0sNCgRzs
;
SIzURRR:H5VRIk8F0C_soo2RCsMCN
0CRRRRRRRRbOsFCR##5mW_B,piRkIF0C_so2_#RoLCHRM
RRRRRRRRRHRRVWR5_pmBiRR='R4'NRM8WB_mpCi'P0CM2ER0CRM
RRRRRRRRRRRRRWRR_z7ma=R<RkIF0C_so;_#
RRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMRFbsO#C#;R
RRMRC8CRoMNCs0zCRU
I;RRRRzRgIRH:RVMR5FI0R80Fk_osC2CRoMNCs0RC
RRRRRRRRRWRR_z7ma=R<RkIF0C_so;_#
RRRR8CMRMoCC0sNCgRzI
;
RRRR-Q-RVsR5Ns88_osC2CRso0H#CqsR7R7)kM#HopRBiR
RR4Rzj:RRRRHV58sN8ss_CRo2oCCMsCN0
RRRRRRRRFbsO#C#R_5)miBp,qR)727)RoLCHRM
RRRRRRRRRHRRV)R5_pmBiRR='R4'NRM8)B_mpCi'P0CM2ER0CRM
RRRRRRRRRRRRRsRRNs8_C#o_RR<=)7q7)85N8HsI8-0E4FR8IFM0R;j2
RRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMRFbsO#C#;R
RRMRC8CRoMNCs0zCR4
j;RRRRzR44:VRHRF5M0NRs8_8ss2CoRMoCC0sNCR
RRRRRRRRRRNRs8C_soR_#<)=Rq)77;R
RRMRC8CRoMNCs0zCR4
4;
RRRRR--Q5VRI8N8sC_sos2RC#oH0RCsq)77RHk#MBoRpRi
RzRR4R.R:VRHRN5I8_8ss2CoRMoCC0sNCR
RRRRRRsRbF#OC#BR5pRi,W7q7)L2RCMoH
RRRRRRRRRRRRRHV5iBpR'=R4N'RMB8RpCi'P0CM2ER0CRM
RRRRRRRRRRRRRIRRNs8_C#o_RR<=W7q7)85N8HsI8-0E4FR8IFM0R;j2
RRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMRFbsO#C#;R
RRMRC8CRoMNCs0zCR4
.;RRRRzR4d:VRHRF5M0NRI8_8ss2CoRMoCC0sNCR
RRRRRRRRRRNRI8C_soR_#<W=Rq)77;R
RRMRC8CRoMNCs0zCR4
d;RRRRRRRR
RRRRR--tCCMsCN0RC0ERv)qRDOCDN#RM#8RCODC0FRDo
HORRRRzR4c:FRVsRRHH5MRM_klODCD_Rnc-2R4RI8FMR0FjCRoMNCs0RC
R-RR-VRQR85N8HsI8R0E>2R6RCMC8FR0RCOsNR0CI0sHCMRCNCLDR8NMR0FkbRk0CLMND#CRCODC0FRDo
HORRRRRRRRzR46:VRHR85N8HsI8R0E>2RnRMoCC0sNCR
RRRRRRRRRRRRRRFRskC0_M5_#H<2R=4R''ERIC5MRs_N8s_Co#85N8HsI8-0E4FR8IFM0RRn2=2RHR#CDCjR''S;
SISSF_k0C#M_5RH2<'=R4I'RERCM58IN_osC_N#58I8sHE80-84RF0IMF2RnRH=R2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0C#M_5RH2<W=R ERIC5MRI_N8s_Co#85N8HsI8-0E4FR8IFM0RRn2=2RHR#CDCjR''R;
RRRRRCRRMo8RCsMCNR0Cz;46
RRRRR--Q5VRNs88I0H8E=R<RR62MIFRsCH0RNCMLRDCFFsRkk0b0MRCNCLDRD#CCRO0DHFoOCRMC88C
RRRRRRRRnz4RH:RVNR58I8sHE80RR<=no2RCsMCN
0CRRRRRRRRRRRRRRRRs0Fk__CM#25HRR<=';4'
SSSSkIF0M_C_H#52=R<R''4;R
RRRRRRRRRRRRRRsRI0M_C_H#52=R<R;W 
RRRRRRRR8CMRMoCC0sNC4RznR;
R-RR-CRtMNCs00CRE)CRqOvRC#DDR8NMRH0s-N#00
C#RRRRRRRRzR4(:FRVsRR[H5MRI0H8ERR-482RF0IMFRRjoCCMsCN0
RRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVzv)qn:cRRLDNCHDR#1R"7Ra"&MRH0CCosl'HN5oCI0H8E&2RR""7RH&RMo0CCHs'lCNo5nH*c&2RR""WRH&RMo0CCHs'lCNo5R[2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50E54H+2c*n,CR8b20E2RR&"RX"&MRH0CCosl'HN5oC[2+4;R
RRRRRRRRRRCRLo
HMRRRRRRRRRRRRzv)qn:cRRqX)vXnc4
7RRRRRRRRRRRRRRRRRb0FsRblNRR57=H>RMC_so5_#[R2,q=jR>FRDIN_I8_8s#25j,4RqRR=>D_FII8N8s5_#4R2,q=.R>FRDIN_I8_8s#25.,R
RRRRRRRRRRRRRRRRRRRRRRRRRq=dR>FRDIN_I8_8s#25d,cRqRR=>D_FII8N8s5_#cR2,q=6R>FRDIN_I8_8s#256,SR
SSSSS7RRuj)qRR=>D_FIs8N8s5_#jR2,7qu)4>R=RIDF_8sN8#s_5,42R)7uq=.R>FRDIN_s8_8s#25.,S
SSSSSRuR7)Rqd=D>RFsI_Ns88_d#527,Ruc)qRR=>D_FIs8N8s5_#cR2,7qu)6>R=RIDF_8sN8#s_5,62RS
SSSSSR RWRR=>I_s0C#M_5,H2RpWBi>R=RiBp,uR7m>R=RksF0k_L#c_n#,5H[R2,1Rum=I>RF_k0L_k#n5c#H2,[2R;
RRRRRRRRRRRRRsRRF_k0s_Co#25[RR<=s0Fk_#Lk_#nc5[H,2ERIC5MRs0Fk__CM#25HR'=R4R'2CCD#R''Z;S
SSFSIks0_C#o_5R[2<I=RF_k0L_k#n5c#H2,[RCIEMIR5F_k0C#M_5RH2=4R''C2RDR#C';Z'
RRRRRRRR8CMRMoCC0sNC4Rz(R;
RRRRCRM8oCCMsCN0Rcz4;RRRRRRRRRRRRR
RRRRR
RRRRR--tCCMsCN0RdNR.FRIs88RCRCb)RqvODCDRRHVNsbbFHbsNR0CRRRRRRRRRRRRRRR
RzRR4:URRRHV5lMk_DOCD._dR4=R2CRoMNCs0RC
R-RR-VRQR85N8HsI8R0E>2R(RCMC8FR0RCOsNR0CI0sHCMRCNCLDR8NMR0FkbRk0CLMND#CRCODC0FRDo
HORRRRRRRRzN4gRH:RVNR58I8sHE80Rn>R2CRoMNCs0RC
RRRRRRRRRRRRRsRRF_k0CdM_.=R<R''4RCIEM5R5s_N8s_Co#85N8HsI8-0E4FR8IFM0RRn2=kRMlC_ODnD_cN2RM58Rs_N8s_Co#256R'=Rj2'2R#CDCjR''S;
SISSF_k0CdM_.=R<R''4RCIEM5R5I_N8s_Co#85N8HsI8-0E4FR8IFM0RRn2=kRMlC_ODnD_cN2RM58RI_N8s_Co#256R'=Rj2'2R#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_M._dRR<=WI RERCM5N5I8C_so5_#Ns88I0H8ER-48MFI0nFR2RR=M_klODCD_2ncR8NMRN5I8C_so5_#6=2RR''j2C2RDR#C';j'
RRRRRRRR8CMRMoCC0sNC4Rzg
N;RRRRRRRRzL4gRH:RVNR58I8sHE80Rn=RR8NMRlMk_DOCDc_nRj=R2CRoMNCs0RC
RRRRRRRRRRRRRsRRF_k0CdM_.=R<R''4RCIEM5R5s_N8s_Co#256R'=Rj2'2R#CDCjR''S;
SISSF_k0CdM_.=R<R''4RCIEM5R5I_N8s_Co#256R'=Rj2'2R#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_M._dRR<=WI RERCM5N5I8C_so5_#6=2RR''j2C2RDR#C';j'
RRRRRRRR8CMRMoCC0sNC4RzgRL;R-RR-VRQR85N8HsI8R0E<6=R2FRMRHIs0CCRMDNLCsRFR0FkbRk0CLMND#CRCODC0FRDoRHOM8CCCR8
RRRRRzRR.:jRRRHV58N8s8IH0<ER=2R6RMoCC0sNCR
RRRRRRRRRRRRRRFRskC0_M._dRR<=';4'
SSSSkIF0M_C_Rd.<'=R4
';RRRRRRRRRRRRRRRRI_s0CdM_.=R<R;W 
RRRRRRRR8CMRMoCC0sNC.RzjR;
R-RR-CRtMNCs00CRE)CRqOvRCRDDNRM80-sH#00NCR
RRRRRR.Rz4RR:VRFs[MRHRH5I8R0E-2R4RI8FMR0FjCRoMNCs0RC
RRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)Rzq.vdRD:RNDLCRRH#"a17"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloMC5kOl_C_DDnnc*c&2RR""WRH&RMo0CCHs'lCNo5R[2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50EM_klODCD_*ncn+cRR,d.Rb8C02E2R"&RX&"RR0HMCsoC'NHlo[C5+;42
RRRRRRRRRRRRoLCHRM
RRRRRRRRRzRR)dqv.RR:Xv)qd4.X7RR
RRRRRRRRRRRRRbRRFRs0lRNb5=7R>MRH_osC_[#52q,Rj>R=RIDF_8IN8#s_5,j2RRq4=D>RFII_Ns88_4#52q,R.>R=RIDF_8IN8#s_5,.2
RRRRRRRRRRRRRRRRRRRRRRRRqRRd>R=RIDF_8IN8#s_5,d2RRqc=D>RFII_Ns88_c#52
,RSSSSSRSR7qu)j>R=RIDF_8sN8#s_5,j2R)7uq=4R>FRDIN_s8_8s#254,uR7)Rq.=D>RFsI_Ns88_.#52S,
SSSSS7RRud)qRR=>D_FIs8N8s5_#dR2,7qu)c>R=RIDF_8sN8#s_5,c2RS
SSSSSR RWRR=>I_s0CdM_.W,RBRpi=B>RpRi,7Rum=s>RF_k0L_k#d5.#M_klODCD_,d.[R2,1Rum=I>RF_k0L_k#d5.#M_klODCD_,d.[;22
RRRRRRRRRRRRRRRRksF0C_so5_#[<2R=FRskL0_kd#_.M#5kOl_C_DDd[.,2ERIC5MRs0Fk__CMd=.RR''42DRC#'CRZ
';SSSSI0Fk_osC_[#52=R<RkIF0k_L#._d#k5MlC_ODdD_.2,[RCIEMIR5F_k0CdM_.RR='24'R#CDCZR''R;
RRRRRRRRCRM8oCCMsCN0R4z.;R
RRCRRMo8RCsMCNR0Cz;4URRRRRRRRR
R
RRRR-t-RCsMCNR0CNnR4RsIF8CR8C)bRqOvRCRDDHNVRbFbsbNsH0RCRRRRRRRRRRRRRRR
RR.Rz.RR:H5VRM_klODCD_R4n=2R4RMoCC0sNCR
RR-R-RRQV58N8s8IH0>ERRR62M8CCRR0FONsC0ICRsCH0RNCMLRDCNRM8Fbk0kC0RMDNLCCR#D0CORoDFHRO
RRRRRzRR.RdN:VRHR85N8HsI8R0E>RRnNRM8M_klODCD_Rd.=2R4RMoCC0sNCR
RRRRRRRRRRRRRRFRskC0_Mn_4RR<='R4'IMECRs55Ns8_C#o_58N8s8IH04E-RI8FMR0Fn=2RRlMk_DOCDc_n2MRN8sR5Ns8_C#o_5R62=4R''N2RM58Rs_N8s_Co#25cR'=Rj2'2R#CDCjR''S;
SISSF_k0C4M_n=R<R''4RCIEM5R5I_N8s_Co#85N8HsI8-0E4FR8IFM0RRn2=kRMlC_ODnD_cN2RM58RI_N8s_Co#256R'=R4R'2NRM858IN_osC_c#52RR='2j'2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0C4M_n=R<RRW IMECRI55Ns8_C#o_58N8s8IH04E-RI8FMR0Fn=2RRlMk_DOCDc_n2MRN8IR5Ns8_C#o_5R62=4R''N2RM58RI_N8s_Co#25cR'=Rj2'2R#CDCjR''R;
RRRRRCRRMo8RCsMCNR0CzN.d;R
RRRRRR.Rzd:LRRRHV58N8s8IH0>ERRNnRMM8RkOl_C_DDd/.R=2R4RMoCC0sNCR
RRRRRRRRRRRRRRFRskC0_Mn_4RR<='R4'IMECRs55Ns8_C#o_58N8s8IH04E-RI8FMR0Fn=2RRlMk_DOCDc_n2MRN8sR5Ns8_C#o_5R62=jR''N2RM58Rs_N8s_Co#25cR'=Rj2'2R#CDCjR''S;
SISSF_k0C4M_n=R<R''4RCIEM5R5I_N8s_Co#85N8HsI8-0E4FR8IFM0RRn2=kRMlC_ODnD_cN2RM58RI_N8s_Co#256R'=RjR'2NRM858IN_osC_c#52RR='2j'2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0C4M_n=R<RRW IMECRI55Ns8_C#o_58N8s8IH04E-RI8FMR0Fn=2RRlMk_DOCDc_n2MRN8IR5Ns8_C#o_5R62=jR''N2RM58RI_N8s_Co#25cR'=Rj2'2R#CDCjR''R;
RRRRRCRRMo8RCsMCNR0CzL.d;R
RRRRRR.Rzd:ORRRHV58N8s8IH0=ERRNnRMM8RkOl_C_DDd=.RRR42oCCMsCN0
RRRRRRRRRRRRRRRRksF0M_C_R4n<'=R4I'RERCM5N5s8C_so5_#6=2RR''42MRN8sR5Ns8_C#o_5Rc2=jR''R22CCD#R''j;S
SSFSIkC0_Mn_4RR<='R4'IMECRI55Ns8_C#o_5R62=4R''N2RM58RI_N8s_Co#25cR'=Rj2'2R#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_Mn_4RR<=WI RERCM5N5I8C_so5_#6=2RR''42MRN8IR5Ns8_C#o_5Rc2=jR''R22CCD#R''j;R
RRRRRRMRC8CRoMNCs0zCR.;dO
RRRRRRRRdz.8RR:H5VRNs88I0H8ERR=6MRN8kRMlC_ODdD_.=R/RR42oCCMsCN0
RRRRRRRRRRRRRRRRksF0M_C_R4n<'=R4I'RERCM5N5s8C_so5_#Ns88I0H8ER-48MFI0cFR2RR=M_klODCD_2d.2DRC#'CRj
';SSSSI0Fk__CM4<nR=4R''ERIC5MR58IN_osC_N#58I8sHE80-84RF0IMF2RcRM=RkOl_C_DDd2.2R#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_Mn_4RR<=WI RERCM5N5I8C_so5_#Ns88I0H8ER-48MFI0cFR2RR=M_klODCD_2d.2DRC#'CRj
';RRRRRRRRCRM8oCCMsCN0Rdz.8R;RR-R-RRQV58N8s8IH0<ER=2R6RRMFI0sHCMRCNCLDRRFsFbk0kC0RMDNLCCR#D0CORoDFHMORCCC88R
RRRRRR.RzcRR:H5VRNs88I0H8E=R<RRc2oCCMsCN0
RRRRRRRRRRRRRRRRksF0M_C_R4n<'=R4
';SSSSI0Fk__CM4<nR=4R''R;
RRRRRRRRRRRRRIRRsC0_Mn_4RR<=W
 ;RRRRRRRRCRM8oCCMsCN0Rcz.;R
RR-R-RMtCC0sNCER0CqR)vCRODNDRM08Rs#H-0CN0
RRRRRRRR6z.RV:RF[sRRRHM58IH0-ERRR428MFI0jFRRMoCC0sNCR
RRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqz)vR4n:NRDLRCDH"#R1"7aRH&RMo0CCHs'lCNo58IH0RE2&7R""RR&HCM0o'CsHolNCk5MlC_ODnD_cc*nRM+RkOl_C_DDdd.*.&2RR""WRH&RMo0CCHs'lCNo5R[2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50EM_klODCD_*ncn+cRRlMk_DOCD._d*Rd.+nR4,CR8b20E2RR&"RX"&MRH0CCosl'HN5oC[2+4;R
RRRRRRRRRRCRLo
HMRRRRRRRRRRRRzv)q4:nRRv)q44nX7RR
RRRRRRRRRRRRRbRRFRs0lRNb5=7R>MRH_osC_[#52q,Rj>R=RIDF_8IN8#s_5,j2RRq4=D>RFII_Ns88_4#52q,R.>R=RIDF_8IN8#s_5,.2
RRRRRRRRRRRRRRRRRRRRRRRRqRRd>R=RIDF_8IN8#s_5,d2R)7uq=jR>FRDIN_s8_8s#25j,uR7)Rq4=D>RFsI_Ns88_4#527,Ru.)qRR=>D_FIs8N8s5_#.
2,SSSSSRSR7qu)d>R=RIDF_8sN8#s_5,d2RRW =I>RsC0_Mn_4,BRWp=iR>pRBi7,Ru=mR>FRskL0_k4#_nM#5kOl_C_DD4[n,21,Ru=mR>FRIkL0_k4#_nM#5kOl_C_DD4[n,2
2;RRRRRRRRRRRRRRRRs0Fk_osC_[#52=R<RksF0k_L#n_4#k5MlC_OD4D_n2,[RCIEMsR5F_k0C4M_nRR='24'R#CDCZR''S;
SISSF_k0s_Co#25[RR<=I0Fk_#Lk_#4n5lMk_DOCDn_4,R[2IMECRF5IkC0_Mn_4R'=R4R'2CCD#R''Z;R
RRRRRRMRC8CRoMNCs0zCR.
6;RRRRCRM8oCCMsCN0R.z.;RRRRR
RCRM8oCCMsCN0Rczc;M
C8sRNO0EHCkO0sMCRFI_s_COEO
	;

------
----NRp#H0RlCbDl0CMNF0HM#RHRV8CN0kD
----CR#D0CO_lsN
ONsECH0Os0kCCR#D0CO_lsNRRFV)_qv)_Wu)#RH
MVkOF0HMCRo0M_C8C_8b50E#CHxRH:RMo0CC;sRRb8C0:ERR0HMCsoC2CRs0MksR0HMCsoCR
H#PHNsNCLDRMlH_x#HCRR:HCM0oRCs:j=R;C
Lo
HMRHRlMH_#x:CR=CR8b;0E
HRRV#R5HRxC<CR8b20ERC0EMR
RRHRlMH_#x:CR=HR#x
C;RMRC8VRH;R
RskC0slMRH#M_H;xC
8CMR0oC_8CM_b8C0
E;O#FM00NMRlMk_DOCD:#RR0HMCsoCRR:=5C58bR0E-2R4/24n;RRRRRRRRRRRRR--yVRFRv)q44nX7CRODRD#M8CCC08
$RbCF_k0L_k#0C$bRRH#NNss$MR5kOl_C#DDRI8FMR0FjI,RHE80-84RF0IMF2RjRRFV#_08DHFoO#;
HNoMDFRskL0_k:#RR0Fk_#Lk_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$FsVR_k8F0HR5M0bkRR0F0-sH#00NC
#2#MHoNsDRF_k0C:MRR8#0_oDFHPO_CFO0sk5MlC_ODRD#8MFI0jFR2R;RRRRRRR--CLMNDRC#VRFs0-sH#00NC##
HNoMDFRIkC0_MRR:#_08DHFoOC_POs0F5lMk_DOCD8#RF0IMF2Rj;H
#oDMNRkIF0k_L#RR:F_k0L_k#0C$b;RRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RV_RI80FkRM5HbRk000FRs#H-0CN0##2
HNoMDsRI0M_CR#:R0D8_FOoH_OPC05FsM_klODCD#FR8IFM0R;j2RRRRRRRR-I-RsCH0RNCML#DCRsVFROCNEFRsIVRFRv)qRDOCD##
HNoMDMRH_osCR#:R0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2R;RRRRRRRRR-k-R#RC80sFRC#oH0RCs7RQh
o#HMRNDs0Fk_osCR#:R0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2R;RRRRRR-R-RCk#8FR0RosCHC#0s_R)7amz
o#HMRNDI0Fk_osCR#:R0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2R;RRRRRR-R-RCk#8FR0RosCHC#0s_RW7amz
o#HMRNDs_N8sRCo:0R#8F_Do_HOP0COFNs58I8sHE80-84RF0IMF2Rj;RRRR-R-RCk#8FR0RosCHC#0sqR)7
7)#MHoNIDRNs8_C:oRR8#0_oDFHPO_CFO0s85N8HsI8-0E4FR8IFM0R;j2RRRRRR--k8#CRR0FsHCo#s0CR7Wq7#)
HNoMDFRDIN_s8R8s:0R#8F_Do_HOP0COFds5RI8FMR0FjR2;RRRRRRRRRRRR-s-RNs88R0LH#MRHbRk00)FRqOvRC#DDRR5cL#H0RJsCkCHs8#2
HNoMDFRDIN_I8R8s:0R#8F_Do_HOP0COFds5RI8FMR0FjR2;RRRRRRRRRRRR-I-RNs88R0LH#MRHbRk00)FRqOvRC#DDRR5cL#H0RJsCkCHs8N2
0H0sLCk0Rs\3NFl_VCV#0:\RRs#0H;Mo
C
Lo
HM
RRRRR--QNVR8I8sHE80Rc<RR#N#HRoM'Rj'0kFRMCk#8HRL0R#
RzRR4:RRRRHV58N8s8IH0=ERRR42oCCMsCN0
RRRRRRRRIDF_8sN8<sR=jR"jRj"&NRs8C_so25j;R
RRRRRRFRDIN_I8R8s<"=Rj"jjRI&RNs8_Cjo52R;
RCRRMo8RCsMCNR0Cz
4;RRRRzR.R:VRHR85N8HsI8R0E=2R.RMoCC0sNCR
RRRRRRFRDIN_s8R8s<"=RjRj"&NRs8C_soR548MFI0jFR2R;
RRRRRDRRFII_Ns88RR<=""jjRI&RNs8_C4o5RI8FMR0Fj
2;RRRRCRM8oCCMsCN0R;z.
RRRRRzdRH:RVNR58I8sHE80Rd=R2CRoMNCs0RC
RRRRRDRRFsI_Ns88RR<='Rj'&NRs8C_soR5.8MFI0jFR2R;
RRRRRDRRFII_Ns88RR<='Rj'&NRI8C_soR5.8MFI0jFR2R;
RCRRMo8RCsMCNR0Cz
d;RRRRzRcR:VRHR85N8HsI8R0E>2RdRMoCC0sNCR
RRRRRRFRDIN_s8R8s<s=RNs8_Cdo5RI8FMR0Fj
2;RRRRRRRRD_FII8N8s=R<R8IN_osC58dRF0IMF2Rj;R
RRMRC8CRoMNCs0zCRc
;
RRRR-Q-RV8R5HsM_CRo2sHCo#s0CRh7QRHk#MBoRpRi
RzRR6:RRRRHV5M8H_osC2CRoMNCs0RC
RRRRRbRRsCFO#5#RB,piRh7Q2CRLo
HMRRRRRRRRRRRRH5VRBRpi=4R''MRN8pRBiP'CC2M0RC0EMR
RRRRRRRRRRRRRRMRH_osCRR<=7;Qh
RRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMRFbsO#C#;R
RRMRC8CRoMNCs0zCR6R;
RzRRn:RRRRHV50MFRM8H_osC2CRoMNCs0RC
RRRRRRRRRHRRMC_so=R<Rh7Q;R
RRMRC8CRoMNCs0zCRn
;
RRRR-Q-RVsR5F_k0s2CoRosCHC#0smR7zkaR#oHMRpmBiR
RR(Rzs:RRRRHV5Fs8ks0_CRo2oCCMsCN0
RRRRRRRRFbsO#C#R_5)miBp,FRsks0_CRo2LHCoMR
RRRRRRRRRRVRHR_5)miBpR'=R4N'RM)8R_pmBiP'CC2M0RC0EMR
RRRRRRRRRRRRRR_R)7amzRR<=s0Fk_osC;R
RRRRRRRRRRMRC8VRH;R
RRRRRRMRC8sRbF#OC#R;
RCRRMo8RCsMCNR0Cz;(s
RRRRszURRR:H5VRMRF0sk8F0C_soo2RCsMCN
0CRRRRRRRRRRRR)m_7z<aR=FRsks0_C
o;RRRRCRM8oCCMsCN0RszU;R

R-RR-VRQRF5sks0_CRo2sHCo#s0CRz7ma#RkHRMomiBp
RRRRIz(RRR:H5VRIk8F0C_soo2RCsMCN
0CRRRRRRRRbOsFCR##5mW_B,piRkIF0C_soL2RCMoH
RRRRRRRRRRRRRHV5mW_BRpi=4R''MRN8_RWmiBp'CCPMR020MEC
RRRRRRRRRRRRRRRR7W_mRza<I=RF_k0s;Co
RRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMRFbsO#C#;R
RRMRC8CRoMNCs0zCR(
I;RRRRzRUIRH:RVMR5FI0R80Fk_osC2CRoMNCs0RC
RRRRRRRRRWRR_z7ma=R<RkIF0C_soR;
RCRRMo8RCsMCNR0Cz;UI
R
RR-R-RRQV58sN8ss_CRo2sHCo#s0CR7)q7k)R#oHMRpmBiR
RRgRzRRR:H5VRs8N8sC_soo2RCsMCN
0CRRRRRRRRbOsFCR##5m)_B,piR7)q7R)2LHCoMR
RRRRRRRRRRVRHR_5)miBpR'=R4N'RM)8R_pmBiP'CC2M0RC0EMR
RRRRRRRRRRRRRRNRs8C_so=R<R7)q7N)58I8sHE80-84RF0IMF2Rj;R
RRRRRRRRRRMRC8VRH;R
RRRRRRMRC8sRbF#OC#R;
RCRRMo8RCsMCNR0Cz
g;RRRRzR4j:VRHRF5M0NRs8_8ss2CoRMoCC0sNCR
RRRRRRRRRRNRs8C_so=R<R7)q7
);RRRRCRM8oCCMsCN0Rjz4;R
RRRRRRRR
R-RR-VRQRN5I8_8ss2CoRosCHC#0sqRW7R7)kM#HopRBiR
RR4Rz6:RRRRHV58IN8ss_CRo2oCCMsCN0
RRRRRRRRFbsO#C#Rp5BiW,Rq)772CRLo
HMRRRRRRRRRRRRH5VRBRpi=4R''MRN8pRBiP'CC2M0RC0EMR
RRRRRRRRRRRRRRNRI8C_so=R<R7Wq7N)58I8sHE80-84RF0IMF2Rj;R
RRRRRRRRRRMRC8VRH;R
RRRRRRMRC8sRbF#OC#R;
RCRRMo8RCsMCNR0Cz;46
RRRRnz4RH:RVMR5FI0RNs88_osC2CRoMNCs0RC
RRRRRRRRRIRRNs8_C<oR=qRW7;7)
RRRR8CMRMoCC0sNC4Rzn
;
RRRR-t-RCsMCNR0C0REC)RqvODCD#MRN8CR#D0CORoDFHRO
RzRR4:4RRsVFRHHRMkRMlC_ODRD#8MFI0jFRRMoCC0sNCR
RRRRRR-R-RRQV58N8s8IH0>ERRRc2M8CCRR0FONsC0ICRsCH0RNCMLRDCNRM8Fbk0kC0RMDNLCCR#D0CORoDFHRO
RRRRRzRR4:.RRRHV58N8s8IH0>ERRRc2oCCMsCN0
RRRRRRRRRRRRRRRRksF0M_C5RH2<'=R4I'RERCM58sN_osC58N8s8IH04E-RI8FMR0Fc=2RRRH2CCD#R''j;R
RRRRRRRRRRRRRRFRIkC0_M25HRR<='R4'IMECRN5I8C_so85N8HsI8-0E4FR8IFM0RRc2=2RHR#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=WI RERCM58IN_osC58N8s8IH04E-RI8FMR0Fc=2RRRH2CCD#R''j;R
RRRRRRMRC8CRoMNCs0zCR4
.;RRRRRRRR-Q-RVNR58I8sHE80RR<=cM2RFsRIHR0CCLMNDFCRskRF00bkRNCMLRDC#CCDOD0RFOoHRCMC8
C8RRRRRRRRzR4d:VRHR85N8HsI8R0E<c=R2CRoMNCs0RC
RRRRRRRRRRRRRsRRF_k0CHM52=R<R''4;R
RRRRRRRRRRRRRRFRIkC0_M25HRR<=';4'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RW;R
RRRRRRRRRRMRC8CRoMNCs0zCR4
d;RRRR-t-RMNCs00CRE)CRqOvRC#DDR8NMRH0s-N#00
C#RRRRRRRRzR4c:FRVsRR[H5MRI0H8ERR-482RF0IMFRRjoCCMsCN0
RRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVzv)qRD:RNDLCRRH#"a17"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloHC5*24nR"&RW&"RR0HMCsoC'NHlo[C52RR&"R "&MRH0CCosl'HN5oCo_C0C_M880CbEH55+*424Rn,80CbER22&XR""RR&HCM0o'CsHolNC+5[4
2;RRRRRRRRRRRRLHCoMR
RRRRRRRRRR)RzqRv:)4qvn7X4RR
RRRRRRRRRRRRRRFRbsl0RN5bR7>R=R_HMs5Co[R2,q=jR>FRDIN_I858sjR2,q=4R>FRDIN_I858s4R2,q=.R>FRDIN_I858s.
2,RRRRRRRRRRRRRRRRRRRRRRRRRdRqRR=>D_FII8N8s25d,uR7)Rqj=D>RFsI_Ns885,j2R)7uq=4R>FRDIN_s858s4R2,
RRRRRRRRRRRRRRRRRRRRRRRR7RRu.)qRR=>D_FIs8N8s25.,uR7)Rqd=D>RFsI_Ns885,d2RRW =I>RsC0_M25H,RR
RRRRRRRRRRRRRRRRRRRRRRRRRpWBi>R=RiBp,uR7m>R=RksF0k_L#,5H[R2,1Rum=I>RF_k0L5k#H2,[2R;
RRRRRRRRRsRRF_k0s5Co[<2R=FRskL0_kH#5,R[2IMECRF5skC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRFRIks0_C[o52=R<RkIF0k_L#,5H[I2RERCM5kIF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRR8CMRMoCC0sNC4RzcR;
RRRRRCRRMo8RCsMCNR0Cz;44
RRRRRRRRRRRRRRRRRRRRRRRRRRRRCR
MN8RsHOE00COkRsC#CCDOs0_N
l;
