--
@ER--B$FbsEHo0OR52gR4g-cRRj.jd$R1MHbDO$H0ROQM
R--fN]C8:CsR#//$DMbH0OH$N/lb0DN.Uj4J4.b/blNb#Cs/0N0/LDH/MoC_OFsN/6o#Dlk0E3P8Ry4f-
-
-

-*R**************************************************************R*R---
-HR1o8MCRDvk0DHbH
Cs-a-RNCso0RR:p0N0HROCmNsOR-6
--
-R3R4RoDFH-ORRsRNsRN$l0kDHHbDCIsRHR0EbCHbL#kVRM5HR#ONCVRFRbbHCMDHH2Mo
R--
R--RR.3LODF	RR-kM#HosRmO6NRRFADOv	RkHD0bCDHsvR5z4paUUX42-
-
R--RbBF$osHE50RO.2Rj,jjRj.j4$R1MHbDO$H0,MRQO-3
-qRRDsDRH0oE#CRs#PCsC
83---
-*R**************************************************************R*R-
-
-*-R*************************************************************R**R
---#-RCODC0MHFR0#CRV8CH0MHH3FMR-R
-sRNOHED#=0RRoDFHLORD	FO_Dlk0-
-R****************************************************************-RR--

-*R**************************************************************R*R---
-HRwsu#0skF8O50#qA,R,ARq2-
-
R--W0H8E-qRR8IH0FERVRRqHkMb0-
-R8WH0REA-HRI8R0EFAVRRbHMk-0
--R
-ARqRL-RHN0IHR#CqRh7FNVRDHDRM0bk#-
-R-
-R****************************************************************-RR-D

HNLssH$RC;CCR#
kCCRHC#C30D8_FOoH_n44cD3ND
;
DsHLNRs$FNsOdk;
#FCRsdON3OFsNlOFbD3ND
;
DsHLNRs$#b$MD$HV;#
kC$R#MHbDVN$30H0sLCk0#D3ND
;
CHM00w$RH0s#u8sFk#O0R
H#RoRRCsMCH
O5RRRRRHRI8q0ERH:RMo0CC
s;RRRRRHRI8A0ERH:RMo0CCRs
R;R2
RRRb0FsRR5
RRRRRRqR:MRHR0R#8F_Do_HOP0COFIs5HE80qR-48MFI0jFR2R;
RRRRRRAR:MRHR0R#8F_Do_HOP0COFIs5HE80AR-48MFI0jFR2R;
RRRRRRqA:kRF00R#8F_Do_HOP0COFIs5HE80AH*I8q0E-84RF0IMF2Rj
RRRR-RR-RRA*
RqR2RR;M
C8HRwsu#0skF8O;0#
s
NO0EHCkO0sNCRs4OERRFVw#Hs0Fus80kO##RH
R
RRo#HMRNDNk_NGRR:#_08DHFoOC_POs0F58IH0-Eq4FR8IFM0R;j2
RRR#MHoNLDR_GNkR#:R0D8_FOoH_OPC05FsI0H8E4A-RI8FMR0Fj
2;LHCoMR
RRsVFNqM8:FRVsNRHRRHMjFR0R8IH0-Eq.CRoMNCs0RC
RRRRRsVFNAM8:FRVsLRHRRHMjFR0R8IH0-EA.CRoMNCs0RC
RRRRRRRRqIA5HE80AN*HRH+RL<2R=5RNHRN2NRM8LL5H2R;
RRRRR8CMRMoCC0sNCFRVs8NMAR;
RRRRR_HVCRJ:H5VRH=NRRRj2oCCMsCN0
RRRRRRRRARq58IH0-EA4<2R=5RNjN2RML8R58IH0-EA4
2;RRRRRMRC8CRoMNCs0HCRVJ_C;R
RRRRRHMV_CRJ:H5VRH/NR=2RjRMoCC0sNCR
RRRRRRqRRAH5I8A0E*+HNI0H8E4A-2=R<RF5M05RNH2N2R8NMRIL5HE80A2-4;R
RRRRRCRM8oCCMsCN0R_HVM;CJ
RRRCRM8oCCMsCN0RsVFNqM8;R
RRsVFNAM8:FRVsLRHRRHMjFR0R8IH0-EA.CRoMNCs0RC
RRRRR5qAI0H8E5A*I0H8E4q-2RR+HRL2<N=R58IH0-Eq4N2RM58RMRF0LL5H2
2;RCRRMo8RCsMCNR0CVNFsM;8A
RRRRqRRAH5I8A0E*H5I8q0E-R42+HRI8A0E-R42<N=R58IH0-Eq4N2RML8R58IH0-EA4
2;CRM8NEsO4
;
-*-R*************************************************************R**R
---N-R8C8so,5qRRA,)2C#

---v-RF#PCRosCHC#0s0#RFCRsbODNCHRbbkCLV
'#-
-R-*-R*************************************************************R**R
--
LDHs$NsRCHCC
;RkR#CHCCC38#0_oDFH4O_43ncN;DD
Ck#RCHCC03#8F_Do_HOkHM#o8MC3DND;D

HNLssF$RsdON;#
kCsRFO3NdFNsOObFl3DND;D

HNLss#$R$DMbH;V$
Ck#RM#$bVDH$03N0LsHk#0C3DND;C

M00H$8RN8osCR
H#RoRRCsMCH
O5RRRRRHRI8R0ERH:RMo0CC
s;RRRRRHRI8q0ERH:RMo0CC
s;RRRRRMRH8RCGRH:RMo0CC
s;RRRRRkRMlsLCRH:RMo0CC
s;RRRRRCRsoRRRRH:RMo0CC-sR-NRhlFCRVER0CCRDP
CDR2RR;R
RRsbF0
R5RRRRRHRBMRR:H#MR0D8_FOoH;R
RRRRRqRRR:MRHR8#0_oDFHPO_CFO0sH5I8-0E4FR8IFM0R;j2
RRRRARRR:RRRRHM#_08DHFoOC_POs0F58IH04E-RI8FMR0Fj
2;RRRRRCR)#RR:FRk0#_08DHFoOC_POs0F58IH04E-RI8FMR0FjR2
R;R2
RRRNs00H0LkC3R\s	NM\RR:HCM0o;Cs
RRRNs00H0LkC3R\sFClPMC_FN_IsRM\:MRH0CCosC;
MN8R8C8so
;
NEsOHO0C0CksRONsEF4RV8RN8osCR
H#
RRR#MHoN)DRCD#k0RR:#_08DHFoOC_POs0F58IH04E-RI8FMR0Fj
2;
oLCHRM
RCR)#0kDRR<=qRR+ARR+O;HM
RRRHjV_:VRHRM5H8RCG>2R4RMoCC0sNCRR
RRRRRsVFDbFFjV:RFHsRRRHMjFR0R8IH0-Eq4CRoMNCs0RC
RRRRRRRRNs00H0LkC3R\s	NM\VRFRosC#RR:DCNLD#RHRosC;R
RRRRRRNRR0H0sLCk0Rs\3CPlFCF_M_sINMF\RVCRso:#RRLDNCHDR#;R4
RRRRLRRCMoH
RRRRRRRRCRsoR#:bCHbL
kVRRRRRRRRRRRRb0FsRblN5R
RRRRRRRRRRRRRRRRRQ>R=R#)Ck5D0H
2,RRRRRRRRRRRRRRRRRRRm=)>RCH#52R
RRRRRRRRRR;R2
RRRRCRRMo8RCsMCNR0CVDFsFjFb;R
RR8CMRMoCC0sNCHRRV;_j
R
RR_HV4H:RVHR5MG8CR4=R2CRoMNCs0
CRRRRRRFRVsFDFbR.:VRFsHMRHR0jRFHRI8q0E-o4RCsMCN
0CRRRRRRRRR0N0skHL0\CR3MsN	F\RVCRsoR#q:NRDLRCDHs#RC
o;RRRRRRRRR0N0skHL0\CR3lsCF_PCMIF_N\sMRRFVs#CoqRR:DCNLD#RHR
4;RRRRRCRLo
HMRRRRRRRRRosC#Rq:bCHbL
kVRRRRRRRRRRRRb0FsRblN5R
RRRRRRRRRRRRRRRRRQ>R=R#)Ck5D0H
2,RRRRRRRRRRRRRRRRRRRm=)>RCH#52R
RRRRRRRRRR;R2
RRRRCRRMo8RCsMCNR0CVDFsF.Fb;R
RR8CMRMoCC0sNCHRRV;_4
R
RR_HV.H:RV.R5*8HMC=GRRlMkL2CsRMoCC0sNCRR
RRRRRsVFDbFFdV:RFHsRRRHMI0H8E0qRFHRI8-0E4CRoMNCs0RC
RRRRRRRRNs00H0LkC3R\s	NM\VRFRosC#:ARRLDNCHDR#CRsoR;
RRRRRRRRNs00H0LkC3R\sFClPMC_FN_IsRM\FsVRCAo#RD:RNDLCRRH#4R;
RRRRRoLCHRM
RRRRRRRRs#CoAb:RHLbCkRV
RRRRRRRRRbRRFRs0l5Nb
RRRRRRRRRRRRRRRRQRRRR=>)kC#DH052R,
RRRRRRRRRRRRRRRRR=mR>CR)#25H
RRRRRRRRRRRR
2;RRRRRMRC8CRoMNCs0VCRFFsDF;bd
RRRCRM8oCCMsCN0RVRH_
.;
RRRHdV_:VRHR*5.HCM8GRR<MLklCRs2oCCMsCN0RR
RRRRRVDFsFcFb:FRVsRRHHIMRHE80qFR0R8IH04E-RMoCC0sNCR
RRRRRRNRR0H0sLCk0Rs\3N\M	RRFVs#CoBRR:DCNLD#RHRosC;R
RRRRRRNRR0H0sLCk0Rs\3CPlFCF_M_sINMF\RVCRsoR#B:NRDLRCDH4#R;R
RRRRRLHCoMR
RRRRRRsRRCBo#:HRbbkCLVR
RRRRRRRRRRFRbsl0RN
b5RRRRRRRRRRRRRRRRRRRQ=)>RCD#k025H,R
RRRRRRRRRRRRRRRRRm>R=R#)C5
H2RRRRRRRRRRRR2R;
RRRRR8CMRMoCC0sNCFRVsFDFb
c;RCRRMo8RCsMCNR0CR_HVdC;
MN8Rs4OE;-

-*R**************************************************************R*R---
--
-RFVDFQs5M0bk,kRm00bk2-
-
R--****************************************************************R-R-
H
DLssN$CRHCRC;
Ck#RCHCC03#8F_Do_HO4c4n3DND;#
kCCRHC#C30D8_FOoH_HNs0NE3D
D;kR#CHCCC38#0_oDFHkO_Mo#HM3C8N;DD
H
DLssN$sRFO;Nd
Ck#ROFsNFd3sOONF3lbN;DD
M
C0$H0RFVDFHsR#R
RRRRRoCCMsRHO5R
RRRRRRRRRRHRI8Q0Eh:RRR0HMCsoCRR:=g
j;RRRRRRRRRRRRI0H8EamzRH:RMo0CC:sR=cR6;R
RRRRRRRRRRkRMlsLCR:RRR0HMCsoCRR:=6R;
RRRRRRRRRIRRHE80qRRR:MRH0CCos=R:R
6;RRRRRRRRRRRRHCM8GRRRRRR:HCM0oRCs:
=4RRRRR;R2
RRRRbRRFRs05R
RRRRRRRRRRMRQbRk0RR:RH#MR0D8_FOoH_OPC05FsI0H8E-Qh4FR8IFM0R;j2
RRRRRRRRRRRR0mkbRk0:kRF00R#8F_Do_HOP0COFIs5HE80m-za4FR8IFM0R
j2RRRRR;R2
RRRRNRR0H0sLCk0Rs\3N\M	RH:RMo0CC
s;SNRR0H0sLCk0Rs\3CPlFCF_M_sINM:\RR0HMCsoC;M
C8DRVF;Fs
s
NO0EHCkO0sNCRs4OERRFVVFDFs#RHRR

RORRFFlbM0CMR8N8s
CoRRRRRMoCCOsHRR5
RRRRRRRRI0H8E:RRR0HMCsoC;R
RRRRRRIRRHE80qRR:HCM0o;Cs
RRRRRRRRMRH8RCGRH:RMo0CC
s;RRRRRRRRRlMkLRCs:MRH0CCosR;
RRRRRRRRsRCoR:RRR0HMCsoCRR--hCNlRRFV0RECDCCPDR
RR2RR;R
RRbRRFRs05R
RRRRRBRHM:MRHR8#0_oDFH
O;RRRRRRRqRRR:H#MR0D8_FOoH_OPC05FsR8IH04E-RI8FMR0Fj
2;RRRRRRRARRR:H#MR0D8_FOoH_OPC05FsR8IH04E-RI8FMR0Fj
2;RRRRRCR)#RR:FRk0#_08DHFoOC_POs0F58IH04E-RI8FMR0FjR2
RRRR2R;
RMRC8FROlMbFC;M0
R
RRb0$CER#H_V00DNLC#RHRsNsN5$RMLklC.s/RI8FMR0FjF2RVMRH0CCos
;
RVRRk0MOHRFM#VEH0sxCFM5H8RCG:MRH0CCoss2RCs0kMER#H_V00DNLC#RH
RRRRPRRNNsHLRDC#b0CRH:RMo0CC
s;RRRRRNRPsLHND0CRNCLD_sPNRRR:#VEH0N_0L;DC
RRRLHCoMR
RRRRR#b0CRR:=4R;
RRRRRsVFRHHRMRR40HFRMG8C-D4RF
FbRRRRRRRRRC#0b=R:RC#0bRR*.R;
RRRRR8CMRFDFbR;
RRRRRsVFRHHRMRRj0MFRkClLsR/.DbFF
RRRRRRRRNR0L_DCP5NsH:2R=0R#C*bRR*5.H2+4;R
RRRRRCRM8DbFF;R
RRRRRskC0s0MRNCLD_sPN;R
RR8CMRH#EVC0xs
F;
RRRO#FM00NMRMDCoR0E:MRH0CCos=R:R8IH0MEQ/lMkL;Cs
RRRO#FM00NMR8IH0REA:MRH0CCos=R:RMDCoR0E-HRI8q0E;R

RFROMN#0M#0RE0HVNC88sRR:#VEH0N_0LRDC:#=RE0HVxFCs58HMC;G2
C
Lo
HMRVRRFFsDF4b_:FRVsRR[H4MRRR0FMLklC.s/RMoCC0sNCR
RRoLCHRM
RRRRRosC#Rq:Ns88CRo
RRRRRMoCCOsHRblNRR5
RRRRR8IH0=ER>CRDMEo0-H#EV80N85Cs[2-4-
4,RRRRRHRI8q0ERR=>I0H8E
q,RRRRRMRH8RCG=[>R,R
RRRRRMLklC=sR>kRMlsLC,R
RRRRRsRCoR>R=R8HMCRG
RRRRRR2
RRRRRsbF0NRlbR5
RRRRRRRRRHRBM>R=RbQMkD05C0MoE.*5*4[-2R2,
RRRRRRRRRRq=Q>RM0bk5MDCo*0E5[.*--424FR8IFM0RMDCo*0E.[*5-+42#VEH08N8C[s5-+424
2,RRRRRRRRR=AR>MRQb5k0DoCM0.E**4[-RI8FMR0FDoCM05E*.-*[4#2+E0HVNC88s-5[442+2R,
RRRRRRRR)RC#=m>Rkk0b0C5DMEo0*4[-RI8FMR0FDoCM05E*[2-4+H#EV80N85Cs[2-4+
42RRRRR;R2
RRRR-RR-NROsRs$VRFs0RECM0CGRFVDFRs
RRRRRsVFDbFF_Rj:VRFsHMRHR0jRFER#HNV08s8C54[-2E-#HNV08s8C5Rj2oCCMsCN0
RRRRRRRRRRRRRRRmbk0kD05C0MoE[*5-+42RRH2<'=Rj
';RRRRRMRC8CRoMNCs0VCRFFsDFjb_;R

RRRRRR--NCDsNR8$oCCMsCN08R
RRRRRVDFsF_FbNV:RFHsRRRHMjFR0RH#EV80N85Csj42-RMoCC0sNCR
RRRRRRNRR0H0sLCk0Rs\3N\M	RRFVs#CoRD:RNDLCRRH#HCM8GR;
RRRRRRRRNs00H0LkC3R\sFClPMC_FN_IsRM\FsVRCRo#:NRDLRCDH4#R;R
RRRRRLHCoMR
RRRRRRsRRC:o#RbbHCVLk
RRRRRRRRRRRRRRRb0FsRblN5R
RRRRRRRRRRRRRRRRRRQRRRR=>QkMb0C5DMEo0*5.*[2-4+H#EV80N85Cs[2-4-H#EV80N85Csj42++,H2
RRRRRRRRRRRRRRRRRRRRRRm=m>Rkk0b0C5DMEo0*-5[4H2++H#EV80N85Cs[2-4-H#EV80N85Csj42+2R
RRRRRRRRRRRRRRRRRR2RR;R
RRRRRCRM8oCCMsCN0RsVFDbFF_
N;
RRRCRM8oCCMsCN0RsVFDbFF_
4;
RRRH#V_FNk#:VRHRk5MlsLCR8lFR=.RRR42oCCMsCN0
RRRRNRR0H0sLCk0Rs\3N\M	RRFVsOCoN$ss#RR:DCNLD#RHR8HMC
G;RRRRR0RN0LsHkR0C\C3slCFP__MFIMNs\VRFRosCOsNs$:#RRLDNCHDR#;R4
RRRLHCoMR
RRRRRVDFsF_FbdV:RFHsRRRHM4FR0RCRDMEo0-H#EV80N85CsMLklC.s/2+-4#VEH08N8Cjs52CRoMNCs0RC
RRRRR0N0skHL0\CR3MsN	F\RVCRso:#RRLDNCHDR#MRH8;CG
RRRRNRR0H0sLCk0Rs\3CPlFCF_M_sINMF\RVCRso:#RRLDNCHDR#;R4
RRRRLRRCMoH
RRRRRRRRCRsoR#:bCHbL
kVRRRRRRRRRsbF0NRlbR5
RRRRRRRRRQRRRR=>QkMb0H5I8Q0Eh2-H,R
RRRRRRRRRRRRm=m>Rkk0b0H5I8m0EzHa-2R
RRRRRR2RR;R
RRRRRCRM8oCCMsCN0RsVFDbFF_
d;RRRRRCRsosONs:$#RbbHCVLk
RRRRRRRRFRbsl0RN
b5RRRRRRRRRRRRQ>R=RbQMkI05HE80QDh-C0MoE
2,RRRRRRRRRRRRm>R=R0mkb5k0I0H8Eamz-MDCo20E
RRRRRRRR;R2
RRRRmRRkk0b0H5I8m0EzDa-C0MoEE+#HNV08s8C5lMkL/Cs.#2-E0HVNC88s25jRI8FMR0FI0H8Eamz-MDCo+0E4<2R=RR
RRRRRRRRRRRRRMRQb5k0I0H8E-QhDoCM0#E+E0HVNC88sk5MlsLC/-.2#VEH08N8Cjs52FR8IFM0R8IH0hEQ-MDCo+0E4R2;
RRRCRM8oCCMsCN0R_HV##FkNC;
MN8Rs4OE;D

HNLssH$RC;CCR#
kCCRHC#C30D8_FOoH_n44cD3NDk;
#HCRC3CC#_08DHFoOs_NH30EN;DD
Ck#RCHCC03#8F_Do_HOkHM#o8MC3DND;D

HNLssF$RsdON;#
kCsRFO3NdFNsOObFl3DND;C

M00H$DRVF_FsNC88s#RH
RRRRoRRCsMCH5OR
RRRRRRRRRRRR8IH0hEQRRR:HCM0oRCs:g=RjR;
RRRRRRRRRIRRHE80mRza:MRH0CCos=R:R;6c
RRRRRRRRRRRRlMkLRCsRRR:HCM0oRCs:6=R
RRRR2RR;R
RRRRRb0FsRR5
RRRRRRRRRQRRM0bkRRR:RRHM#_08DHFoOC_POs0F58IH0hEQ-84RF0IMF2Rj;R
RRRRRRRRRRkRm00bkRF:Rk#0R0D8_FOoH_OPC05FsI0H8Eamz-84RF0IMF2Rj
RRRR2RR;M
C8DRVF_FsNC88s
;
NEsOHO0C0CksRONsEF4RVDRVF_FsNC88s#RHRR
RRMOF#M0N0CRDMEo0RH:RMo0CC:sR=HRI8Q0EMk/MlsLC;C
Lo
HMRVRRFFsDF4b_:FRVsRR[H4MRRR0FMLklC.s/RMoCC0sNCR
RRRRRmbk0kD05C0MoE-*[4FR8IFM0RMDCo*0E54[-22+4RR<=RbQMkD05C0MoE.*5*4[-2R-48MFI0DFRC0MoE**.54[-22+4
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR+MRQb5k0DoCM0.E**4[-RI8FMR0FDoCM05E*.-*[442+2R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRQ+RM0bk5MDCo*0E5[.*-242;R

RRRRR0mkb5k0DoCM05E*[2-42=R<R''j;R
RR8CMRMoCC0sNCFRVsFDFb;_4
R
RR_HV##FkNH:RVMR5kClLsFRl8RR.=2R4RMoCC0sNCR
RRRRRmbk0kI05HE80m-za4FR8IFM0R8IH0zEmaC-DMEo02=R<RbQMkI05HE80Q4h-RI8FMR0FI0H8E-QhDoCM0;E2RR
RR8CMRMoCC0sNCVRH_k#F#
N;
8CMRONsE
4;
LDHs$NsRCHCC
;RkR#CHCCC38#0_oDFH4O_43ncN;DD
Ck#RCHCC03#8F_Do_HON0sHED3NDk;
#HCRC3CC#_08DHFoOM_k#MHoCN83D
D;
0CMHR0$NC88sCasCH.R#R
RRMoCCOsH5R
RRRRRI0H8E:qRR0HMCsoC;R
RRRRRI0H8E:ARR0HMCsoC;R
RRRRR0CsCR:RRR0HMCsoC
RRR2R;
RFRbs50R
RRRRqRR,lRq,RRA:MRHR8#0_oDFH
O;RRRRRARqRRR:H#MR0D8_FOoH_OPC05FsI0H8EIA*HE80qR-48MFI0jFR2R;
RRRRRFbs80kORF:Rk#0R0D8_FOoH_OPC05FsI0H8EIA+HE80qR-48MFI0jFR2R
RRRRR-A-RRq*R
RRR2C;
MN8R8s8CaCsC.R;

ONsECH0Os0kCsRNORE4FNVR8s8CaCsC.#RH
RRRO#FM00NMRC0EEEHoR#:R0D8_FOoH_OPC05Fs486RF0IMF2RjRR:=Bemh_71a_tpmQeB_ mBa)H5I8q0E-R4,4;n2
RRRObFlFMMC0DRVF
FsRRRRRCRoMHCsO
R5RRRRRRRRR8IH0hEQRRR:HCM0oRCs;R
RRRRRRIRRHE80mRza:MRH0CCos
R;RRRRRRRRRlMkLRCsRRR:HCM0oRCs;R
RRRRRRIRRHE80qRRR:MRH0CCos
R;RRRRRRRRR8HMCRGRRRR:HCM0o
CsRRRRR;R2
RRRRRRRb0FsRR5
RRRRRRRRRRRRRbQMkR0R:MRHR8#0_oDFHPO_CFO0sH5I8Q0EhR-48MFI0jFR2R;
RRRRRRRRRRRRR0mkbRk0:kRF00R#8F_Do_HOP0COFIs5HE80m-za4FR8IFM0R
j2RRRRR2RR;R
RR8CMRlOFbCFMM
0;
RRRObFlFMMC0DRVF_FsNC88sR
RRRRRoCCMsRHO5R
RRRRRRIRRHE80QRhR:MRH0CCos
R;RRRRRRRRR8IH0zEmaRR:HCM0oRCs;R
RRRRRRMRRkClLsRRR:MRH0CCosR
RRRRR2R;
RRRRRFRbs50R
RRRRRRRRRRRRQRRM0bkRRR:H#MR0D8_FOoH_OPC05FsI0H8E-Qh4FR8IFM0R;j2
RRRRRRRRRRRRmRRkk0b0RR:FRk0#_08DHFoOC_POs0F58IH0zEmaR-48MFI0jFR2R
RRRRRR
2;RCRRMO8RFFlbM0CM;R

RkRVMHO0F8MRCEb0W0H8ECRs0MksR0HMCsoCR
H#RLRRCMoH
RRRRFRVsRRHH4MR6FR8IFM0RDjRF
FbRHRRV0R5EHCEoHE52RR='24'RC0EMR
RRRRRskC0sHMR+
4;RCRRMH8RVR;
RRRRCRM8DbFF;R
RRsRRCs0kM;Rj
RRRCRM880CbE8WH0
E;
RRRO#FM00NMRb8C0:ERR0HMCsoCRR:=80CbE8WH0
E;RORRF0M#NRM0I0H8E:0RR0HMCsoCRR:=I0H8EIA+HE80q;+.
RRR0C$bRlDH##RHRsNsN5$R80CbER+48MFI0jFR2VRFR0HMCsoC;

RRVRRk0MOHRFMOONDhLklCRs#skC0sDMRHRl#HR#
RRRRRsPNHDNLCER0Ck_MlsLC#RR:D#Hl;R
RRoLCHRM
RRRRRC0E_lMkL#Cs5Rj2:I=RHE80qR;
RRRRRsVFRHHRMRR408FRCEb0+D4RF
FbRRRRRRRRRC0E_lMkL#Cs5RH2:0=REMC_kClLsH#5-/42.RR+5C0E_lMkL#Cs54H-2FRl82R.;R
RRRRRCRM8DbFF;R
RRRRRskC0s0MREMC_kClLs
#;RRRRCRM8OONDhLklC;s#
RR
RFROMN#0MM0RkClLs:#RRlDH#=R:RDONOlhkL#Cs;

RRVRRk0MOHRFMOONDpRHlskC0sDMRHRl#HR#
RRRRRsPNHDNLCER0CH_Dl:#RRlDH#R;
RRRRRsPNHDNLCkRMl:LRR0HMCsoC;R
RRoLCHRM
RRRRRC0E_lDH#25jRR:=jR;
RRRRRlMkL=R:R8IH0;Eq
RRRRVRRFHsRRRHM4FR0Rb8C04E+RFDFbR
RRC0E_lDH#25HRR:=0_ECD#Hl54H-2RR+MLkl*8IH0;E0
RRRMLklRR:=MLkl/+.RRk5MllLRF.8R2R;
RRRRR8CMRFDFbR;
RRRRR0sCkRsM0_ECD#Hl;R
RRMRC8NRODHOplR;

RRRO#FM00NMROPCDRHl:HRDl:#R=NRODHOplR;
RHR#oDMNRoLH0CsCR#:R0D8_FOoH_OPC05FsPDCOH8l5CEb0+-424FR8IFM0R;j2
RRR#MHoNODRN$ss,HR#oRM,#MHo4RR:#_08DHFoO
;
LHCoMRR
RVRH_C	Cb8_N8aCss:CCRRHV5C0sCRR=jo2RCsMCNR0C-k-R#VCRFbsRHDbCHMMHoMRN8FRDIFRO#
0
RRRRRHR#o<MR=RRqGRFsAR;
RRRRRo#HM<4R=RRqFAsR;R
RRRRROsNs$=R<RF5M0lRq2MRN8;RA
RRRRLRRHso0CIC5HE800R-48MFI0jFR2=R<RmRBh1e_ap7_mBtQ_Be a5m)jI,RHE80qR2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRO&RN$ss
RRRRRRRRRRRRRRRRRRRRRRRRRRRR&RRR5qAI0H8E4A-RI8FMR0FjR2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRB&Rm_he1_a7pQmtB _eB)am5Rj,4
2;
RRRRVRRFMsN8Rq:VRFsHHNRMRR40IFRHE80qR-doCCMsCN0
RRRRRRRRHRLoC0sCH55N2+4*8IH0-E04FR8IFM0R*HNI0H8ER02<R=RBemh_71a_tpmQeB_ mBa),5jR8IH0+Eq4N-H2R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR&ARq58IH0*EA5+HN442-RI8FMR0FI0H8EHA*NR2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRB&Rm_he1_a7pQmtB _eB)am5Rj,H4N+2R;
RRRRR8CMRMoCC0sNCFRVs8NMqR;
RRRRRR--FRMCLFCVs0CREDCRNR#0P0COFRs
RRRRRoLH0CsC5H5I8q0E-*42I0H8E40-RI8FMR0F58IH0-Eq.I2*HE800<2R=BRRm_he1_a7pQmtB _eB)am5Rj,.R2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR&RRRo#HMR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR&qIA5HE80AI*5HE80q2-4-84RF0IMFHRI8A0E*H5I8q0E-2.2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRB&Rm_he1_a7pQmtB _eB)am5Rj,I0H8E4q-2R;
RRRRRR--D0N#ROPC0
FsRRRRRHRLoC0sCH5I8q0E*8IH0-E04FR8IFM0RH5I8q0E-*42I0H8ER02<
=RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRBemh_71a_tpmQeB_ mBa),5jR
42RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR#&RH4oM
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR&qIA5HE80AH*I8q0E-84RF0IMFHRI8A0E*H5I8q0E-242
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR&Bemh_71a_tpmQeB_ mBa),5jR8IH0-Eq4R2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR&;Rq
R
RRRRRVDFsF.Fb:sVFRH[RMRR408FRCEb0RMoCC0sNCR
RRRRRRlRR4R:RVFDFsR
RRRRRRRRRRCRoMHCsONRlb
R5RRRRRRRRRRRRRRRRRRRRR8IH0hEQR>R=ROPCD5Hl[-2RROPCD5Hl[2-4,R
RRRRRRRRRRRRRRRRRRIRRHE80mRza=P>RCHODl+5[4-2RROPCD5Hl[
2,RRRRRRRRRRRRRRRRRRRRRlMkLRCsR>R=RlMkL#Cs54[-2R,
RRRRRRRRRRRRRRRRRRRRI0H8ERqRRR=>I0H8E
q,RRRRRRRRRRRRRRRRRRRRR8HMCRGRR>R=RR[
RRRRRRRRR2RR
RRRRRRRRRRRRsbF0NRlb
R5RRRRRRRRRRRRRRRRRRRRRbQMkR0RR>R=RoLH0CsC5OPCD5Hl[42-RI8FMR0FPDCOH[l5-242,R
RRRRRRRRRRRRRRRRRRmRRkk0b0RRR=L>RHso0CPC5CHODl+5[442-RI8FMR0FPDCOH[l52R2
RRRRRRRRR2RR;R
RRRRRCRM8RMoCC0sNCFRVsFDFb
.;RCRRMo8RCsMCNR0CH	V_C_CbNC88sCasC
;
RHRRVF_M0C	Cb8_N8aCss:CCRRHV5C0sCRR=4o2RCsMCNR0C-k-R#HCRV8RN8RCsNCV0sER0CkRlDb0HDsHC
RRRR-RR-HRI8q0ERR>=cR
RRRRR#MHoR=R<RGqRFAsR;R
RRRRR#MHo4=R<RFqRs;RA
RRRRORRN$ssRR<=50MFR2qlR8NMR
A;RRRRRHRLoC0sCH5I800E-84RF0IMF2RjRR<=RhBmea_17m_pt_QBea Bmj)5,HRI8q0E2R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR&NROs
s$RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR&qIA5HE80AR-48MFI0jFR2R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR&mRBh1e_ap7_mBtQ_Be a5m)j4,R2
;
RRRRRVRH_8IH0:EqRRHV58IH0REq>2RdRMoCC0sNCR
RRRRRRLRRHso0C.C5*8IH0-E04FR8IFM0R8IH02E0RR<=RhBmea_17m_pt_QBea Bmj)5,HRI8q0E2R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRq&RA*5.I0H8E4A-RI8FMR0FI0H8E
A2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR&RRRRq
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR&q
;
RRRRRRRRRsVFNqM8:FRVsNRHRRHM.FR0R8IH0-EqdCRoMNCs0RC
RRRRRRRRRLRRHso0C5C5H4N+2H*I800E-84RF0IMFNRH*8IH02E0RR<=RhBmea_17m_pt_QBea Bmj)5,HRI8q0E+H4-NR2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR&ARq58IH0*EA5+HN442-RI8FMR0FI0H8EHA*NR2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR&
RqRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRB&Rm_he1_a7pQmtB _eB)am5Rj,H;N2
RRRRRRRRMRC8CRoMNCs0VCRFMsN8
q;RRRRRRRRRR--FRMCLFCVs0CREDCRNR#0P0COFRs
RRRRRRRRL0Hos5CC58IH0-Eq4I2*HE800R-48MFI05FRI0H8E.q-2H*I800E2=R<RmRBh1e_ap7_mBtQ_Be a5m)j.,R2R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR#&RH
oMRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR&RRR5qAI0H8E5A*I0H8E4q-2R-48MFI0IFRHE80AI*5HE80q2-.2R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRq&R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR&mRBh1e_ap7_mBtQ_Be a5m)jI,RHE80q2-.;R
RRRRRCRM8oCCMsCN0R_HVI0H8E
q;
RRRRHRRVH_I8q0E_Rj:H5VRI0H8E=qRRRd2oCCMsCN0
RRRRRRRR-R-RCFMRVLCFRsC0RECD0N#ROPC0
FsRRRRRRRRRoLH0CsC5I.*HE800R-48MFI0IFRHE800<2R=BRRm_he1_a7pQmtB _eB)am5Rj,.R2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR&#MHo
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR&ARq5I.*HE80AR-48MFI0IFRHE80AR2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR&qR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRq&R;R

RRRRR8CMRMoCC0sNCVRH_8IH0_EqjR;
RRRRRR--D0N#ROPC0
FsRRRRRHRLoC0sCH5I8q0E*8IH0-E04FR8IFM0RH5I8q0E-*42I0H8ER02<R=RBemh_71a_tpmQeB_ mBa),5jR
42RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR#&RH4oM
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR&qIA5HE80AH*I8q0E-84RF0IMFHRI8A0E*H5I8q0E-242
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR&qR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR&RRRhBmea_17m_pt_QBea Bmj)5,HRI8q0E-;42
R
RRRRRVDFsFdFb:sVFRH[RMRR408FRCEb0RMoCC0sNCR
RRRRRRlRR4R:RVFDFs8_N8
CsRRRRRRRRRRRRoCCMsRHOlRNb5R
RRRRRRRRRRRRRRRRRRIRRHE80QRhR=P>RCHODl25[RP-RCHODl-5[4
2,RRRRRRRRRRRRRRRRRRRRR8IH0zEma>R=ROPCD5Hl[2+4RP-RCHODl25[,R
RRRRRRRRRRRRRRRRRRMRRkClLsRRR=M>RkClLs[#5-
42RRRRRRRRRRRR2R
RRRRRRRRRRFRbsl0RN5bR
RRRRRRRRRRRRRRRRRRRRMRQbRk0R=RR>HRLoC0sCC5POlDH5-[24FR8IFM0ROPCD5Hl[2-42R,
RRRRRRRRRRRRRRRRRRRRmbk0kR0RRR=>L0Hos5CCPDCOH[l5+-424FR8IFM0ROPCD5Hl[
22RRRRRRRRRRRR2R;
RRRRR8CMRCRoMNCs0VCRFFsDF;bd
RRRCRM8oCCMsCN0R_HVM	F0C_CbNC88sCasC
;
RbRRskF8O<0R=HRLoC0sCC5POlDH5b8C04E+2R-.8MFI0PFRCHODlC58b20E+;42RC

MN8Rs4OE;D

HNLssH$RC;CC
Ck#RCHCC03#8F_Do_HO4c4n3DND;#
kCCRHC#C30D8_FOoH_HNs0NE3D
D;kR#CHCCC38#0_oDFH#O_HCoM8D3ND
;
DsHLNRs$FNsOdk;
#FCRsdON3OFsNlOFbD3ND
;
DsHLNRs$#b$MD$HV;#
kC$R#MHbDVN$30H0sLCk0#D3ND
;
CHM00#$RlDNDv0kDR
H#RoRRCsMCH
O5RRRRRIRNHE80RH:RMo0CC:sR=;Rg
RRRRLRRI0H8ERR:HCM0oRCs:g=R;R
RRRRRI0H8E:RRR0HMCsoCRR:=4RU
R;R2
RRRb0FsRR5
RRRRRRqRRRR:HRMR#_08DHFoOC_POs0F5HNI8-0E4FR8IFM0R;j2
RRRRARRRRRR:MRHR0R#8F_Do_HOP0COFLs5I0H8ER-48MFI0jFR2R;
RRRRRmu)7RR:FRk0#_08DHFoOC_POs0F58IH04E-RI8FMR0FjR2
RRRRRR--ARR*qR
RR
2;RNRR0H0sLCk0Rs\3CPlFCF_M_sINM:\RR0HMCsoC;R
RR0N0skHL0\CR3MsN	:\RR0HMCsoC;M
C8lR#NvDDk;D0
s
NO0EHCkO0sNCRs4OERRFV#DlNDDvk0#RH
R
RRMVkOF0HMkR#bH5I8N0E,HRI8L0ERH:RMo0CCRs2skC0sHMRMo0CCHsR#R
RRoLCHRM
RRRRRRHV58IH0REN>HRI8L0E2ER0CRM
RsRRCs0kMHRI8N0E;R
RRRRRCCD#
RRRR0sCkRsMI0H8E
L;RRRRRMRC8VRH;R
RR8CMRb#k;R

RkRVMHO0FHMRMIV5HE80NI,RHE80LRR:HCM0o2CsR0sCkRsMHCM0oRCsHR#
RCRLo
HMRRRRRVRHRH5I8N0ERI<RHE80L02RE
CMRRRRskC0sIMRHE80NR;
RRRRR#CDCR
RR0sCkRsMI0H8E
L;RRRRRMRC8VRH;R
RR8CMRVHM;R

RFROMN#0MI0RHE80qRR:HCM0oRCs:H=RMNV5I0H8EL,RI0H8E
2;RORRF0M#NRM0I0H8E:ARR0HMCsoCRR:=#5kbN8IH0RE,L8IH0;E2
R
RRlOFbCFMMw0RH0s#u8sFk#O0
oSSCsMCH
O5SISSHE80qRR:HCM0o;Cs
SSSI0H8E:ARR0HMCsoC
SSS2S;
SsbF0
R5SqSSRRR:HRMR#_08DHFoOC_POs0F5HNI8-0E4FR8IFM0R;j2
SSSA:RRRRHMR8#0_oDFHPO_CFO0sI5LHE80-84RF0IMF2Rj;S
SSRqA:kRF00R#8F_Do_HOP0COFLs5I0H8EI*NHE80-84RF0IMF2Rj
SSS-A-RRq*R
SSS2R;
RMRC8FROlMbFC;M0
R
RRlOFbCFMMN0R8s8CaCsC.S
SoCCMs5HO
SSSI0H8E:qRR0HMCsoC;S
SS8IH0REA:MRH0CCosS;
SsS0CRCRRH:RMo0CCSs
S;S2
bSSFRs05S
SSRq,qRl,ARR:H#MR0D8_FOoH;S
SSRqARH:RM0R#8F_Do_HOP0COFLs5I0H8EI*NHE80-84RF0IMF2Rj;S
SSFbs80kORF:Rk#0R0D8_FOoH_OPC05FsL8IH0NE+I0H8ER-48MFI0jFR2S
SSR--ARR*qS
SS
2;RCRRMO8RFFlbM0CM;R

RHR#oDMNRNN_k:GRR8#0_oDFHPO_CFO0sH5I8q0E-84RF0IMF2Rj;R
RRo#HMRNDLk_NGRR:#_08DHFoOC_POs0F58IH0-EA4FR8IFM0R;j2
RRR#MHoNNDRLRRRR#:R0D8_FOoH_OPC05FsN8IH0LE*I0H8ER-48MFI0jFR2R;
RHR#oDMNR#)Ck:D0R8#0_oDFHPO_CFO0sI5NHE80+HLI8-0E4FR8IFM0R;j2
oLCH
MRR-RR-IR1NqbRR8NMRHARVCRMO#C#N
s$RHRRVNqDssoCAH:RVNR5I0H8ERR>L8IH0RE2oCCMsCN0
RRRRVRRFFsDF:b.RsVFRHHRMRRj0LFRI0H8ER-4oCCMsCN0
RRRRRRRR0RN0LsHkR0C\N3sMR	\FsVRCqo#RD:RNDLCRRH#jR;
RRRRRRRRNs00H0LkC3R\sFClPMC_FN_IsRM\FsVRCqo#RD:RNDLCRRH#4R;
RRRRRRRRNs00H0LkC3R\s	NM\VRFRosC#:ARRLDNCHDR#;Rj
RRRRRRRR0RN0LsHkR0C\C3slCFP__MFIMNs\VRFRosC#:ARRLDNCHDR#;R4
RRRRLRRCMoH
RRRRsRRCqo#:HRbbkCLVR
RRRRRb0FsRblN5R
RRRRRRQRRRR=>A25H,R
RRRRRRmRRRR=>Nk_NG25H
RRRR2RR;R
RRRRRs#CoAb:RHLbCkRV
RRRRRsbF0NRlbR5
RRRRRRRRQ>R=RHq52R,
RRRRRRRRm>R=RNL_kHG52R
RRRRR2R;
RRRRR8CMRMoCC0sNCFRVsFDFb
.;RRRRRFRVsFDFbR4:VRFsHMRHRHLI8R0E0NFRI0H8ER-4oCCMsCN0
RRRRRRRR0RN0LsHkR0C\N3sMR	\FsVRCAo#RD:RNDLCRRH#jR;
RRRRRRRRNs00H0LkC3R\sFClPMC_FN_IsRM\FsVRCAo#RD:RNDLCRRH#4R;
RRRRRoLCHRM
RRRRRosC#RA:bCHbL
kVRRRRRFRbsl0RN
b5RRRRRRRRR=QR>5RqH
2,RRRRRRRRR=mR>_RLN5kGHR2
RRRRR
2;RRRRRMRC8CRoMNCs0VCRFFsDF;b4
RRRCRM8oCCMsCN0RqHVDoNsC;sA
R
RRqHV#DlNDACs:VRHRI5NHE80RR<=L8IH0RE2oCCMsCN0
RRRRVRRFFsDF:bNRsVFRHHRMRRj0NFRI0H8ER-4oCCMsCN0
RRRRRRRR0RN0LsHkR0C\N3sMR	\FsVRCBo#RD:RNDLCRRH#jR;
RRRRRRRRNs00H0LkC3R\sFClPMC_FN_IsRM\FsVRCBo#RD:RNDLCRRH#4R;
RRRRRRRRNs00H0LkC3R\s	NM\VRFRosC#:1RRLDNCHDR#;Rj
RRRRRRRR0RN0LsHkR0C\C3slCFP__MFIMNs\VRFRosC#:1RRLDNCHDR#;R4
RRRRLRRCMoH
RRRRsRRCBo#:HRbbkCLVR
RRRRRb0FsRblN5R
RRRRRRQRRRR=>q25H,R
RRRRRRmRRRR=>Nk_NG25H
RRRR2RR;R
RRRRRs#Co1b:RHLbCkRV
RRRRRsbF0NRlbR5
RRRRRRRRQ>R=RHA52R,
RRRRRRRRm>R=RNL_kHG52R
RRRRR2R;
RRRRR8CMRMoCC0sNCFRVsFDFb
N;RRRRRFRVsFDFbRL:VRFsHMRHRHNI8R0E0LFRI0H8ER-4oCCMsCN0
RRRRRRRR0RN0LsHkR0C\N3sMR	\FsVRC7o#RD:RNDLCRRH#jR;
RRRRRRRRNs00H0LkC3R\sFClPMC_FN_IsRM\FsVRC7o#RD:RNDLCRRH#4R;
RRRRRoLCHRM
RRRRRosC#R7:bCHbL
kVRRRRRFRbsl0RN
b5RRRRRRRRR=QR>5RAH
2,RRRRRRRRR=mR>_RLN5kGHR2
RRRRR
2;RRRRRMRC8CRoMNCs0VCRFFsDF;bL
RRRCRM8oCCMsCN0RqHV#DlNDACs;R

RHRws1#00:CbRswH#s0uFO8k0R#
RCRoMHCsONRlb
R5RRRRRHRI8q0ERR=>I0H8E
q,RRRRRHRI8A0ERR=>I0H8ERA
R
R2RbRRFRs0lRNb5R
RRRRRq>R=RNN_k
G,RRRRRRRA=L>R_GNk,R
RRRRRq=AR>LRN
RRR2
;
RqRR8s8CaCsCRN:R8s8CaCsC.R
RRMoCCOsHRblNRR5
RRRRR8IH0REq=I>RHE80qR,
RRRRR8IH0REA=I>RHE80AR,
RRRRRC0sCRRR=j>RRRRRR-RR-RR4HNVR8s8CR0NVC0sRElCRkHD0bCDHsj,RR#CDCR
RRR2
RFRbsl0RN5bR
RRRRqRRl>R=RNN_kjG52R,
RRRRRRqR=N>R_GNk58IH0-Eq4
2,RRRRRRRARR=>Lk_NGH5I8A0E-,42
RRRRqRRA>R=R,NL
RRRRbRRskF8O=0R>CR)#0kD
RRR2
;
RHRRVF_I:VRHRH5I8R0E<I=RHE80qRR+I0H8ERA2oCCMsCN0
RRRRuRR)Rm7<)=RCD#k0H5I8-0E4FR8IFM0R;j2
RRRCRM8oCCMsCN0R_HVI
F;RHRRV4_I:VRHRH5I8R0E>HRI8q0ERI+RHE80Ao2RCsMCN
0CRRRRR)RumI75HE80qH+I8A0E-84RF0IMF2RjRR<=)kC#DI05HE80qH+I8A0E-84RF0IMF2Rj;R
RRRRRV_FsDbFF_RI:VRFsHMRHR8IH0+EqI0H8E0ARFHRI8-0E4CRoMNCs0RC
RRRRRRRRu7)m5RH2<)=RCD#k0H5I8q0E+8IH0-EA4
2;RRRRRMRC8CRoMNCs0VCRFDs_F_FbIR;
RMRC8CRoMNCs0HCRV4_I;M
C8sRNO;E4
-
-R****************************************************************-RR--
-RAe.pimB5Rq,Au,R)2m7

---N-RI0H8ERR-I0H8EVRFRHqRM0bk
R--L8IH0-ERR8IH0FERVRRAHkMb0-
-R-
-Rmu)7RR-aRECVDkDRFbs80kORI5NHE80RL+RI0H8EHRI8RC2VlsFRFLDOl	RkHD0bCDHsR#3
R--
R--****************************************************************R-R-
H
DLssN$CRHC
C;kR#CHCCC38#0_oDFH4O_43ncN;DD
Ck#RCHCC03#8F_Do_HON0sHED3NDk;
#HCRC3CC#_08DHFoOM_k#MHoCN83D
D;
LDHs$NsROFsN
d;kR#CFNsOds3FOFNOlNb3D
D;
0CMHR0$ep.AmRBiHS#
oCCMsRHO5S
SSHNI8R0E:MRH0CCosS;
SISLHE80RH:RMo0CC
s;SMSSC_C8bCHbL#kVRH:RMo0CC;s2
FSbs50R
qSSRRRR:MRHR0R#8F_Do_HOP0COFNs5I0H8ER-48MFI0jFR2S;
SRARRRR:HRMR#_08DHFoOC_POs0F5HLI8-0E4FR8IFM0R;j2
uSS)Rm7:kRF00R#8F_Do_HOP0COFNs5I0H8EI+LHE80-84RF0IMF2Rj2S;
Ns00H0LkC3R\s	NM\RR:HCM0o;Cs
0SN0LsHkR0C\C3slCFP__MFIMNs\RR:HCM0o;Cs
0SN0LsHkR0C\C3Lo_HM0CsC\RR:HCM0o;Cs
0SN0LsHkR0C\M3H0MCsNHD_MN#0MN0H0\C8RH:RMo0CC
s;CRM8ep.Am;Bi
s
NO0EHCkO0sLCRD	FO#VRFRAe.pimBR
H#
-S-RlqRNlGHkVlRk0MOHRFMM8CCCI8RERCMN8IH0HER#FRM0JRCkRND0LFRI0H8E-
S-kRbs#bFCV:RHRM80REC#NJksNCRs$sNR8IH0VERsRFl0RECHkMb0kRL#HR#x
C#RVRRk0MOHRFMlN$lGPR5NCDkNP,RNCDkLRR:HCM0o2Cs
sSSCs0kMMRH0CCos#RH
CSLoRHMRR--lN$lGS
SHPVRNCDkNRR>PkNDC0LRE
CMSsSSCs0kMNRPDNkC;S
SCCD#
SSSskC0sPMRNCDkLS;
S8CMR;HV
MSC8$Rll;NG
-
S-kRbs#bFCB:RNkDODCN0RC0ER8HMCHGRMER0CsRuFO8k0sRqsRN$F0VRECCRM$0s
-S-RN0E0CR80lCsH#MCRC0ERo#HMHRL0FRVsER0CkROsMsC0FRsI
3RRVRRk0MOHRFM1MHoAODF	
R5RRRRRFROMN#0MI0RH,8NR8IHLH,R8:GRR0HMCsoC2S
SskC0sHMRMo0CCHsR#L
SCMoHR-R-Ro1HMFADOS	
SRHV58IHN2-4-GH8RI<RHR8L0MEC
SSSskC0s5MR58IHL2+4*H5I84N-28-HG
2;SDSC#SC
SCSs0MksRH5I85L*ILH8+GH822-4;S
SCRM8H
V;S8CMRo1HMFADO
	;
RRRObFlFMMC0zRvpUa4X_4U Rv
RRRRRsbF0
R5S4Sq(q,R4Rn,q,46Rcq4,4Rqdq,R4R.,q,44Rjq4,gRqRRRRRRRRRH:RM0R#8F_DoRHO;S
SqRU,qR(,qRn,qR6,qRc,qRd,qR.,qR4,qSjSSRSRRH:RM0R#8F_DoRHO;S
SA,4(RnA4,4RA6A,R4Rc,A,4dR.A4,4RA4A,R4Rj,ARgRRRRRR:RRRRHM#_08DHFoO
R;SUSA,(RA,nRA,6RA,cRA,dRA,.RA,4RA,jRASSSSR:RRRRHM#_08DHFoO
R;
RSRRdRu6u,RdRc,u,ddR.ud,dRu4u,RdRj,u,.gRUu.,.Ru(RRRRRRRRF:Rk#0R0D8_FOoHRS;
Snu.,.Ru6u,R.Rc,u,.dR.u.,.Ru4u,R.Rj,u,4gRUu4SRSRRF:Rk#0R0D8_FOoHRS;
S(u4,4Runu,R4R6,u,4cRdu4,4Ru.u,R4R4,u,4jRRugRRRRRRRR:kRF00R#8F_DoRHO;S
SuRU,uR(,uRn,uR6,uRc,uRd,uR.,uR4,uSjSSRSRRF:Rk#0R0D8_FOoHRS
S2S;
CRM8ObFlFMMC0
;
RORRF0M#NRM0WRzvR:RRR0HMCsoCRR:=4R(;-I-RHE80RRFVFNsOd#kMHCoM8DRLFRO	l0kDHHbDCRs
RFROMN#0MW0R1RvRRRR:HCM0oRCs:4=RU-;R-HRI8R0EFFVRsdON#MHoCL8RD	FORDlk0DHbH
Cs
RRRO#FM00NMR)Z mR4(:0R#8F_Do_HOP0COF:sR=jR"jjjjjjjjjjjjjjjj"
;
SMOF#M0N0HRI8RNRRH:RMo0CC:sR=5R5N8IH0WE+z.v-2z/WvR2;RR--#MHoR0LHRRH#8bsFb
C8RORRF0M#NRM0ILH8R:RRR0HMCsoCRR:=5I5LHE80+vWz-/.2W2zv;-RR-HR#oLMRHH0R#sR8FCbb8R
RRMOF#M0N0bRIsR8RRH:RMo0CC:sR=HRI8+NRR8IHLR;R-I-RHE80RRFVb8sFk
O0SMOF#M0N0NRIsRsRRH:RMo0CC:sR=HRI8*NRR8IHLR;R-I-RHE80RRFVu0NsHRNDu8sFkRO0NNss$R
RRMOF#M0N0lRINRGRRH:RMo0CC:sR=$Rll5NGINH8,HRI8;L2
-
S-ERaCMRHb#k0RCNsRD#bHH0RMR0F4L(-HO0RE	kM#0,RERCMCENORkOEMH	R#HR#oCMRGM0C8
C8R0RR$RbCqb0$C#RHRsNsN5$RjFR0R8IHN2-4RRFV#_08DHFoOC_POs0F5WRR14v-RI8FMR0Fj
2;R0RR$RbCAb0$C#RHRsNsN5$RjFR0R8IHL2-4RRFV#_08DHFoOC_POs0F5WRR14v-RI8FMR0Fj
2;R-
S-ER0CDRCCMlC0F#RVER0CNRusN0HDkR1lFR)IN#Rs4CR(H-L0I#RH
8CR0RR$RbC1b0$C#RHRsNsN5$RjFR0RsIb82-4RRFV#_08DHFoOC_POs0F5WRRz4v-RI8FMR0Fj
2;
-S-RC0ERsbN0DHNRFbs80kO#sRNCnRd-0LH#HRI8RC
R$R0buCR0C$bRRH#NNss$jR5RR0FIsNs-R42F#VR0D8_FOoH_OPC05Fs.1*WvR-48MFI0jFR2
;
SR--aRECHkMb0H#RMRRNINH8RsNsNF$RVUR4-0LHRkOEM
	#So#HMRNDqsNsNR$RRRR:qb0$CS;
#MHoNADRNNss$RRRRA:R0C$b;S

-0-REuCRNHs0NuDRskF8ON0Rs$sNRRN#NNRIsNsRs$sNRRFVdLn-HO0RE	kM#R
RRo#HMRNDuVLkRRRRRRR:ub0$CR;
RHR#oDMNRFus8sqsN:$RR$u0b
C;SC
LoRHMRR--LODF	
#
SR--a#ECCIR0FsRbF#OC#RC#OMENo0CREPCRNNsHLRDCI0H8EMRHb#k0R0HMFHRVGRC8I0H8EMRHb#k03-
S-ERaCHRI8R0EF0VREHCRM0bk#sRNCMRHRvW1RFoskRb#VRFsLEF03]RRFPICCRs,0REC4LU-HS0
-o-RsbFk#NRCOOERFNM0H4MR(HRL0V#RsRFl0RECFosHHDMN,GRCO0CbRsVFRC0ER#lF0-
S-HR#oVMHHMON0sRoFRkb00ENR#NDFNRE#ER0CHR#oLMRHF0RVER0CsRFHMoHN
D3RsRRCx#HC:_NRFbsO#C#R25q
NSPsLHND CRGe0qNRDSR#:R0D8_FOoH_OPC05FsW-1v4FR8IFM0R;j2
CSLoRHMRR--bOsFCR##sHC#xNC_
RRRRVRRFHsR8HGRMRRj0WFR14v-RFDFbS
SSRHV58IHN2-4*vWz+GH8<HNI8R0E0MECR-R-RbOF$sRFHMoHNLDRH
0#SSSS qG0e5NDH28GRR:=q555INH8-*42W2zv+GH82S;
SDSC#SCRS-R-Ro#HMGRC08CM
SSSS0 GqDeN5GH82=R:Rqq5'VDC0
2;SCSSMH8RVS;
S8CMRFDFbR;R-H-R8SG
SsqNs5N$INH8-R42< =RGe0qN
D;S-S-RR8FMRF0#MHoR0CGCRM8pR1AoksFbS#
SsVFRGH8RRHMjFR0R8IHNR-.DbFF
SSSqsNsNH$58RG2<'=Rj&'RRWq5z5v*H+8G442-RI8FMR0FW*zvH28G;R
RRRRRCRM8DbFF;C
SMb8RsCFO#s#RCx#HC;_N
R
RR#sCH_xCLb:RsCFO#5#RAS2
PHNsNCLDR0 GADeNS:RRR8#0_oDFHPO_CFO0s15WvR-48MFI0jFR2R;
RCRLoRHMRR--bOsFCR##sHC#xLC_
RRRRVRRFHsR8HGRMRRj0WFR14v-RFDFbS
SSRHV58IHL2-4*vWz+GH8<HLI8R0E0MECR-R-RbOF$sRFHMoHNLDRH
0#SSSS AG0e5NDH28GRR:=A555ILH8-*42W2zv+GH82S;
SDSC#SCRS-R-Ro#HMGRC08CM
SSSS0 GADeN5GH82=R:RAA5'VDC0
2;SCSSMH8RVS;
S8CMRFDFbR;R-H-R8SG
SsANs5N$ILH8-R42< =RGe0AN
D;S-S-RR8FMRF0#MHoR0CGCRM8pR1AoksFbR#
RRRRRsVFRGH8RRHMjFR0R8IHLR-.DbFF
SSSAsNsNH$58RG2<'=Rj&'RRWA5z5v*H+8G442-RI8FMR0FW*zvH28G;S
SCRM8DbFF;-RR-8RHGR
RR8CMRFbsO#C#R#sCH_xCL
;
SR--oCCMsCN0RC0ERsuN0DHNRFus80kORsNsNL$R$kRlDb0HDM$HoER0CUR4-0LHRkOEMR	#FSV
-0-REHCRM0bk#FR0RsVFlnRd-0LHRsuN0DHNRFus80kO#R3R
o
SCkMlD:0NRsVFRRNGHjMRRR0FINH8-o4RCsMCN
0CSCSoMDlk0RL:VRFsLHGRMRRj0IFRH-8L4CRoMNCs0SC
S0SN0LsHkR0C\M3H0MCsNHD_MN#0MN0H0\C8RRFVl0kDG:GRRLDNCHDR#;R4
LSSCMoH
SSSl0kDG:GRRpvzaX4U4 U_vR
RRRRRb0FsRblNRR5
RRRRRRRRqR4(=q>RNNss$G5N2(542R,
RRRRRRRRqR4n=q>RNNss$G5N2n542R,
RRRRRRRRqR46=q>RNNss$G5N26542R,
RRRRRRRRqR4c=q>RNNss$G5N2c542R,
RRRRRRRRqR4d=q>RNNss$G5N2d542R,
RRRRRRRRqR4.=q>RNNss$G5N2.542R,
RRRRRRRRqR44=q>RNNss$G5N24542R,
RRRRRRRRqR4j=q>RNNss$G5N2j542R,
RRRRRRRRq=gR>NRqs$sN52NG5,g2
RRRRRRRRURqRR=>qsNsNN$5GU252R,
RRRRRRRRq=(R>NRqs$sN52NG5,(2
RRRRRRRRnRqRR=>qsNsNN$5Gn252R,
RRRRRRRRq=6R>NRqs$sN52NG5,62
RRRRRRRRcRqRR=>qsNsNN$5Gc252R,
RRRRRRRRq=dR>NRqs$sN52NG5,d2
RRRRRRRR.RqRR=>qsNsNN$5G.252R,
RRRRRRRRq=4R>NRqs$sN52NG5,42
RRRRRRRRjRqRR=>qsNsNN$5Gj252R,
RRRRRRRRAR4(=A>RNNss$G5L2(542R,
RRRRRRRRAR4n=A>RNNss$G5L2n542R,
RRRRRRRRAR46=A>RNNss$G5L26542R,
RRRRRRRRAR4c=A>RNNss$G5L2c542R,
RRRRRRRRAR4d=A>RNNss$G5L2d542R,
RRRRRRRRAR4.=A>RNNss$G5L2.542R,
RRRRRRRRAR44=A>RNNss$G5L24542R,
RRRRRRRRAR4j=A>RNNss$G5L2j542R,
RRRRRRRRA=gR>NRAs$sN52LG5,g2
RRRRRRRRURARR=>AsNsNL$5GU252R,
RRRRRRRRA=(R>NRAs$sN52LG5,(2
RRRRRRRRnRARR=>AsNsNL$5Gn252R,
RRRRRRRRA=6R>NRAs$sN52LG5,62
RRRRRRRRcRARR=>AsNsNL$5Gc252R,
RRRRRRRRA=dR>NRAs$sN52LG5,d2
RRRRRRRR.RARR=>AsNsNL$5G.252R,
RRRRRRRRA=4R>NRAs$sN52LG5,42
RRRRRRRRjRARR=>AsNsNL$5Gj252R,
RRRRRRRRuRd6=u>RL5kV5*NGILH82G+L265d2R,
RRRRRRRRuRdc=u>RL5kV5*NGILH82G+L2c5d2R,
RRRRRRRRuRdd=u>RL5kV5*NGILH82G+L2d5d2R,
RRRRRRRRuRd.=u>RL5kV5*NGILH82G+L2.5d2R,
RRRRRRRRuRd4=u>RL5kV5*NGILH82G+L245d2R,
RRRRRRRRuRdj=u>RL5kV5*NGILH82G+L2j5d2R,
RRRRRRRRuR.g=u>RL5kV5*NGILH82G+L2g5.2R,
RRRRRRRRuR.U=u>RL5kV5*NGILH82G+L2U5.2R,
RRRRRRRRuR.(=u>RL5kV5*NGILH82G+L2(5.2R,
RRRRRRRRuR.n=u>RL5kV5*NGILH82G+L2n5.2R,
RRRRRRRRuR.6=u>RL5kV5*NGILH82G+L265.2R,
RRRRRRRRuR.c=u>RL5kV5*NGILH82G+L2c5.2R,
RRRRRRRRuR.d=u>RL5kV5*NGILH82G+L2d5.2R,
RRRRRRRRuR..=u>RL5kV5*NGILH82G+L2.5.2R,
RRRRRRRRuR.4=u>RL5kV5*NGILH82G+L245.2R,
RRRRRRRRuR.j=u>RL5kV5*NGILH82G+L2j5.2R,
RRRRRRRRuR4g=u>RL5kV5*NGILH82G+L2g542R,
RRRRRRRRuR4U=u>RL5kV5*NGILH82G+L2U542R,
RRRRRRRRuR4(=u>RL5kV5*NGILH82G+L2(542R,
RRRRRRRRuR4n=u>RL5kV5*NGILH82G+L2n542R,
RRRRRRRRuR46=u>RL5kV5*NGILH82G+L26542R,
RRRRRRRRuR4c=u>RL5kV5*NGILH82G+L2c542R,
RRRRRRRRuR4d=u>RL5kV5*NGILH82G+L2d542R,
RRRRRRRRuR4.=u>RL5kV5*NGILH82G+L2.542R,
RRRRRRRRuR44=u>RL5kV5*NGILH82G+L24542R,
RRRRRRRRuR4j=u>RL5kV5*NGILH82G+L2j542R,
RRRRRRRRu=gR>LRuk5V5NIG*H28L+2LG5,g2
RRRRRRRRURuRR=>uVLk5G5N*8IHLL2+GU252R,
RRRRRRRRu=(R>LRuk5V5NIG*H28L+2LG5,(2
RRRRRRRRnRuRR=>uVLk5G5N*8IHLL2+Gn252R,
RRRRRRRRu=6R>LRuk5V5NIG*H28L+2LG5,62
RRRRRRRRcRuRR=>uVLk5G5N*8IHLL2+Gc252R,
RRRRRRRRu=dR>LRuk5V5NIG*H28L+2LG5,d2
RRRRRRRR.RuRR=>uVLk5G5N*8IHLL2+G.252R,
RRRRRRRRu=4R>LRuk5V5NIG*H28L+2LG5,42
RRRRRRRRjRuRR=>uVLk5G5N*8IHLL2+Gj252S
S2
;
SHSSVH_bb:L4RRHV5CMC8H_bbkCLV=#RRR42oCCMsCN0
SSSSVLkb:bHRsVFRHHRMRRj0.FR*vW1-o4RCsMCN
0CSSSSS0N0skHL0\CR3MsN	F\RVCRso:#RRLDNCHDR#;R4
SSSS0SN0LsHkR0C\C3Lo_HM0CsC\VRFRosC#RR:DCNLD#RHR
4;SSSSS0N0skHL0\CR3lsCF_PCMIF_N\sMRRFVs#CoRD:RNDLCRRH#4S;
SLSSCMoHRS
SSsSSC:o#RHRbbkCLVS
SSbSSFRs0l5Nb
SSSSSSSQ>R=RkuLVN55GH*I8+L2L5G2H
2,SSSSSmSSRR=>u8sFqNss$N55GH*I8+L2L5G2H;22
SSSS8CMRMoCC0sNCkRLVHbb;S
SS8CMRMoCC0sNCVRH_bbHL
4;SHSSVH_bb:LjRRHV5CMC8H_bbkCLV=#RRRj2oCCMsCN0
SSSSFus8sqsN5$5NIG*H28L+2LGRR<=uVLk5G5N*8IHLL2+G
2;SCSSMo8RCsMCNR0CHbV_HjbL;S
SCRM8oCCMsCN0RMoCl0kDLS;
CRM8oCCMsCN0RMoCl0kDN
;
SR--aCN	RC0ERsuN0DHNRFus80kORsNsNN$RML8Rk8HDRC0ER8N8C0sRs3CCRRRqsMkMHRMo#
klSR--HH#RMNH0DCHx80,RERCMFC0EsFRsIF#RVER0CNRbsN0HDsRbFO8k0sRNC8RN83C8
-S-RswFRNCGlCbD,VRHRHqR#UR6-0LH#HRI8NCRMA8RRRH#.Lc-HR0#ICH8,ER0CqMRR0VH#MRHRSc
-4-R(H-L0EROk#M	R8NMRVARHR0#H.MRR-4(LRH0OMEk	R#3RCaERsNsNI$RHRDDHDMOkR8Cc=*.
-S-RlURkHD0bCDHsV#RFHslMUoRR-dnLRH0u0NsHRNDu8sFk#O03aRREVCRkRDDb8sFkRO0IDHDRRLC
-S-R.c+=4nR(H-L0EROk#M	R8IHCR3RaREC)1kMkHlR#MRHHN0HDCHx8FR0:-
S-RRRRo1HM0 G,RRR1MHo ,G0RuRRu,544H2E,uRu544,2,DFR5uuj2,jERH,uju5,Dj2F-
S-ERaCFMR0sECRIsF#sRNCFRVs8lCR#LNCF8RMER0CHRI8R0EFqVRRRHM4L(-HO0RE	kM#MRN8-
S-ER0CHRI8R0EFAVRRRHM4L(-HO0RE	kM#R3RwRFs0RECClGNb:DC
-S-RCaER''qRFDFb4R5RR0FdS2
-R-RRHR1oGM 0R,RR5uu.2,4ERH,u.u5,D42Fu,Ru,54jH2E,uRu5j4,2,DFR#j'
-S-RRRRudu5,E42Hu,Ru,5d4F2D,uRu5j.,2,EHR5uu.2,jDRF,j,'#RRRRRjRR'S#
-R-RRHR1oGM 0R,RR5uud2,jERH,udu5,Dj2Fj,R'R#,RRRRR'Rj#R,RRRRRR#j'
-S-RCaER''ARFDFb4R5RR0F4S2
-R-RRHR1oGM 0R,RRo1HM0 G,RRR1MHo ,G0RuRRu,5j4H2E,uRu54j,2,DFR#j'
-S-RswFRlNRFRsC0sEFFEkoRbCGDNNM0MHF,CR#CER0CHResG0C-RQQAODF	kRvDb0HDsHC
-S-RC#bOHHVOHN0FRM3
R
RR8N8b8sF:sRbF#OC#uR5sqF8s$sN2S
SPHNsNCLDRM)k1RklR:RRR8#0_oDFHPO_CFO0sb5IsW8*z4v+RI8FMR0Fj:2R=FR50sEC#>R=R''j2R;
RRRRRsPNHDNLCkR1lI)FeRCO:0R#8F_Do_HOP0COFIs5b*s8W+zv4FR8IFM0R;j2
RRRRPRRNNsHLRDC1)klFRIRRRR:1b0$CR;
RRRRRsPNHDNLCHRN8RGRRRRR:MRH0CCosR;
RRRRRsPNHDNLCHRL8RGRRRRR:MRH0CCosR;
RRRRRsPNHDNLCRR[RRRRRRRR:MRH0CCosR;
RRRRRsPNHDNLCRR	RRRRRRRR:MRH0CCosS;
LHCoM-RR-sRbF#OC#8RN8Fbs8S
S-Q-RMHH0NxDHCER0CkRsMMMHokR#l)R5kkM1lR2
RRRRRsVFRRNGHjMRRR0FIGlN-D4RF
FbSLSSHR8G:N=RGS;
SRS[R:RR=*R.N
G;S	SSRRRR:[=RR4+R;S
SSRHVN>GRR8IHNR-4FLsRHR8G>HRI84L-RC0EMS
SSVSHR<[RRsIb8ER0CRMRS-SR-HR#oCMRGM0C8S
SS1SSkFl)I25[RR:=5EF0CRs#=u>RsqF8s$sN5o1HMFADOI	5H,8NILH8,2j25W.*1.v-2
2;SSSSCRM8H
V;SSSSH	VRRI<RbRs80MECRSRSRR--#MHoR0CGC
M8SSSSSl1k)5FI	:2R=FR50sEC#>R=RFus8sqsN1$5HAoMD	FO58IHNH,I8jL,2.25*vW1-2.2;S
SSMSC8VRH;S
SS#CDCS
SSkS1lI)F5R[2:u=RsqF8s$sN5*NGILH8+8LHGR25RvWz-84RF0IMFRRRj
2;RRRRRRRRRRRRH	VRRI<RbRs80MEC
SSSSkS1lI)F5R	2:u=RsqF8s$sN5*NGILH8+8LHG.25*vWz-84RF0IMFzRWv
2;SSSSCRM8H
V;SCSSMH8RVS;
S-S-RMOFP0CsRC0ERsNsNF$RVEROk#M	R0HMFMRNRsNsNF$RVHRL0S#
SFSVsLRHGMRHR0jRFbRIs48-RFDFbS
SSFSVsGRDRRHMjFR0RvWz-D4RF
FbSSSSSM)k15klH*LGW+zvDRG2:1=RkFl)IL5HGD25G
2;SSSSCRM8DbFF;-RR-GRD
SSSCRM8DbFF;-RR-LRHGS
SSR--H0MHHHNDx0CRE#CRHRoML#H0
SSS)1kMkIl5b*s8W+zv4FR8IFM0RsIb8z*Wv:2R=FR50sEC#>R=RFus8sqsN1$5HAoMD	FO58IHNH,I8jL,2.25*vW1-2.2;S
SCRM8DbFF;-RR-GRN
-SS-FRpFFbRMER0CRRqHCM8GS
SVRFsHR8GH4MRRR0FINH8-D4RF
FbRRRRRRRRRsVFRRNGHjMRRR0FIGlN-D4RF
FbSSSSLGH8RR:=N-GRRGH8;S
SSRS[R:RR=GRNRL+RH;8G
SSSSR	RR=R:R+[RR
4;SSSSHNVRGRR>INH8-F4RsHRL8>GRR8IHLR-40MEC
RRRRRRRRRRRRRRRH[VRRI<RbRs80MECRSRSRR--#MHoR0CGC
M8SSSSSkS1lI)F5R[2:5=RFC0Es=#R>uR5sqF8s$sN5o1HMFADOI	5H,8NILH8,GH82.25*vW1-2.22S;
SSSSCRM8H
V;SSSSSRHV	RR<I8bsRC0EMSRRS-R-Ro#HMGRC08CM
SSSS1SSkFl)I25	RR:=5EF0CRs#=5>Ru8sFqNss$H51oDMAF5O	INH8,8IHL8,HG522.1*Wv2-.2
2;SSSSS8CMR;HV
SSSS#CDHLVRHR8G<RRj0MEC
SSSSVSHR<[RR0jRERCMRSSSRR--Nk8[#00REHCRMH8OCl#RFD8kFlRINSG
SSSSS:[R=RR[+*R.IGlN;R
RRRRRRRRRRRRRR8CMR;HV
RRRRRRRRRRRRRRRH	VRRj<RRC0EMS
SSSSS	=R:R+	RRI.*l;NG
SSSSMSC8VRH;S
SSHSSVRR[<GRNRC0EMS
SSSSS1)klF[I52=R:R)Z m;4(
SSSSDSC#RHV[RR<I8bsRC0EMSRRS-R-Ro#HMGRC08CM
SSSS1SSkFl)I25[RR:=5EF0CRs#=5>Ru8sFqNss$H51oDMAF5O	INH8,8IHL8,HG522.1*Wv2-.2
2;SSSSS8CMR;HV
SSSS-S-REF0CHsI#RC,0RECHCM8G#RHR0MFRRHM0REC1)klFRI,8MFRFH0EMSo
SSSSH	VRRR<=N0GRE
CMSSSSSkS1lI)F5R	2:Z=R 4)m(R;
RRRRRRRRRRRRRDRC#RHV	RR<I8bsRC0EMSRRS-R-Ro#HMGRC08CM
SSSS1SSkFl)I25	RR:=5EF0CRs#=5>Ru8sFqNss$H51oDMAF5O	INH8,8IHL8,HG522.1*Wv2-.2
2;SSSSSR--FC0Es#IHC0,REHCRMG8CRRH#MRF0H0MRE1CRkFl)I8,RFFRM0MEHoS
SSCSSMH8RVS;
SCSSDR#CRSSSSSSSRR--MlFsNbDRskF8O00RC
slSSSSSl1k)5FI[:2R=sRuFs8qs5N$NIG*H+8LLGH82R5RW-zv4FR8IFM0RjRR2S;
SSSSH	VRRI<RbRs80MEC
SSSS1SSkFl)I25	RR:=u8sFqNss$G5N*8IHLH+L85G2.z*WvR-48MFI0WFRz;v2
SSSSMSC8VRH;S
SSMSC8VRH;S
SS8CMRFDFbR;R-N-RGS
SSR--OPFMCRs00RECNNss$VRFRkOEMR	#HFM0RRNMNNss$VRFR0LH#R
RRRRRRVRRFHsRLHGRMRRj0IFRb-s84FRDFSb
SVSSFDsRGMRHR0jRFzRWvR-4DbFF
SSSSkS1lI)Fe5COH*LGW+zvDRG2:1=RkFl)IL5HGD25G
2;SSSSCRM8DbFF;-RR-GRD
SSSCRM8DbFF;-RR-LRHGS
SSR--1RC00REC#MHoR0LH#FRVsER0Hs#RFRI
RRRRRRRR1)klFCIeOb5IsW8*z4v+RI8FMR0FI8bs*vWz2=R:RFR50sEC#>R=RFus8sqsN1$5HAoMD	FO58IHNH,I8HL,82G25W.*1.v-2
2;S-SS-8Rq8ER0CFRsIkR[#O0Rs0CNC08RFER0CkRsMMMHokR#lR
RRRRRR)RRkkM1l=R:RM)k1Rkl+kR1lI)Fe;CO
CSSMD8RF;FbR-R-RGH8
-SS-FRpFFbRMER0CRRAHCM8GS
SVRFsHRxGH4MRRR0FILH8-D4RF
FbRRRRRRRRRsVFRRLGHjMRRR0FIGlN-D4RF
FbSSSSNGH8RR:=L-GRRGHx;S
SSRS[R:RR=HRN8+GRR;LG
SSSSR	RR=R:R+[RR
4;SSSSHLVRGRR>ILH8-F4RsHRN8>GRR8IHNR-40MEC
RRRRRRRRRRRRRRRH[VRRI<RbRs80MECRSRSRR--#MHoR0CGC
M8SSSSSkS1lI)F5R[2:5=RFC0Es=#R>uR5sqF8s$sN5o1HMFADOI	5H,8NILH8,x-HG522.1*Wv2-.2
2;SSSSS8CMR;HV
SSSSVSHR<	RRsIb8ER0CRMRS-SR-HR#oCMRGM0C8S
SSSSS1)klF	I52=R:R05FE#CsRR=>5Fus8sqsN1$5HAoMD	FO58IHNH,I8-L,H2xG2*5.W-1v.222;S
SSCSSMH8RVS;
SCSSDV#HR8NHGRR<jER0CSM
SSSSH[VRRj<RRC0EMSRRS-SR-8RN[0k#RC0ER8HMO#HCR8lFkRDFIGlN
SSSS[SSRR:=[RR+.l*IN
G;SSSSS8CMR;HV
SSSSVSHR<	RR0jRE
CMSSSSSRS	:	=RR.+R*NIlGS;
SSSSCRM8H
V;SSSSSRHV[RR<L0GRE
CMSSSSSkS1lI)F5R[2:Z=R 4)m(R;
RRRRRRRRRRRRRDRC#RHV[RR<I8bsRC0EMSRRS-R-Ro#HMGRC08CM
SSSS1SSkFl)I25[RR:=5EF0CRs#=5>Ru8sFqNss$H51oDMAF5O	INH8,8IHLH,-x2G25W.*1.v-2;22
SSSSMSC8VRH;S
SSHSSVRR	<L=RGER0CSM
SSSSSl1k)5FI	:2R= RZ)(m4;R
RRRRRRRRRRRRRR#CDH	VRRI<RbRs80MECRSRSRR--#MHoR0CGC
M8SSSSSkS1lI)F5R	2:5=RFC0Es=#R>uR5sqF8s$sN5o1HMFADOI	5H,8NILH8,x-HG522.1*Wv2-.2
2;SSSSS8CMR;HV
SSSS#CDCS
SS1SSkFl)I25[RR:=u8sFqNss$H5N8IG*H+8LL5G2RzRWvR-48MFI0RFRR;j2
SSSSVSHR<	RRsIb8ER0CSM
SSSSSl1k)5FI	:2R=sRuFs8qs5N$NGH8*8IHLG+L2*5.W-zv4FR8IFM0RvWz2S;
SSSSCRM8H
V;SSSSCRM8H
V;SCSSMD8RF;FbR-R-R
LGS-SS-FROMsPC0ER0CsRNsRN$FOVRE	kM#MRH0NFRMsRNsRN$FLVRH
0#RRRRRRRRRsVFRGHNRRHMjFR0RsIb8R-4DbFF
SSSSsVFRRDGHjMRRR0FW-zv4FRDFSb
SSSS1)klFCIeON5HGz*WvG+D2=R:Rl1k)5FIH2NG52DG;S
SSMSC8FRDFRb;RR--DSG
SMSC8FRDFRb;RR--H
NGS-SS-CR10ER0CHR#oLMRHR0#VRFs0#EHRIsF
RRRRRRRRkR1lI)Fe5COI8bs*vWz+84RF0IMFbRIsW8*zRv2:R=R5EF0CRs#=u>RsqF8s$sN5o1HMFADOI	5H,8NILH8,x-HG522.1*Wv2-.2S;
S-S-R8q8RC0ERIsFR#[k0sROCCN08FR0RC0ERMskMoHMRl#k
RRRRRRRRkR)Ml1kRR:=)1kMk+lRRl1k)eFIC
O;SMSC8FRDFRb;RR--H
xGRRRRR)Rum<7R=kR)Ml1k5HNI8+0EL8IH04E-RI8FMR0Fj
2;S8CMRFbsO#C#R8N8b8sF;C

ML8RD	FO#
;
-*-R*************************************************************R**R
---
-R- -RM00H$CR7OsDNNF0HMFRVsHR#o8MCRDlk0DHbH
Cs-
-R-a-RERH#H0#RElCRNRHMCHM00V$RF0sRE#CRHCoM8kRlDb0HDsHC3aRRE0CRINFRsHOE00COk#sC
R--8HCVMRC8LFCDI#RkCER0CMRC0HH0CN#RLCFP,MRN8kRl#L0RCNRD#H0RMER0HV#RH3DCRERaC-
-RF0IRONsECH0Os0kCN#Rs0CREDCRFOoHRsPC#MHFR8NMRC0ERFLDOP	RCHs#F
M3-
-R-*-R*************************************************************R**R
--
LDHs$NsRCHCCk;
#HCRC3CC#_08DHFoO4_4nNc3D
D;kR#CHCCC38#0_oDFHNO_sEH03DND;#
kCCRHC#C30D8_FOoH_#kMHCoM8D3ND
;
DsHLNRs$FNsOdk;
#FCRsdON3OFsNlOFbD3ND
;
DsHLNRs$#b$MD$HV;#
kC$R#MHbDVN$30H0sLCk0#D3ND
;
CHM001$RvazpR
H#RRRRoCCMs5HO
RRRRRRRI0H8E:RRR0HMCsoCRR:=.
c;RRRRRNRRI0H8ERR:HCM0oRCs:4=R.R;
RRRRRIRLHE80RH:RMo0CC:sR=.R4
RSS2R;
RbRRF5s0
RSSqRRRRH:RM0R#8F_Do_HOP0COFNs5I0H8E4R-RI8FMR0Fj
2;SASRRRRR:MRHR8#0_oDFHPO_CFO0sI5LHE80RR-48MFI0jFR2S;
S)Rum:7RR0FkR8#0_oDFHPO_CFO0sH5I8R0E-84RF0IMF2Rj
RRRRRRR2R;
R0RN0LsHkR0C\N3sMR	\:MRH0CCosR;
R0RN0LsHkR0C\F3l8CkD\RR:#H0sM
o;RNRR0H0sLCk0Rb\3Fl8C\RR:HCM0o;Cs
RRRNs00H0LkC3R\bCF8l#Lk\RR:#H0sM
o;RNRR0H0sLCk0RC\3M08_s\CCRH:RMo0CC
s;RNRR0H0sLCk0RL\3CMoH_C0sC:\RR0HMCsoC;R
RR0N0skHL0\CR3lsCF_PCMIF_N\sMRH:RMo0CC
s;CRM81pvza
;
-*-R*************************************************************R**R
---
-R-D-RFOoHRONsECH0Os0kCV#RFFsRsdON
R--
R--****************************************************************R-R-
s
NO0EHCkO0sDCRFOoHRRFV1pvza#RH
R
RRMVkOF0HMNROD8IH0REL5MOF#M0N0NRI,LRIRH:RMo0CCRs2skC0sHMRMo0CCHsR#R
RRRRRPHNsNCLDRMsO0RR:HCM0o;Cs
RRRLHCoMR
RRRRRH5VRI<LR=NRI2ER0CRM
RRRRRRRRs0OMRR:=I;LR
RRRRCRRDR#C
RRRRRRRRORsM:0R=NRIRR;
RRRRR8CMR;HV
RRRRsRRCs0kMORsM
0;RCRRMO8RNHDI8L0E;R

RkRVMHO0FOMRNHDI8N0ERF5OMN#0MI0RNI,RLRR:HCM0o2CsR0sCkRsMHCM0oRCsHR#
RRRRRsPNHDNLCORsM:0RR0HMCsoC;R
RRoLCHRM
RRRRRRHV5RIL<I=RN02RE
CMRRRRRRRRRMsO0=R:RRIN;R
RRRRRCCD#RR
RRRRRRsRRORM0:I=RL
R;RRRRRMRC8VRH;R
RRRRRskC0ssMRO;M0
RRRCRM8OINDHE80N
;
RORRF0M#NRM0I0H8E:NRR0HMCsoCRR:=OINDHE80NI5NHE80,IRLHE802R;
RFROMN#0MI0RHE80LRR:HCM0oRCs:O=RNHDI8L0E5HNI8,0ERHLI820E;R

RFROlMbFCRM0#DlNDDvk0R
RRRRRoCCMs5HO
RRRRRRRRIRNHE80RH:RMo0CC;sR
RRRRRRRRIRLHE80RH:RMo0CC;sR
RRRRRRRRHRI8R0ERH:RMo0CCRs
RRRRR
2;RRRRRFRbs50R
RRRRRRRRRRqR:RRRRHMR8#0_oDFHPO_CFO0sI5NHE80-84RF0IMF2Rj;R
RRRRRRARRRRRR:MRHR0R#8F_Do_HOP0COFLs5I0H8ER-48MFI0jFR2R;
RRRRRRRRu7)mRF:Rk#0R0D8_FOoH_OPC05FsR8IH04E-RI8FMR0FjR2
RRRRR
2;RCRRMO8RFFlbM0CM;R

RHR#oDMNRNN_kRGR:0R#8F_Do_HOP0COFIs5HE80NR-48MFI0jFR2R;R
RRR#MHoNLDR_GNkRRR:#_08DHFoOC_POs0F58IH0-EL4FR8IFM0R;j2RR
RRo#HMRND)kC#D:0RR8#0_oDFHPO_CFO0sI5RHE80-84RF0IMF2Rj;C
Lo
HMR-RR-CRp0R'##bIN
RRRQIw_Nk_#bL_I:VRHRI5NHE80RR>=L8IH0RE2oCCMsCN0
RRRRNRR_GNkRR<=NR;
RRRRRNL_k<GR=;RL
RRRCRM8oCCMsCN0R_QwI#N_kIb_L
;
RQRRwL_I_b#k_:INRRHV5HLI8R0E>IRNHE802CRoMNCs0RC
RRRRRNN_k<GR=;RL
RRRRLRR_GNkRR<=NR;
RMRC8CRoMNCs0QCRwL_I_b#k_;IN
H
SV4_I:VRHRH5I8L0ER4=R2CRoMNCs0SC
So#HMRNDObFlDCClMR0,0OIFFRlb:0R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj;S
SLHCoMS
SV_FsDbFF:FRVsRRHHjMRRR0FI0H8E4N-RMoCC0sNCS
SSlOFblDCC5M0H<2R=FRM0_RNN5kGHR2;
CSSMo8RCsMCNR0CV_FsDbFF;S
SSlOFblDCC5M0I0H8E2-4RR<=MRF0Nk_NGH5I8N0E-;42
SSS0OIFFRlb<O=RFDlbCMlC0RR+';4'
sSSCD#k0=R<RhBmea_17m_pt_QBea Bmj)5,HRI8N0E+8IH02ELRCIEMLR5_GNk5Rj2=jR''S2
SCSSDR#C0OIFF;lb

SSS)Sum<7R=CRs#0kD58IH04E-RI8FMR0Fj
2;S8CMRMoCC0sNCVRH_;I4
R
RR_HVIRj:H5VRI0H8E=LRRR.2oCCMsCN0
RRRR#RRHNoMDFROlCbDl0CM,IR0FlOFbRR:#_08DHFoOC_POs0F58IH0-EN4FR8IFM0R;j2
RRRLHCoMR
RRRRRV_FsDbFF:FRVsRRHHjMRRR0FI0H8E4N-RMoCC0sNCR
RRRRRRORRFDlbCMlC025HRR<=MRF0Nk_NG25H;RR
RRRRR8CMRMoCC0sNCFRVsF_DF
b;RRRRRIR0FlOFb=R<RlOFblDCCRM0+4R''
;
RRRRRCR)#0kDRR<=Bemh_71a_tpmQeB_ mBa),5jRHNI8+0EL8IH0RE2IMECR_5LN5kGj=2RR''j2R
RRRRRRRRRRDRC#0CRIFFOlIb5HE80L2-4R0&RIFFOlIb5HE80L2-4R0&RIFFOlIbRERCM5NL_k4G52RR='24'
RRRRRRRRRRRR#CDC_RNN5kGI0H8E4L-2RR&Nk_NGH5I8L0E-R42&_RNNRkG;R

RRRRRmu)7=R<R#)Ck5D0I0H8ER-48MFI0jFR2R;
RMRC8CRoMNCs0HCRVj_I;R

RVRH_4.I:VRHRH5I8L0ER.>R2CRoMNCs0RC
RRRRRDlk0R4:RN#lDzDvpRa
RRRRRRRRRoRRCsMCHlORN5bR
RRRRRRRRRRRRRRRRRRRRIRNHE80RR=>I0H8E
N,RRRRRRRRRRRRRRRRRRRRRHLI8R0E=I>RHE80LR,
RRRRRRRRRRRRRRRRRRRRI0H8E=RR>HRI8
0ERRRRRRRRRRRR2R
RRRRRRRRRRFRbsl0RN5bR
RRRRRRRRRRRRRRRRRRRRRRq=N>R_GNk,R
RRRRRRRRRRRRRRRRRRARRRR=>Lk_NGR,
RRRRRRRRRRRRRRRRRRRRu7)mRR=>u7)m
RRRRRRRRRRRR
2;RCRRMo8RCsMCNR0CH.V_I
4;
8CMRoDFH
O;
R--****************************************************************R-R-
R--
R--LODF	k_lDN0RsHOE00COk#sCRsVFROFsN-d
--R
-*R**************************************************************R*R-
-
NEsOHO0C0CksRFLDOl	_kRD0F1VRvazpR
H#
-S-RsbkbCF#:CRs0Mks#ER0CCRMIHRI8R0ELCN#8MRFROCGCR##L#H0RHLCMboRsCC#MR0
RkRVMHO0FbMRNW##HE80RR5
RRRRRMOF#M0N0FRl88IH0:ERR0HMCsoC;R
RRRRRO#FM00NMR8FDW0H8ERR:HCM0o2Cs
sSSCs0kMMRH0CCos#RH
CSLoRHMRR--b#N#W0H8ER
RRRRRHlVRFH8I8R0E>RR.0MECR-RS-FRl#00RNR	C0#EHRNLsM
OESsSSCs0kMDRF88WH0
E;SDSC#RHVlIF8HE80R.=RRC0EMS
SS0sCkRsMFWD8HE80-
.;SDSC#RHVlIF8HE80R4=RRC0EMS
SS0sCkRsMFWD8HE80-
4;SDSC#RHVlIF8HE80Rj=RRC0EMS
SS0sCkRsMFWD8HE80;S
SCCD#RSRSSSSS-0-RERH#H##RksbCVFDkkS#
SCSs0MksR8FDW0H8ES;
S8CMR;HV
MSC8NRb#H#W8;0E
-
S-CRs0MksRH4RVNROMHRbbHCDM0CRElCRkHD0bCDHsV
Sk0MOHRFMM8CC__0FbCHbDCHM5HNI8,0ERHLI8R0E:MRH0CCoss2RCs0kMMRH0CCos#RH
CSLo
HMSVSHRN55I0H8ERR>4R(2NRM85HLI8R0E>(R4202RE
CMSsSSCs0kM;R4
CSSMH8RVS;
S0sCkRsMjS;
CRM8M8CC__0FbCHbDCHM;R

R-R-RMVH8ER0ClR#NCDDsHRI8R0E58IH0FERsIRNHE802R
RRMVkOF0HMMRHVH5I8,0ERHNI8R0E:MRH0CCoss2RCs0kMMRH0CCos#RH
RRRLHCoMR
RRRRRH5VRI0H8ERR<N8IH0RE20MEC
RRRRRRRRCRs0MksR8IH0
E;RRRRRDRC#RC
RRRRRRRRskC0sNMRI0H8ER;
RRRRR8CMR;HV
RRRCRM8H;MV
R
RRMVkOF0HMHR#o8MCl5F8I0H8ERR:HCM0o2CsR0sCkRsMHCM0oRCsHS#
LHCoMSRRSSSSSSSS
RRRRHRRVHRI8<0E40gRESCMRR--4HgR#zRWvRR+.S
SS0sCkRsMI0H8ER;RRR--4H(R#zRWv4,R6#RHRvWz-R.
RRRRR#CDCS
SS0sCkRsM58IH04E-25-55H5I8+0E4/624-(2442*(
2;SRSRCRM8HRV;RC
SM#8RHCoM88lF;R

RFROMN#0MW0RzRvRRH:RMo0CC:sR=(R4;SRRRR--I0H8EVRFR#kMHCoM8kRlDb0HDsHC
R
RRMOF#M0N0IRNHR8C:MRH0CCos=R:RVHM58IH0RE,N8IH0;E2
FSOMN#0ML0RICH8RH:RMo0CC:sR=MRHVH5I8,0ERHLI820E;R

RFROMN#0MN0RlRF8RH:RMo0CC:sR=HR#o8MCl5F8N8IHC
2;RORRF0M#NRM0L8lFRRR:HCM0oRCs:#=RHCoM88lF5HLI8;C2
R
RRMOF#M0N0IRNH:8RR0HMCsoCRR:=b#N#W0H8El5NFR8,N8IHC
2;RORRF0M#NRM0L8IHRH:RMo0CC:sR=NRb#H#W850EL8lF,IRLH28C;S

O#FM00NMRCMC8H_bbkCLV:#RR0HMCsoCRR:=M8CC__0FbCHbDCHM5HNI8,0ERHLI820E;S

#MHoNCDR4RRRR:RRR8#0_oDFHPO_CFO0sR548MFI0jFR2S;
#MHoNCDR.RRRR:RRR8#0_oDFHPO_CFO0sR548MFI0jFR2S;
SSSSRRR
RHR#oDMNRsq0HRlRR#:R0D8_FOoH_OPC05FsN8IHCR-48MFI0jFR2R;
RHR#oDMNRsA0HRlRR#:R0D8_FOoH_OPC05FsL8IHCR-48MFI0jFR2
;
R#RRHNoMDbRqsCHlRRR:#_08DHFoOC_POs0F5HNI8R-48MFI0jFR2R;
RHR#oDMNRsAbHRlCR#:R0D8_FOoH_OPC05FsL8IH-84RF0IMF2Rj;R
RRo#HMRND1sEF0RuR:0R#8F_Do_HOP0COFNs5I+H8L8IH-84RF0IMF2RjRR:=5EF0CRs#='>Rj;'2
R
RRo#HMRND)kC#DR04:0R#8F_Do_HOP0COFNs5ICH8+HLI84C-RI8FMR0Fj
2;R#RRHNoMDCR)#0kDGRR:#_08DHFoOC_POs0F5HNI8LC+ICH8-84RF0IMF2Rj;R
RRo#HMRND)kC#DR0N:0R#8F_Do_HOP0COFNs5ICH8+HLI84C-RI8FMR0Fj
2;R#RRHNoMDCR)#0kDLRR:#_08DHFoOC_POs0F5HNI8LC+ICH8-84RF0IMF2Rj;R
RRo#HMRND)kC#DR0C:0R#8F_Do_HOP0COFNs5ICH8+HLI84C-RI8FMR0Fj
2;
RRR#MHoNuDRs4F8,sRuF_84N,kGRFus8s4_CR#RR#:R0D8_FOoH_OPC05FsN8IHCI+LH-8C4FR8IFM0R;j2
RRR#MHoNuDRs.F8R:RRR8#0_oDFHPO_CFO0sH5I8-0E4FR8IFM0R;j2
O
SFFlbM0CMRAe.pimB
oSSCsMCH5OR
SSSN8IH0:ERR0HMCsoCRR:=N8IH;S
SSHLI8R0E:MRH0CCos=R:RHLI8S;
SCSMCb8_HLbCkRV#:MRH0CCos
2;SFSbs50R
SSSqRRRRH:RM#RR0D8_FOoH_OPC05FsN8IH-84RF0IMF2Rj;S
SSRARRRR:HRMR#_08DHFoOC_POs0F5HLI8R-48MFI0jFR2S;
S)Sum:7RR0FkR8#0_oDFHPO_CFO0sI5NHL8+I-H84FR8IFM0R2j2;C
SMO8RFFlbM0CM;L

CMoHR-R-RFLDOl	_k
D0
-S-RsbkbCF#:NR0	OCRNRsCF0VRE4CRR8NMRL.-HO0RN##C
-S-Rb0$CRRR:FROlMLHNF0HM
NDSR--HkMb0:#RRRq,A-
S-kRF00bk#u:R)
m7SR--0lsHRC0ERbHMkR0#0LFRCFRMR8IHC0sRERNM0RECFbk0kS0
HbV_H4bC:VRHRC5MCb8_HLbCkRV#=2R4RMoCC0sNCS
S0lsHHq0_:FRVsRRHHjMRRR0FN8IHCR-4oCCMsCN0
SSSNs00H0LkC3R\s	NM\VRFRosC#:qRRLDNCHDR#;Rj
SSSNs00H0LkC3R\bCF8lF\RVCRsoR#q:NRDLRCDHH#R;S
SS0N0skHL0\CR38bFCklL#F\RVCRsoR#q:NRDLRCDH"#Rq
";SNSS0H0sLCk0Rl\3FD8kCF\RVCRsoR#q:NRDLRCDH"#R1pvza
";SNSS0H0sLCk0Rs\3CPlFCF_M_sINMF\RVCRsoR#q:NRDLRCDH4#R;S
SLHCoMS
SSosC#Rq:RbbHCVLk
SSSb0FsRblN5S
SSQSSRR=>q25H,S
SSmSSRR=>qH0sl25H2S;
S8CMRMoCC0sNCsR0H0lH_
q;
0SSsHHl0RA:VRFsHMRHR0jRFIRLH-8C4CRoMNCs0SC
S0SN0LsHkR0C\N3sMR	\FsVRCAo#RD:RNDLCRRH#jS;
S0SN0LsHkR0C\F3b8\ClRRFVs#CoARR:DCNLD#RHR
H;SNSS0H0sLCk0Rb\3Fl8CL\k#RRFVs#CoARR:DCNLD#RHR""A;S
SS0N0skHL0\CR38lFk\DCRRFVs#CoARR:DCNLD#RHRv"1z"pa;S
SS0N0skHL0\CR3lsCF_PCMIF_N\sMRRFVs#CoARR:DCNLD#RHR
4;SCSLo
HMSsSSCAo#:bRRHLbCkSV
SbSSFRs0l5Nb
SSSSQSSRR=>A25H,S
SSSSSm>R=RsA0HHl52
2;SMSC8CRoMNCs00CRsHHl0
A;S8CMRMoCC0sNCVRH_bbHC
4;S_HVbCHbjH:RVMR5C_C8bCHbL#kVRj=R2CRoMNCs0SC
Ssq0H<lR=5RqN8IHCR-48MFI0jFR2S;
SsA0H<lR=5RAL8IHCR-48MFI0jFR2S;
CRM8oCCMsCN0R_HVbCHbj
;
SR--sFClP0CRECCRGN0sR0LH#0RNRC0ERAp1R8CM
RRRbMskC:H0RFbsO#C#R05qs,HlRsA0H
l2SoLCHRMR-b-RsCFO#b#RsCkMHS0
SRHVN8lFR4=RRC0EMS
SSRC4<'=Rj&'RRsq0Hjl52S;
SbSqsCHlRR<=qH0slI5NH-8C4FR8IFM0R;42
CSSDV#HRFNl8RR=.ER0CRM
RRRRRRRRC<4R=0Rqs5Hl4FR8IFM0R;j2
SSSqHbsl<CR=0Rqs5HlN8IHCR-48MFI0.FR2R;
RRRRR#CDCS
SSRC4<'=Rj&'RR''j;S
SSsqbHRlC<q=R0lsH;S
SCRM8H
V;
HSSVlRLF=8RR04RE
CMSCSS.=R<R''jRA&R0lsH5;j2
SSSAHbsl<CR=0RAs5HlL8IHCR-48MFI04FR2S;
S#CDHLVRlRF8=RR.0MEC
RRRRRRRR.RCRR<=AH0slR548MFI0jFR2S;
SbSAsCHlRR<=AH0slI5LH-8C4FR8IFM0R;.2
RRRRCRRD
#CSCSS.=R<R''jR'&Rj
';SASSblsHC=R<RsA0H
l;SMSC8VRH;C
SMb8RsCFO#b#RsCkMH
0;
-S-RDvk0DHb$$RLRC0ER0CGsLNRHR0#HIVRCNREPFCRMFCRsIR0FGRC0RsNL#H0RRFVqH
SV4_N:VRHRl5NF48=2CRoMNCs0SC
S_HVNj4L:VRHRl5LF<8R=RRjFLsRlRF8>2R.RMoCC0sNCS
SS#)CkND0RR<=Bemh_71a_tpmQeB_ mBa),5jRHNI8LC+ICH82ERIC5MRCj452RR='2j'RS
SSSSSRDRC#1CRXAa5blsHCN,RICH8+HLI8;C2
RRRRCRRMo8RCsMCNR0CHNV_4;Lj
HSSV4_NLR4:H5VRL8lFR4=R2CRoMNCs0SC
SCS)#0kDN=R<RhBmea_17m_pt_QBea Bmj)5,IRNH+8CL8IHCI2RERCM55C4j=2RR''j2SR
SSSSSCRRDR#C15XaAHbsl&CRR''j,IRNH+8CL8IHC
2;RRRRRMRC8CRoMNCs0HCRV4_NL
4;SVSH_LN4.H:RVLR5lRF8=2R.RMoCC0sNCS
SS#)CkND0RR<=Bemh_71a_tpmQeB_ mBa),5jRHNI8LC+ICH82ERIC5MRCj452RR='2j'RS
SSSSSRDRC#1CRXAa5blsHCRR&'Rj'&jR''N,RICH8+HLI8;C2
RRRRCRRMo8RCsMCNR0CHNV_4;L.
MSC8CRoMNCs0HCRV4_N;H
SV.NM:VRHRl5NF.8=R8NMRHNI8>0E.o2RCsMCNR0CRR--zQh1t7h 
RRRR#RRHNoMDFRM1VEH0#,RE0HVCR8,NC888RR:#_08DHFoOC_POs0F5HNI8LC+ICH8-84RF0IMF2Rj;L
SCMoH
HSSV.NMLRj:H5VRL8lFRR<=jsRFRFLl8RR>.o2RCsMCN
0CRSRRS1MFE0HVRR<=15XaAHbslRC,N8IHCI+LH28C;R
RRRRRCRM8oCCMsCN0RNHVMj.L;S
SHMVN.:L4RRHV5FLl8RR=4o2RCsMCN
0CRSRRS1MFE0HVRR<=15XaAHbsl&CRR''j,IRNH+8CL8IHC
2;RRRRRMRC8CRoMNCs0HCRV.NML
4;SVSHNLM..H:RVLR5lRF8=2R.RMoCC0sNCR
RRMSSFH1EV<0R=XR1ab5AsCHlR'&Rj&'RR''j,IRNH+8CL8IHC
2;RRRRRMRC8CRoMNCs0HCRV.NML
.;SES#HCV08=R<R1MFE0HV5HNI8LC+ICH8-8.RF0IMF2RjR'&Rj
';RRRRR8RN8RC8R=R<R1MFE0HVR#+RE0HVC
8;SCS)#0kDN=R<RhBmea_17m_pt_QBea Bmj)5,HNI8LC+ICH82ERIC5MRC=4RRj"j"S2
SSSSRDRC#MCRFH1EVI0RERCM5RC4=jR"4
"2SSSSSCRRDR#C#VEH0RC8IMECR45CR"=R42j"
SSSSRSRCCD#R8N8CS8;RR--R45CR"=R424"
MSC8CRoMNCs0HCRV.NM;H
SV._N:VRHRl5NF.8=R8NMRHNI8=0E.o2RCsMCNR0CRR--1hQt S7
So#HMRNDMEF1H,V0RlOFblDCC,M0RF0IObFlR#:R0D8_FOoH_OPC05FsN8IHCI+LH-8C4FR8IFM0R;j2
CSLo
HMSVSH_LN.jH:RVLR5lRF8<j=RRRFsL8lFR.>R2CRoMNCs0RC
RSRRS1MFE0HVRR<=15XaAHbslRC,N8IHCI+LH28C;R
RRRRRCRM8oCCMsCN0R_HVNj.L;S
SHNV_.:L4RRHV5FLl8RR=4o2RCsMCN
0CRSRRS1MFE0HVRR<=15XaAHbsl&CRR''j,IRNH+8CL8IHC
2;RRRRRMRC8CRoMNCs0HCRV._NL
4;SVSH_LN..H:RVLR5lRF8=2R.RMoCC0sNCR
RRMSSFH1EV<0R=XR1ab5AsCHlR'&Rj&'RR''j,IRNH+8CL8IHC
2;RRRRRMRC8CRoMNCs0HCRV._NL
.;SFSOlCbDl0CMRR<=MRF0MEF1H;V0
0SSIFFOl<bR=FROlCbDl0CMR'+R4
';RRRRRCR)#0kDN=R<RhBmea_17m_pt_QBea Bmj)5,IRNH+8CL8IHCI2RERCM5RC4=jR"j
"2SSSSSCRRDR#CMEF1HRV0IMECR45CR"=Rj24"
SSSSRSRCCD#RF0IObFlRCIEMCR54RR=""442S
SSRSSR#CDCIR0FlOFbI5NH+8CL8IHCR-.8MFI0jFR2RR&';j'R-R-RCIEMCR54RR=""4j2C
SMo8RCsMCNR0CHNV_.
;
SR--v0kDH$bDRRL$0RECCsG0NHRL0H#RVCRIRPENCMRFCsRFRF0IR0CGsLNRHR0#FAVR
VSH_:L4RRHV5FLl82=4RMoCC0sNCR
RRRRRHLV_4:NjRVRHRl5NF<8R=RRjFNsRlRF8>2R.RMoCC0sNCS
SS#)CkLD0RR<=Bemh_71a_tpmQeB_ mBa),5jRHNI8LC+ICH82ERIC5MRCj.52RR='2j'RS
SSSSSRDRC#1CRXqa5blsHCN,RICH8+HLI8;C2
RRRRCRRMo8RCsMCNR0CHLV_4;Nj
HSSV4_LNR4:H5VRN8lFR4=R2CRoMNCs0SC
SCS)#0kDL=R<RhBmea_17m_pt_QBea Bmj)5,IRNH+8CL8IHCI2RERCM55C.j=2RR''j2SR
SSSSSCRRDR#C15XaqHbsl&CRR''j,IRNH+8CL8IHC
2;RRRRRMRC8CRoMNCs0HCRV4_LN
4;SVSH_NL4.H:RVNR5lRF8=2R.RMoCC0sNCS
SS#)CkLD0RR<=Bemh_71a_tpmQeB_ mBa),5jRHNI8LC+ICH82ERIC5MRCj.52RR='2j'RS
SSSSSRDRC#1CRXqa5blsHCRR&'Rj'&jR''N,RICH8+HLI8;C2
RRRRCRRMo8RCsMCNR0CHLV_4;N.
MSC8CRoMNCs0HCRV4_L;R
RRLHVMR.:H5VRL8lF=N.RML8RI0H8E2>.RMoCC0sNC-RR-hRz1hQt R7
RRRRRo#HMRNDMEF1H,V0RH#EV80C,8RN8RC8:0R#8F_Do_HOP0COFNs5ICH8+HLI84C-RI8FMR0Fj
2;SoLCHSM
SLHVMj.N:VRHRl5NF<8R=RRjFNsRlRF8>2R.RMoCC0sNCR
RRMSSFH1EV<0R=XR1ab5qsCHl,IRNH+8CL8IHC
2;RRRRRMRC8CRoMNCs0HCRV.LMN
j;SVSHLNM.4H:RVNR5lRF8=2R4RMoCC0sNCR
RRMSSFH1EV<0R=XR1ab5qsCHlR'&RjR',N8IHCI+LH28C;R
RRRRRCRM8oCCMsCN0RLHVM4.N;S
SHMVL.:N.RRHV5FNl8RR=.o2RCsMCN
0CRSRRS1MFE0HVRR<=15XaqHbsl&CRR''jR'&RjR',N8IHCI+LH28C;R
RRRRRCRM8oCCMsCN0RLHVM..N;S
S#VEH0RC8<M=RFH1EVN05ICH8+HLI8.C-RI8FMR0Fj&2RR''j;R
RRRRRNC888RRR<M=RFH1EV+0RRH#EV80C;S
S)kC#DR0L<B=Rm_he1_a7pQmtB _eB)am5Rj,N8IHCI+LH28CRCIEMCR5.RR=""jj2S
SSRSSR#CDCFRM1VEH0ERIC5MRC=.RR4"j"S2
SSSSRDRC##CRE0HVCI8RERCM5RC.=4R"j
"2SSSSSCRRDR#CNC888R;RRR--R.5CR"=R424"
MSC8CRoMNCs0HCRV.LM;H
SV._L:VRHRl5LF.8=R8NMRHLI8=0E.o2RCsMCNR0CRR--1hQt S7
So#HMRNDMEF1H,V0RlOFblDCC,M0RF0IObFlR#:R0D8_FOoH_OPC05FsN8IHCI+LH-8C4FR8IFM0R;j2
CSLo
HMRRRRRVRH_NL.jR:RH5VRN8lFRR<=jsRFRFNl8RR>.o2RCsMCN
0CRRRRRRRRR1MFE0HVRR<=15XaqHbslRC,N8IHCI+LH28C;S
SCRM8oCCMsCN0R_HVLj.N;S
SHLV_.:N4RRHV5FNl8RR=4o2RCsMCN
0CRSRRS1MFE0HVRR<=15XaqHbsl&CRR''j,IRNH+8CL8IHC
2;RRRRRMRC8CRoMNCs0HCRV._LN
4;SVSH_NL..H:RVNR5lRF8=2R.RMoCC0sNCR
RRMSSFH1EV<0R=XR1ab5qsCHlR'&Rj&'RR''j,IRNH+8CL8IHC
2;RRRRRMRC8CRoMNCs0HCRV._LN
.;SFSOlCbDl0CMRR<=MRF0MEF1H;V0
0SSIFFOl<bR=FROlCbDl0CMR'+R4
';SCS)#0kDL=R<RhBmea_17m_pt_QBea Bmj)5,IRNH+8CL8IHCI2RERCM5RC.=jR"j
"2SSSSSCRRDR#CMEF1HRV0IMECR.5CR"=Rj24"
SSSSRSRCCD#RF0IObFlRCIEMCR5.RR=""442S
SSRSSR#CDCIR0FlOFbI5NH+8CL8IHCR-48MFI0jFR2RR&';j'R-R-RCIEMCR5.RR=""4j2C
SMo8RCsMCNR0CHLV_.
;
SR--v0kDH$bDRC0ER0CGsLNRHR0#HIVRCNREPCCRGN0s#MRHR0CHERCsqMRN8
RAS_HVCR#:H5VR5FNl8RR=4sRFRFNl8RR=.N2RM58RL8lFR4=RRRFsL8lFR.=R2o2RCsMCN
0CSCS)#0kDC25dRR<=R5C44N2RMC8R425jR8NMR5C.4N2RMC8R.25j;S
S)kC#D50C.<2R=CR54254R8NMRF5M04RC52j2R8NMR5C.4R22FSs
SSSSS5RRC4452MRN8.RC5R42NRM850MFR5C.j222;S
S)kC#D50C4<2R=CR54254R8NMRF5M04RC52j2R8NMR5C.jR22FSs
SSSSS5RR50MFR5C44R22NRM8Cj452MRN8.RC5242R
FsSSSSSRSR55C44N2RM58RMRF0C4.52N2RMC8R.25j2sRF
SSSSRSSR45C5Rj2NRM8C4.52MRN8MR5FC0R.25j2
2;SCS)#0kDC25jRR<=R5C4jN2RMC8R.25j;S
SHsV_C:#CRRHV5HNI8LC+ICH8Rc>R2CRoMNCs0SC
SCS)#0kDCI5NH+8CL8IHCR-48MFI0cFR2=R<RhBmea_17m_pt_QBea Bmj)5,IRNH+8CL8IHCRR-c
2;SMSC8CRoMNCs0HCRVC_s#
C;S8CMRMoCC0sNCVRH_;C#
L
Sl0kD:VRHRHNI8>CRRN.RML8RICH8R.>RRMoCC0sNCS
Sl0kDG:GRRAe.pimB
SSSoCCMsRHOlRNb5S
SSSSSN8IH0=ER>IRNH
8,SSSSSISLHE80RR=>L8IH,S
SSSSSM8CC_bbHCVLk#>R=RCMC8H_bbkCLV
#2SbSSFRs0lRNb5S
SSqSSRRRR=q>RblsHCS,
SSSSARRRRR=>AHbsl
C,SSSSSmu)7>R=RF1Es20u;C
SMo8RCsMCNR0CLDlk0
;
RCRRGM0C8:H0RFbsO#C#RE51Fus02L
SCMoHR-R-RFbsO#C#R0CGCHM80R
RRRRR)kC#DR04<1=RX1a5E0FsuN,RICH8+HLI8;C2
MSC8sRbF#OC#GRC08CMH
0;
RRRNFLl8Rj:H5VR5FNl8R>.FNsRl=F8jN2RM58RL8lF>F.RslRLFj8=2o2RCsMCN
0CSCS)#0kDG=R<R#)Ck4D0;C
SMo8RCsMCNR0CNFLl8
j;
RRRNFLl8R4:H5VRN8lF=N4RM58RL8lF>F.RslRLFj8=2F2Rs5R5N8lF>F.RslRNFj8=2MRN8lRLF48=2CRoMNCs0SC
S#)CkGD0RR<=)kC#D504N8IHCI+LH-8C.FR8IFM0RRj2&jR''S;
CRM8oCCMsCN0RlNLF;84
R
RRlNLF:8.RRHV5FNl8R=4NRM8L8lF=R42F5sRN8lF=N.RM58RL8lF>F.RslRLFj8=2F2Rs5R5N8lF>F.RslRNFj8=2MRN8lRLF.8=2CRoMNCs0SC
S#)CkGD0RR<=)kC#D504N8IHCI+LH-8CdFR8IFM0RRj2&jR"j
";S8CMRMoCC0sNCLRNl.F8;R

RLRNldF8:VRHRl5NF.8=R8NMRFLl82=4RRFs5FNl8R=4NRM8L8lF=R.2oCCMsCN0
)SSCD#k0<GR=CR)#0kD4I5NH+8CL8IHCR-c8MFI0jFR2RR&"jjj"S;
CRM8oCCMsCN0RlNLF;8d
R
RRlNLF:8cRRHV5FNl8R=.NRM8L8lF=R.2oCCMsCN0
)SSCD#k0<GR=CR)#0kD4I5NH+8CL8IHCR-68MFI0jFR2RR&"jjjj
";S8CMRMoCC0sNCLRNlcF8;R

S_HVoCCMsCN0:VRHR555N8lFRj>R2MRN8NR5lRF8<2Rd2sRFRL55lRF8>2RjR8NMRl5LF<8RR2d22CRoMNCs0RC
RCRLo
HMSVSH_N#00:C4RRHV5l5NF>8RRRj2NRM85FNl8RR<dN2RM58RL8lFRj>R2MRN8LR5lRF8<2Rd2CRoMNCs0SC
SsSuF_84NRkG<R=R)kC#DR0N+CR)#0kDLRR+)kC#D;0C
CSSMo8RCsMCNR0CH#V_0CN04S;
S_HV#00NCR.:H5VR5FNl8RR>jN2RM58RN8lFRd<R2MRN85R5L8lFR.>R2sRFRl5LF=8RR2j22CRoMNCs0SC
SsSuF_84NRkG<R=R)kC#D;0N
CSSMo8RCsMCNR0CH#V_0CN0.S;
S_HV#00NCRd:H5VR5FLl8RR>jN2RM58RL8lFRd<R2MRN85R5N8lFR.>R2sRFRl5NF=8RR2j22CRoMNCs0SC
SsSuF_84NRkG<R=R)kC#D;0L
CSSMo8RCsMCNR0CH#V_0CN0d
;
SVSH_bbHNR4:H5VRM8CC_bbHCVLk#RR=4o2RCsMCN
0CSbSSHjbC:FRVsRRHHjMRRR0FI0H8ER-4oCCMsCN0
SSSS0N0skHL0\CR3MsN	F\RVCRsoR#1:NRDLRCDH4#R;S
SS0SN0LsHkR0C\C3Lo_HM0CsC\VRFRosC#:1RRLDNCHDR#;R4
SSSS0N0skHL0\CR3lsCF_PCMIF_N\sMRRFVs#Co1RR:DCNLD#RHR
4;SLSSCMoH
SSSSosC#R1:RbbHCVLk
SSSSsbF0NRlbS5
SSSSS=QR>sRuF_84N5kGH
2,SSSSSRSm=u>Rs4F8_#sC52H2;S
SS8CMRMoCC0sNCHRbb;Cj
CSSMo8RCsMCNR0CHbV_H4bN;S
SHbV_HjbN:VRHRC5MCb8_HLbCkRV#=2RjRMoCC0sNCS
SSFus8s4_C<#R=sRuF_84N;kG
CSSMo8RCsMCNR0CHbV_HjbN;C
SMo8RCsMCNR0CHoV_CsMCN;0C
S
RHoV_CsMCN_0C4H:RV5R5N8lFR.>R2MRN8LR5lRF8>2R.2CRoMNCs0SC
SFus8s4_C<#R=BRRm_he1_a7pQmtB _eB)am5Rj,N8IHCI+LH28C;C
SMo8RCsMCNR0CHoV_CsMCN_0C4
;
RuRRs4F8RR<=)kC#DR0G+sRuF_84s;C#
C
SGM0C8Fbs8b:RsCFO#5#Ru8sF4S2
LHCoM-RR-sRbF#OC#GRC08CMb8sF
HSSVHRI8R0E>IRNHR8C+IRLHR8C0MEC
SSSu8sF.=R<Ra1X5Fus8R4,I0H8E
2;SDSC#SC
SsSuFR8.<u=Rs4F858IH04E-RI8FMR0Fj
2;SMSC8VRH;C
SMb8RsCFO#C#RGM0C8Fbs8
;
S_HVbLHb4H:RVMR5C_C8bCHbL#kVR4=R2CRoMNCs0SC
SVLkFbk0kR0:VRFsHMRHR0jRFHRI8-0E4CRoMNCs0SC
S0SN0LsHkR0C\N3sMR	\FsVRC1o#RD:RNDLCRRH#.S;
S0SN0LsHkR0C\M3C8s_0CRC\FsVRC1o#RD:RNDLCRRH#4S;
S0SN0LsHkR0C\F3b8\ClRRFVs#Co1RR:DCNLD#RHR
H;SNSS0H0sLCk0Rb\3Fl8CL\k#RRFVs#Co1RR:DCNLD#RHR)"um;7"
SSSNs00H0LkC3R\sFClPMC_FN_IsRM\FsVRC1o#RD:RNDLCRRH#4S;
SoLCHSM
SCSso:#1RHRbbkCLVS
SSbSSFRs0l5Nb
SSSSSSSQ>R=RFus8H.52S,
SSSSSRSm=u>R)5m7H;22
CSSMo8RCsMCNR0CLFkVkk0b0S;
CRM8oCCMsCN0R_HVbLHb4S;
HbV_HjbL:VRHRC5MCb8_HLbCkRV#=2RjRMoCC0sNCS
Su7)mRR<=u8sF.S;
CRM8oCCMsCN0R_HVbLHbj
;
CRM8LODF	k_lD
0;
