DDggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggDggDggZ}��������ZksspZ��Z�hZ{��Z������Z��������hDggDggZ����Z������Z����Z��Z��Z���������Z����Z��Z�Z���ZkjqphlgksspfZ�Z��������ZDggZ��~�Z������������Z��������hZ����Z������Z����Z���Z���Z��Z������fZ����fZ��ZDggZ��������Z����Z��������Z����Z��Z����Z�������Z�������Z����������Z����Z���Z�DggZ���������Z~���������hZ����Z������Z����Z���Z��Z����Z��Z���������Z����Z��������ZDggZ���Z���Z��Z�����������Z��Z��������Z����Z��Z���Z������Z��Z����Z��Z���ZDggZ��������Z����Z����Z���Z�����Z������Z�������������Z��Z���Z��������Z������Z����hDggZ����Z������Z����Z���Z��Z������Z���Z����������Z���Z�������Z��������Z�����hZDggZ����Z������Z����Z��Z��������Z��Z��Z{�Z��Z�����hZ���Z�Z���������Z{��ZDggZ�{��{���Z�����Z��Z�����~Z��}��~���Z{��Z�{��{���Z��Z��}�{��{|�����ZDggZ{�~Z������Z���Z��Z���Z{Z�{���}��{�Z������hZ���Z����Z��Z���Z������ZDggZ����Z�����Z���������Z���Z����Z�Z��������Z����Z���Z�������Z��Z���������ZDggZ�������Z���Z��Z���Z���Z�������hDggDggZ�����tZZZZZZZ��������Z��~�Z������������Z��������Zb�Z���ZkjqphlgksspfZDggZZZZZZZZZZZZZZ�{����{�cDggDggZ�������tZZZZZ����Z�������Z�����Z��Z��������Z����Z�Z�������DggZZZZZZZZZZZZZZ������������Z�����Z�hDggDggZ~���������tZZ�Z~{�}Z��~�Z������������Z��������Z�������Z�����DggDggZ�������tZZZZZ����Z�������Z�������Z�Z��������Z���Z���������Z��Z���Z��DggZZZZZZZZZZZZZZ����������Z��~�Z������Z����Z����Z���Z��Z������Z�{�Z���������DggZZZZZZZZZZZZZZ���Z������Z�{�Z����������Z������������Z���������hDggDggZ����������tZZ���Z������Z���������Z��Z���Z���������Z��Z����Z�������Z���DggZZZZZZZZZZZZZZ����Z����Z��������Z��Z��������fZ���Z���Z���������Z��Z�������DggZZZZZZZZZZZZZZ��Z����Z����������Z��Z��Z���Z�������Z��������Z��Z�Z���ZkjqpgDggZZZZZZZZZZZZZZkssmhDggDggZ�����tDggZZZZZZZZZZZZZZ��Z������������Z��Z�����������Z�����Z��Z��������Z��fZ��DggZZZZZZZZZZZZZZ��������Z����fZ����Z�������hDggZZZZZZZZZZZZZZ���Z\�������Z�����������\Z�������Z���Z�����fZ��������fZ���DggZZZZZZZZZZZZZZ������������Z��Z�{����{�hDggZZZZZZZZZZZZZZ���Z��������Z������������Z����������Z���Z������������Z�������DggZZZZZZZZZZZZZZ��Z���Z������������Z���������Z����Z���Z����Z��Z����Z��������DggZZZZZZZZZZZZZZ���������Z���Z������Z���������Z��Z���Z��������������Z��Z���DggZZZZZZZZZZZZZZ�{����{�Z�������Z�����������hZZ���Z�������Z��Z���Z�{����{�DggZZZZZZZZZZZZZZ�������Z����Z��Z��Z�������Z�Z���������Z���Z���������������Z��DggZZZZZZZZZZZZZZ������Z�����Z��������������Z��Z�{����{�hZZ����Z����������Z���DggZZZZZZZZZZZZZZ������Z��Z���������Z���Z�������Z����Z��Z���Z����Z���������DggZZZZZZZZZZZZZZ������Z���������Z��Z����hDggDggZgggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggDggZ�������ZZZZtZkhoDggZ~���ZZZZZZZtZlnZ����ZksspDggZgggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggDD�������Z�{����{�Z��DZZZZ��������Z}��������������tZ������DZZZZZZtwZ\}��������ZksspZ�hZ{��Z������Z��������h\uDDZZZZggDZZZZggZ}�������Z~����������DZZZZggDZZZZ��������ZZ�{���ZtZ�{�ZtwZlhqkrlr�krlrn�osjno�lmompuDZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZggZ�����Z��Z�DZZZZ��������ZZ�{���k�����ZtZ�{�ZtwZjhmpqrq�snnkk�qknnl�mlkpjuDZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZggZ�����Z��Zki�DZZZZ��������ZZ�{�����ZtZ�{�ZtwZmhknkos�lpomo�rsqsm�lmrnpuDZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZggZ�����Z��Z��DZZZZ��������ZZ�{���l���ZtZ�{�ZtwZphlrmkr�omjqk�qsorp�nqpsmuDZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZggZ�����Z��Zld��DZZZZ��������ZZ�{���k�������ZtZ�{�ZtwZjhmkrmj�srrpk�rmqsj�pqkonuDZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZggZ�����Z��Zki��DZZZZ��������ZZ�{����������lZtZ�{�ZtwZkhoqjqs�pmlpq�snrsp�pkslmuDZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZggZ�����Z��Z��ilDZZZZ��������ZZ�{����������mZtZ�{�ZtwZkhjnqks�qookk�sposq�qnpkouDZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZggZ�����Z��Z��imDZZZZ��������ZZ�{����������nZtZ�{�ZtwZjhqroms�rkpmm�sqnnr�mjspluDZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZggZ�����Z��Z��inDZZZZ��������ZZ�{���m��������lZtZ�{�ZtwZnhqklmr�rsrjm�rnprs�roqpsuDZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZggZ�����Zmd��ilDZZZZ��������ZZ�{����������lZtZ�{�ZtwZjhpsmkn�qkrjo�ossno�mjsnluDZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZggZ�������Z���Z��ZlDZZZZ��������ZZ�{����������kjZtZ�{�ZtwZlhmjlor�ojsls�snjno�prnjluDZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZggZ�������Z���Z��ZkjDZZZZ��������ZZ�{������l����ZtZ�{�ZtwZkhnnlps�ojnjr�rrspm�njqnuDZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZggZ���Z����ZlZ��Z�DZZZZ��������ZZ�{������kj����tZ�{�ZtwZjhnmnls�nnrks�jmlok�rlqpouDZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZggZ���Z����ZkjZ��Z�DZZZZ��������ZZ�{��������ltZ�{�ZtwZkhnknlk�moplm�qmjso�jnrrjuDZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZggZ������Z����Z��ZlDZZZZ��������ZZ�{���k����������ltZ�{�ZtwZjhqjqkj�pqrkk�rponq�olnnjuDZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZggZ������Z����Z��ZkilDZZZZ��������ZZ�{����������tZ�{�ZtwZkhqqlno�mrojs�jookp�jlqmjuDZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZggZ������Z����Z��Z��DZZZZ��������ZZ�{���~������{~tZ�{�ZtwZjhjkqno�mlslo�kssnm�lsoqquDZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZggZ}���������Z������Z����Z������Z��Z������DZZZZ��������ZZ�{����{~����~�tZ�{�ZtwZoqhlsoqq�sokmj�rlmlj�rqprjuDZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZggZ}���������Z������Z����Z������Z��Z������DDZZZZggDZZZZggZ��������Z~�����������DZZZZggDZZZZ��������Z����Zb�tZ��Z�{�ZcZ������Z�{�uDZZZZZZZZggZ�������tDZZZZZZZZggZZZZZZZZZ�������ZkhjZ��Z�ZxZjhjuZjhjZ��Z�ZwZjhjuZgkhjZ��Z�ZvZjhjDZZZZZZZZggZ�������Z������tDZZZZZZZZggZZZZZZZZZ����DZZZZZZZZggZ~�����tDZZZZZZZZggZZZZZZZZZ�Z��Z�{�DZZZZZZZZggZ����Z����������tDZZZZZZZZggZZZZZZZZZ����DZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZZ{|�b����b�ccZvwZkhjDZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZZ����DDZZZZ��������Z}��Zb�ZtZ��Z�{�ZcZ������Z�{�uDZZZZZZZZggZ�������tDZZZZZZZZggZZZZZZZZZ�������Z��������Z�����Z�����Zb��Z�{�cZ���Z����Z����Z�DZZZZZZZZggZ�������Z������tDZZZZZZZZggZZZZZZZZZ����DZZZZZZZZggZ~�����tDZZZZZZZZggZZZZZZZZZ�Z��Z�{�DZZZZZZZZggZ����Z����������tDZZZZZZZZggZZZZZZZZZ����DZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZZ}��b�cZ��Z��������������Z���������DZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZZ�cZ���������������Z����Z��Z�������Z��Z�����Z���Z������DZZZZZZZZggZZZZZZZZZZZZZZZZ{|�b�cZvZ�{�b�����a����cDDZZZZ��������Z�����Zb�ZtZ��Z�{�ZcZ������Z�{�uDZZZZZZZZggZ�������tDZZZZZZZZggZZZZZZZZZ�������Z�������Z�����Z�����Zb��Z�{�cZ���Z�������Z����Z�DZZZZZZZZggZ�������Z������tDZZZZZZZZggZZZZZZZZZ�����bjhjcZwZjhjDZZZZZZZZggZ~�����tDZZZZZZZZggZZZZZZZZZ�Z��Z�{�DZZZZZZZZggZ����Z����������tDZZZZZZZZggZZZZZZZZZ����DZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZZ�����b�cZ��Z��������������Z���������DZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZZ�cZ���������������Z����Z��Z�������Z��Z�����Z���Z������DZZZZZZZZggZZZZZZZZZZZZZZZZ{|�b�cZvZ�{�b�����a����cDDZZZZ��������Z����~Zb�ZtZ��Z�{�ZcZ������Z�{�uDZZZZZZZZggZ�������tDZZZZZZZZggZZZZZZZZZ������Z�Z��Z���Z�������Z�������Z�����Zb��Z����chZ��Z�Z��DZZZZZZZZggZZZZZZZZZ�������Z�������Z���Z��������fZ��������Z��Z����Z����ZjhjDZZZZZZZZggZ�������Z������tDZZZZZZZZggZZZZZZZZZ����~bjhjcZwZjhjDZZZZZZZZggZ~�����tDZZZZZZZZggZZZZZZZZZ�Z��Z�{�DZZZZZZZZggZ����Z����������tDZZZZZZZZggZZZZZZZZZ����DZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZZ����~b�cZ��Z��������������Z���������DZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZZ�cZ���������������Z����Z��Z�������Z��Z�����Z���Z������DZZZZZZZZggZZZZZZZZZZZZZZZZ{|�b�cZvZ�{�b�����a����cDDZZZZ��������Z����}Zb�ZtZ��Z�{�ZcZ������Z�{�uDZZZZZZZZggZ�������tDZZZZZZZZggZZZZZZZZZ���������Z�Z�������ZjhjZ���Z�������Z���������Z�����DZZZZZZZZggZ�������Z������tDZZZZZZZZggZZZZZZZZZ����}bjhjcZwZjhjDZZZZZZZZggZ~�����tDZZZZZZZZggZZZZZZZZZ�Z��Z�{�DZZZZZZZZggZ����Z����������tDZZZZZZZZggZZZZZZZZZ����DZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZZ����}b�cZ��Z��������������Z���������DZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZZ�cZ���������������Z����Z��Z�������Z��Z�����Z���Z������DZZZZZZZZggZZZZZZZZZZZZZZZZ{|�b�cZvZ�{�b�����a����cDDZZZZ��������Z\��~\Zb�fZ�tZ��Z�{�ZcZ������Z�{�uDZZZZZZZZggZ�������tDZZZZZZZZggZZZZZZZZZ�������Z��������Z�����Z�������Z��Z�i�fZ����Z���Z����Z����Z��DZZZZZZZZggZZZZZZZZZ�fZ���Z��������Z�����Z����Z����Z���Z��������Z�����Z��Z�fZ���DZZZZZZZZggZZZZZZZZZ���Z����Z�����Z�����Z�Z���Z������Z���������Z���Z��������DZZZZZZZZggZZZZZZZZZ�ZwZ�d�ZeZ��~b�f�cDZZZZZZZZggZ�������Z������tDZZZZZZZZggZZZZZZZZZ����DZZZZZZZZggZ~�����tDZZZZZZZZggZZZZZZZZZ�Z��Z�{�uZ�Z��Z�{�Z���Z�ZiwZjhjDZZZZZZZZggZ����Z����������tDZZZZZZZZggZZZZZZZZZ����Z��Z�ZwZjhjDZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZZ{|�b��~b�f�ccZvZ{|�b�cDZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZZ����DDZZZZ��������Z�{��{�Zb�fZ�ZtZ��Z�{�ZcZ������Z�{�uDZZZZZZZZggZ�������tDZZZZZZZZggZZZZZZZZZ�������Z���Z�������������Z������Z��Z�Z���Z�DZZZZZZZZggZ�������Z������tDZZZZZZZZggZZZZZZZZZ�{��{�b�f�cZwZ�Z����Z�ZwZ�DZZZZZZZZggZ~�����tDZZZZZZZZggZZZZZZZZZ�Z��Z�{�uZ�Z��Z�{�DZZZZZZZZggZ����Z����������tDZZZZZZZZggZZZZZZZZZ����DZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZZ�{��{�b�f�cZ��Z��������������Z���������DZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZZ����DDZZZZ��������Z�{����Zb�fZ�ZtZ��Z�{�ZcZ������Z�{�uDZZZZZZZZggZ�������tDZZZZZZZZggZZZZZZZZZ�������Z���Z�������������Z�������Z��Z�Z���Z�DZZZZZZZZggZ�������Z������tDZZZZZZZZggZZZZZZZZZ�{����b�f�cZwZ�Z����Z�ZwZ�DZZZZZZZZggZ~�����tDZZZZZZZZggZZZZZZZZZ�Z��Z�{�uZ�Z��Z�{�DZZZZZZZZggZ����Z����������tDZZZZZZZZggZZZZZZZZZ����DZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZZ�{����b�f�cZ��Z��������������Z���������DZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZZ����DDZZZZ���������Z�������b��������Z�~kf�~lt�����Z�������uZ��������Z�t���Z�{�cuDZZZZZZZZggZ�������tDZZZZZZZZggZZZZZZZZZ�������fZ��Z�fZ�Z������g������Z������Z����Z�������DZZZZZZZZggZZZZZZZZZ������������Z��Z���Z����Z��������ZbjhjfZkhjchDZZZZZZZZggZ�������Z������tDZZZZZZZZggZZZZZZZZZ����DZZZZZZZZggZ~�����tDZZZZZZZZggZZZZZZZZZkZvwZ�~kZvwZlknqnrmopluZkZvwZ�~lZvwZlknqnrmmsrDZZZZZZZZggZ����Z����������tDZZZZZZZZggZZZZZZZZZ����Z��Z�~kZ��Z�~lZ�������Z��Z�����Z������DZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZZjhjZvZ�ZvZkhjDZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZZ�cZ���Z���������Z���Z����Z��������Z���Z���������Z��Z���DZZZZZZZZggZZZZZZZZZZZZ���������Z���������Z��Z������Z�a�����Z��Z\}�������������DZZZZZZZZggZZZZZZZZZZZZ��Z���Z{}�f\Z���hZmkfZ��hZpfZ����ZksrrfZ��hZqnlgqqnhDZZZZZZZZggZZZZZZZZZZZZ���Z���������Z��Z�����Z��Z���Z�����������Z��Z���DZZZZZZZZggZZZZZZZZZZZZ��������������Z������Z������������Z����������Z���Zmlg���DZZZZZZZZggZZZZZZZZZZZZ���������hDZZZZZZZZggDZZZZZZZZggZZZZZZZZZ�cZ|�����Z���Z�����Z����Z��Z�������fZ���Z����Z������DZZZZZZZZggZZZZZZZZZZZZb�~kfZ�~lcZ����Z��Z��Z�����������Z��Z������Z��Z���Z�����DZZZZZZZZggZZZZZZZZZZZZ�kfZlknqnrmopl�Z���Z�kfZlknqnrmmsr�Z������������hZZ���DZZZZZZZZggZZZZZZZZZZZZ����Z������Z���Z��������Z�����Z����Z����Z��Z�������hDZZZZZZZZggDZZZZZZZZggZZZZZZZZZ�cZ����Z������Z������Z���������Z��Z��������Z���Zmlg���DZZZZZZZZggZZZZZZZZZZZZ���������fZ���Z��Z���Z�Z������Z��Z�lhmjorndbkjddkrcZ���Z����DZZZZZZZZggZZZZZZZZZZZZ���Z��Z����Z������hDZZZZZZZZggDZZZZZZZZggZZZZZZZZZ�cZ���Z�����������Z��Z��������Z�����Z���Z���Z���������fZ�����DZZZZZZZZggZZZZZZZZZZZZ��Z���Z�a�����Z�������hDDZZZZ��������Z����Zb�ZtZ��Z�{�ZcZ������Z�{�uDZZZZZZZZggZ�������tDZZZZZZZZggZZZZZZZZZ�������Z������Z����Z��Z�DZZZZZZZZggZ�������Z������tDZZZZZZZZggZZZZZZZZZ����bjhjcZwZjhjDZZZZZZZZggZZZZZZZZZ����bkhjcZwZkhjDZZZZZZZZggZ~�����tDZZZZZZZZggZZZZZZZZZ�ZxwZjhjDZZZZZZZZggZ����Z����������tDZZZZZZZZggZZZZZZZZZ����Z��Z�ZvZjhjDZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZZ����b�cZxwZjhjDZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZZ�cZ���Z�����Z�����Z��Z���Z���������Z�����Z��Z����Z��DZZZZZZZZggZZZZZZZZZZZZ�������������Z�����Z��tDZZZZZZZZggZZZZZZZZZZZZZZZZ����b�cZvwZ����b�{�a����cDDZZZZ��������Z}|��Zb�ZtZ��Z�{�ZcZ������Z�{�uDZZZZZZZZggZ�������tDZZZZZZZZggZZZZZZZZZ�������Z����Z����Z��Z�DZZZZZZZZggZ�������Z������tDZZZZZZZZggZZZZZZZZZ}|��bjhjcZwZjhjDZZZZZZZZggZZZZZZZZZ}|��bkhjcZwZkhjDZZZZZZZZggZZZZZZZZZ}|��bgkhjcZwZgkhjDZZZZZZZZggZ~�����tDZZZZZZZZggZZZZZZZZZ�Z��Z�{�DZZZZZZZZggZ����Z����������tDZZZZZZZZggZZZZZZZZZ����DZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZZ}|��b�cZ��Z��������������Z���������DZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZZ�cZ���Z���������Z�����Z��Z}|��Z��Z�������������Z�����Z��tDZZZZZZZZggZZZZZZZZZZZZZZZZ{|�b}|��b�ccZvwZ}|��b�{�a����cDDZZZZ��������Z\dd\Zb�ZtZ��Z�����uZ�ZtZ��Z�{�cZ������Z�{�uDZZZZZZZZggZ�������tDZZZZZZZZggZZZZZZZZZ�������Z�Z�����Z��Z�ZwwxZZ�dd�DZZZZZZZZggZ�������Z������tDZZZZZZZZggZZZZZZZZZ�ddjhjZwZkhjuZ�ZiwZjDZZZZZZZZggZZZZZZZZZjdd�ZwZjhjuZ�ZxZjhjDZZZZZZZZggZZZZZZZZZ�ddkhjZwZ�{�b�cuZ�ZxwZjDZZZZZZZZggZZZZZZZZZkdd�ZwZkhjDZZZZZZZZggZ~�����tDZZZZZZZZggZZZZZZZZZ�ZxZjDZZZZZZZZggZZZZZZZZZ�ZwZjZ���Z�ZxZjhjDZZZZZZZZggZZZZZZZZZ�ZvZjZ���Z�ZwZjhjDZZZZZZZZggZ����Z����������tDZZZZZZZZggZZZZZZZZZ����Z��Z�ZvZjZ���Z�ZiwZjhjDZZZZZZZZggZZZZZZZZZ����Z��Z�ZwZjZ���Z�ZvwZjhjDZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZZ�dd�ZxwZjhjDZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZZ�cZ���Z�����Z�����Z��Z���Z���������Z�����Z���Z\dd\Z��DZZZZZZZZggZZZZZZZZZZZZ�������������Z�����Z��tDZZZZZZZZggZZZZZZZZZZZZZZZZ�dd�ZvwZ�{�a����DDZZZZ��������Z\dd\Zb�ZtZ��Z�{�uZ�ZtZ��Z�{�cZ������Z�{�uDZZZZZZZZggZ�������tDZZZZZZZZggZZZZZZZZZ�������Z�Z�����Z��Z�ZwwxZZ�dd�DZZZZZZZZggZ�������Z������tDZZZZZZZZggZZZZZZZZZ�ddjhjZwZkhjuZ�ZiwZjhjDZZZZZZZZggZZZZZZZZZjhjdd�ZwZjhjuZ�ZxZjhjDZZZZZZZZggZZZZZZZZZ�ddkhjZwZ�uZ�ZxwZjhjDZZZZZZZZggZZZZZZZZZkhjdd�ZwZkhjDZZZZZZZZggZ~�����tDZZZZZZZZggZZZZZZZZZ�ZxZjhjDZZZZZZZZggZZZZZZZZZ�ZwZjhjZ���Z�ZxZjhjDZZZZZZZZggZZZZZZZZZ�ZvZjhjZ���Z�ZwZjhjDZZZZZZZZggZ����Z����������tDZZZZZZZZggZZZZZZZZZ����Z��Z�ZvZjhjZ���Z�ZiwZjhjDZZZZZZZZggZZZZZZZZZ����Z��Z�ZwZjhjZ���Z�ZvwZjhjDZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZZ�dd�ZxwZjhjDZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZZ�cZ���Z�����Z�����Z��Z���Z���������Z�����Z���Z\dd\Z��DZZZZZZZZggZZZZZZZZZZZZ�������������Z�����Z��tDZZZZZZZZggZZZZZZZZZZZZZZZZ�dd�ZvwZ�{�a����DDZZZZ��������Z��Zb�ZtZ��Z�{�ZcZ������Z�{�uDZZZZZZZZggZ�������tDZZZZZZZZggZZZZZZZZZ�������Z�dd�uZ�����Z�ZwZ�{���DZZZZZZZZggZ�������Z������tDZZZZZZZZggZZZZZZZZZ��bjhjcZwZkhjDZZZZZZZZggZZZZZZZZZ��bkhjcZwZ�{���DZZZZZZZZggZZZZZZZZZ��bgkhjcZwZ�{���k�����DZZZZZZZZggZZZZZZZZZ��b�cZwZjhjZ���Z�ZvwZg���b�{�a����cDZZZZZZZZggZ~�����tDZZZZZZZZggZZZZZZZZZ�Z��Z�{�Z����Z����Z��b�cZvwZ�{�a����DZZZZZZZZggZ����Z����������tDZZZZZZZZggZZZZZZZZZ����Z��Z�ZxZ���b�{�a����cDZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZZ��b�cZxwZjhjDZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZZ�cZ���Z������Z������Z��Z��Z��Z�������������Z�����Z��tDZZZZZZZZggZZZZZZZZZZZZZZZZ�ZvwZ���b�{�a����cDDZZZZ��������Z���Zb�ZtZ��Z�{�ZcZ������Z�{�uDZZZZZZZZggZ�������tDZZZZZZZZggZZZZZZZZZ�������Z�������Z���������Z��Z�DZZZZZZZZggZ�������Z������tDZZZZZZZZggZZZZZZZZZ���bkhjcZwZjhjDZZZZZZZZggZZZZZZZZZ���b�{���cZwZkhjDZZZZZZZZggZ~�����tDZZZZZZZZggZZZZZZZZZ�ZxZjhjDZZZZZZZZggZ����Z����������tDZZZZZZZZggZZZZZZZZZ����Z��Z�ZvwZjhjDZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZZ���b�cZ��Z��������������Z���������DZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZZ�cZ���Z���������Z�����Z��Z���Z��Z�������������Z�����Z��tDZZZZZZZZggZZZZZZZZZZZZZZZZ���bjecZvwZ���b�cZvwZ���b�{�a����cDDZZZZ��������Z���lZb�ZtZ��Z�{�ZcZ������Z�{�uDZZZZZZZZggZ�������tDZZZZZZZZggZZZZZZZZZ�������Z���������Z����ZlZ��Z�DZZZZZZZZggZ�������Z������tDZZZZZZZZggZZZZZZZZZ���lbkhjcZwZjhjDZZZZZZZZggZZZZZZZZZ���lblhjcZwZkhjDZZZZZZZZggZ~�����tDZZZZZZZZggZZZZZZZZZ�ZxZjhjDZZZZZZZZggZ����Z����������tDZZZZZZZZggZZZZZZZZZ����Z��Z�ZvwZjhjDZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZZ���lb�cZ��Z��������������Z���������DZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZZ�cZ���Z���������Z�����Z��Z���lZ��Z�������������Z�����Z��tDZZZZZZZZggZZZZZZZZZZZZZZZZ���lbjecZvwZ���lb�cZvwZ���lb�{�a����cDDZZZZ��������Z���kjZb�ZtZ��Z�{�ZcZ������Z�{�uDZZZZZZZZggZ�������tDZZZZZZZZggZZZZZZZZZ�������Z���������Z����ZkjZ��Z�DZZZZZZZZggZ�������Z������tDZZZZZZZZggZZZZZZZZZ���kjbkhjcZwZjhjDZZZZZZZZggZZZZZZZZZ���kjbkjhjcZwZkhjDZZZZZZZZggZ~�����tDZZZZZZZZggZZZZZZZZZ�ZxZjhjDZZZZZZZZggZ����Z����������tDZZZZZZZZggZZZZZZZZZ����Z��Z�ZvwZjhjDZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZZ���kjb�cZ��Z��������������Z���������DZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZZ�cZ���Z���������Z�����Z��Z���kjZ��Z�������������Z�����Z��tDZZZZZZZZggZZZZZZZZZZZZZZZZ���kjbjecZvwZ���kjb�cZvwZ���kjb�{�a����cDDZZZZ��������Z���Zb�tZ��Z�{�uZ|{�tZ��Z�{�cZ������Z�{�uDZZZZZZZZggZ�������tDZZZZZZZZggZZZZZZZZZ�������Z���������Z����Z|{�Z��Z�DZZZZZZZZggZ�������Z������tDZZZZZZZZggZZZZZZZZZ���bkhjfZ|{�cZwZjhjDZZZZZZZZggZZZZZZZZZ���b|{�fZ|{�cZwZkhjDZZZZZZZZggZ~�����tDZZZZZZZZggZZZZZZZZZ�ZxZjhjDZZZZZZZZggZZZZZZZZZ|{�ZxZjhjDZZZZZZZZggZZZZZZZZZ|{�ZiwZkhjDZZZZZZZZggZ����Z����������tDZZZZZZZZggZZZZZZZZZ����Z��Z�ZvwZjhjDZZZZZZZZggZZZZZZZZZ����Z��Z|{�ZvwZjhjDZZZZZZZZggZZZZZZZZZ����Z��Z|{�ZwZkhjDZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZZ���b�fZ|{�cZ��Z��������������Z���������DZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZZ�cZ����Z|{�ZxZkhjfZ���Z���������Z�����Z��Z���Z��DZZZZZZZZggZZZZZZZZZZZZ�������������Z�����Z��tDZZZZZZZZggZZZZZZZZZZZZZZZZ���bjefZ|{�cZvwZ���b�fZ|{�cZvwZ���b�{�a����fZ|{�cDZZZZZZZZggZZZZZZZZZ�cZ����ZjhjZvZ|{�ZvZkhjfZ���Z���������Z�����Z��Z���Z��DZZZZZZZZggZZZZZZZZZZZZ�������������Z�����Z��tDZZZZZZZZggZZZZZZZZZZZZZZZZ���b�{�a����fZ|{�cZvwZ���b�fZ|{�cZvwZ���bjefZ|{�cDDZZZZ��������ZZ���Zb�ZtZ��Z�{�ZcZ������Z�{�uDZZZZZZZZggZ�������tDZZZZZZZZggZZZZZZZZZ�������Z����Z��Z�uZ�Z��Z�������DZZZZZZZZggZ�������Z������tDZZZZZZZZggZZZZZZZZZ���b�cZwZjhjZ���Z�ZwZ�d�{�����fZ�����Z�Z��Z��Z�����DZZZZZZZZggZZZZZZZZZ���b�cZwZkhjZ���Z�ZwZbnd�ekcd�{����������lfZ�����Z�Z��Z��DZZZZZZZZggZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ�����DZZZZZZZZggZZZZZZZZZ���b�cZwZgkhjZ���Z�ZwZbnd�emcd�{����������lfZ�����Z�Z��Z��DZZZZZZZZggZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ�����DZZZZZZZZggZ~�����tDZZZZZZZZggZZZZZZZZZ�Z��Z�{�DZZZZZZZZggZ����Z����������tDZZZZZZZZggZZZZZZZZZ����DZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZZ{|�b���b�ccZvwZkhjDZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZZ�cZ���Z������Z������Z��Z{|�b�cfZ��������Z��������Z��Z�������hDDZZZZ��������ZZ}��ZbZ�ZtZ��Z�{�ZcZ������Z�{�uDZZZZZZZZggZ�������tDZZZZZZZZggZZZZZZZZZ�������Z������Z��Z�uZ�Z��Z�������DZZZZZZZZggZ�������Z������tDZZZZZZZZggZZZZZZZZZ}��b�cZwZjhjZ���Z�ZwZbld�ekcd�{����������lfZ�����Z�Z��Z��DZZZZZZZZggZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ�����DZZZZZZZZggZZZZZZZZZ}��b�cZwZkhjZ���Z�ZwZbld�cd�{�����fZ�����Z�Z��Z��Z�����DZZZZZZZZggZZZZZZZZZ}��b�cZwZgkhjZ���Z�ZwZbld�ekcd�{�����fZ�����Z�Z��Z��Z�����DZZZZZZZZggZ~�����tDZZZZZZZZggZZZZZZZZZ�Z��Z�{�DZZZZZZZZggZ����Z����������tDZZZZZZZZggZZZZZZZZZ����DZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZZ{|�b}��b�ccZvwZkhjDZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZZ�cZ���Z������Z������Z��Z{|�b�cfZ��������Z��������Z��Z�������hDDZZZZ��������ZZ�{�Zb�ZtZ��Z�{�ZcZ������Z�{�uDZZZZZZZZggZ�������tDZZZZZZZZggZZZZZZZZZ�������Z�������Z��Z�uZ�Z��Z�������DZZZZZZZZggZ�������Z������tDZZZZZZZZggZZZZZZZZZ�{�b�cZwZjhjZ���Z�ZwZ�d�{�����fZ�����Z�Z��Z��Z�����DZZZZZZZZggZ~�����tDZZZZZZZZggZZZZZZZZZ�Z��Z�{�Z���DZZZZZZZZggZZZZZZZZZ�ZiwZbld�ekcd�{����������lfZ�����Z�Z��Z��Z�����DZZZZZZZZggZ����Z����������tDZZZZZZZZggZZZZZZZZZ����Z��Z�ZwZbbld�ekcZdZ�{����������lcfZ�����Z�Z��Z��DZZZZZZZZggZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ�����DZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZZ�{�b�cZ��Z��������������Z���������DZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZZ�cZ���Z������Z������Z��Z{|�b�cfZ��������Z��������Z��Z�������hDDZZZZ��������ZZ{�}���Zb�ZtZ��Z�{�ZcZ������Z�{�uDZZZZZZZZggZ�������tDZZZZZZZZggZZZZZZZZZ�������Z�������Z����Z��Z�DZZZZZZZZggZ�������Z������tDZZZZZZZZggZZZZZZZZZ{�}���bjhjcZwZjhjDZZZZZZZZggZZZZZZZZZ{�}���bkhjcZwZ�{����������lDZZZZZZZZggZZZZZZZZZ{�}���bgkhjcZwZg�{����������lDZZZZZZZZggZ~�����tDZZZZZZZZggZZZZZZZZZ{|�b�cZvwZkhjDZZZZZZZZggZ����Z����������tDZZZZZZZZggZZZZZZZZZ����Z��Z{|�b�cZxZkhjDZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZZ{|�b{�}���b�cZvwZ�{����������lDZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZZ����DDZZZZ��������ZZ{�}}��Zb�ZtZ��Z�{�ZcZ������Z�{�uDZZZZZZZZggZ�������tDZZZZZZZZggZZZZZZZZZ�������Z�������Z������Z��Z�DZZZZZZZZggZ�������Z������tDZZZZZZZZggZZZZZZZZZ{�}}��bkhjcZwZjhjDZZZZZZZZggZZZZZZZZZ{�}}��bjhjcZwZ�{����������lDZZZZZZZZggZZZZZZZZZ{�}}��bgkhjcZwZ�{�����DZZZZZZZZggZ~�����tDZZZZZZZZggZZZZZZZZZ{|�b�cZvwZkhjDZZZZZZZZggZ����Z����������tDZZZZZZZZggZZZZZZZZZ����Z��Z{|�b�cZxZkhjDZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZZjhjZvwZ{�}}��b�cZvwZ�{�����DZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZZ����DDZZZZ��������ZZ{�}�{�Zb�ZtZ��Z�{�cZ������Z�{�uDZZZZZZZZggZ�������tDZZZZZZZZggZZZZZZZZZ�������Z���Z�����Z��Z���Z�����Z��Z�������Z��Z���Z�����DZZZZZZZZggZZZZZZZZbkhjfZ�cfZ�����Z��Z��Z�����������Z�����������DZZZZZZZZggZ�������Z������tDZZZZZZZZggZZZZZZZZZ{�}�{�bjhjcZwZjhjDZZZZZZZZggZ~�����tDZZZZZZZZggZZZZZZZZZ�Z��Z�{�DZZZZZZZZggZ����Z����������tDZZZZZZZZggZZZZZZZZZ����DZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZZ{|�b{�}�{�b�ccZvwZ�{����������lDZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZZ����DDZZZZ��������ZZ{�}�{�Zb�ZtZ��Z�{�uZ�ZtZ��Z�{�cZ������Z�{�uDZZZZZZZZggZ�������tDZZZZZZZZggZZZZZZZZZ�������Z���Z���������Z�����Z��Z���Z�����Z��Z�������Z��DZZZZZZZZggZZZZZZZZZ���Z�����Zb�fZ�cfZ�����Z��Z��Z�����������Z�����������DZZZZZZZZggZ�������Z������tDZZZZZZZZggZZZZZZZZZ{�}�{�bjhjfZ�cZwZjhjZ��Z�ZxZjhjDZZZZZZZZggZZZZZZZZZ{�}�{�bjhjfZ�cZwZ�{�����Z��Z�ZvZjhjDZZZZZZZZggZZZZZZZZZ{�}�{�b�fZjhjcZwZ�{����������lZ��Z�ZxZjhjDZZZZZZZZggZZZZZZZZZ{�}�{�b�fZjhjcZwZg�{����������lZ��Z�ZvZjhjDZZZZZZZZggZ~�����tDZZZZZZZZggZZZZZZZZZ�Z��Z�{�DZZZZZZZZggZZZZZZZZZ�Z��Z�{�fZ�ZiwZjhjZ����Z�ZwZjhjDZZZZZZZZggZ����Z����������tDZZZZZZZZggZZZZZZZZZ����Z��Z�ZwZjhjZ���Z�ZwZjhjDZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZZg�{�����ZvZ{�}�{�b�f�cZvwZ�{�����DZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZZ����DDZZZZ��������Z����Zb�ZtZ��Z�{�cZ������Z�{�uDZZZZZZZZggZ�������tDZZZZZZZZggZZZZZZZZZ�������Z����������Z����Z��Z�DZZZZZZZZggZ�������Z������tDZZZZZZZZggZZZZZZZZZ����bjhjcZwZjhjDZZZZZZZZggZ~�����tDZZZZZZZZggZZZZZZZZZ�Z��Z�{�DZZZZZZZZggZ����Z����������tDZZZZZZZZggZZZZZZZZZ����DZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZZ����b�cZ��Z��������������Z���������DZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZZ�cZ���Z������Z������Z��Z����Z��Z�������������Z�����Z��tDZZZZZZZZggZZZZZZZZZZZZZZZZ{|�b�cZvwZ���b�{�a����cDDDZZZZ��������Z}���Zb�ZtZ��Z�{�cZ������Z�{�uDZZZZZZZZggZ�������tDZZZZZZZZggZZZZZZZZZ�������Z����������Z������Z��Z�DZZZZZZZZggZ�������Z������tDZZZZZZZZggZZZZZZZZZ}���bjhjcZwZkhjDZZZZZZZZggZ~�����tDZZZZZZZZggZZZZZZZZZ�Z��Z�{�DZZZZZZZZggZ����Z����������tDZZZZZZZZggZZZZZZZZZ����DZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZZ}���b�cZxwZkhjDZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZZ�cZ���Z������Z������Z��Z}���Z��Z�������������Z�����Z��tDZZZZZZZZggZZZZZZZZZZZZZZZZ{|�b�cZvwZ���b�{�a����cDDZZZZ��������Z�{��Zb�ZtZ��Z�{�cZ������Z�{�uDZZZZZZZZggZ�������tDZZZZZZZZggZZZZZZZZZ�������Z����������Z�������Z��Z�DZZZZZZZZggZ�������Z������tDZZZZZZZZggZZZZZZZZZ�{��bjhjcZwZjhjDZZZZZZZZggZ~�����tDZZZZZZZZggZZZZZZZZZ�Z��Z�{�DZZZZZZZZggZ����Z����������tDZZZZZZZZggZZZZZZZZZ����DZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZZ{|�b�{��b�ccZvwZkhjDZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZZ����DDZZZZ��������Z{�}����Zb�ZtZ��Z�{�cZ������Z�{�uDZZZZZZZZggZ�������tDZZZZZZZZggZZZZZZZZZ�������Z�������Z����������Z����Z��Z�DZZZZZZZZggZ�������Z������tDZZZZZZZZggZZZZZZZZZ{�}����bjhjcZwZjhjDZZZZZZZZggZ~�����tDZZZZZZZZggZZZZZZZZZ�Z��Z�{�DZZZZZZZZggZ����Z����������tDZZZZZZZZggZZZZZZZZZ����DZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZZ{�}����b�cZ��Z��������������Z���������DZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZZ�cZ���Z���������Z�����Z��Z{�}����Z��Z�������������Z�����Z��tDZZZZZZZZggZZZZZZZZZZZZZZZZ{|�b{�}����b�ccZvwZ���b�{�a����cDDZZZZ��������Z{�}}���Zb�ZtZ��Z�{�cZ������Z�{�uDZZZZZZZZggZ�������tDZZZZZZZZggZZZZZZZZZ�������Z�������Z����������Z������Z��Z�DZZZZZZZZggZ�������Z������tDZZZZZZZZggZZZZZZZZZ{�}}���bkhjcZwZjhjDZZZZZZZZggZ~�����tDZZZZZZZZggZZZZZZZZZ�ZxwZkhjDZZZZZZZZggZ����Z����������tDZZZZZZZZggZZZZZZZZZ����Z��Z�ZvZkhjDZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZZ{�}}���b�cZxwZjhjDZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZZ�cZ���Z�����Z�����Z��Z���Z���������Z�����Z��Z{�}}���Z��DZZZZZZZZggZZZZZZZZZZZZ�������������Z�����Z��tZZZ{�}}���b�cZvwZ���b�{�a����cDDZZZZ��������Z{�}�{��Zb�ZtZ��Z�{�cZ������Z�{�uDZZZZZZZZggZ�������tDZZZZZZZZggZZZZZZZZZ�������Z�������Z����������Z�������Z��Z�DZZZZZZZZggZ�������Z������tDZZZZZZZZggZZZZZZZZZ{�}�{��bjhjcZwZjhjDZZZZZZZZggZ~�����tDZZZZZZZZggZZZZZZZZZ{|�b�cZvZkhjDZZZZZZZZggZ����Z����������tDZZZZZZZZggZZZZZZZZZ����Z��Z{|�b�cZxwZkhjDZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZZ{�}�{��b�cZ��Z��������������Z���������DZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZZ�cZ���Z���������Z�����Z��Z{�}�{��Z��Z�������������Z�����Z��tDZZZZZZZZggZZZZZZZZZZZZZZZZ{|�b{�}�{��b�ccZvZ���b�{�a����cDD���ZZ�{����{�uDDDDggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggDggDggZ}��������ZksspZ��Z�hZ{��Z������Z��������hDDggZ����Z������Z����Z��Z��Z�����������Z����Z��Z�Z���ZkjqphlgksspfZ�Z��������ZDggZ��~�Z������������Z��������hZ����Z������Z����Z���Z���Z��Z������fZ����fZ��ZDggZ��������Z����Z��������Z����Z��Z����Z�������Z�������Z����������Z����Z���Z�DggZ���������Z~���������hZ����Z������Z����Z���Z��Z����Z��Z���������Z����Z��������ZDggZ���Z���Z��Z�����������Z��Z��������Z����Z��Z���Z������Z��Z����Z��Z���ZDggZ��������Z����Z����Z���Z�����Z������Z�������������Z��Z���Z��������Z������Z����hDggZ����Z������Z����Z���Z��Z������Z���Z����������Z���Z�������Z��������Z�����hZDggZ����Z������Z����Z��Z��������Z��Z��Z{�Z��Z�����hZ���Z�Z���������Z{��ZDggZ�{��{���Z�����Z��Z�����~Z��}��~���Z{��Z�{��{���Z��Z��}�{��{|�����ZDggZ{�~Z������Z���Z��Z���Z{Z�{���}��{�Z������hZ���Z����Z��Z���Z������ZDggZ����Z�����Z���������Z���Z����Z�Z��������Z����Z���Z�������Z��Z���������ZDggZ�������Z���Z��Z���Z���Z�������hDDggDggZ�����tZZZZZZZ��������Z��~�Z������������Z��������Zb�Z���ZkjqphlgksspfDggZZZZZZZZZZZZZZ�{����{�cDggDggZ�������tZZZZZ����Z�������Z�����Z��Z��������Z����Z�Z�������DggZZZZZZZZZZZZZZ������������Z�����Z�hDggDggZ~���������tZZ�Z~{�}Z��~�Z������������Z��������Z�������Z�����DggDggZ�������tZZZZZ����Z�������Z����Z��Z�Z������������Z��������������Z��Z���ZDggZZZZZZZZZZZZZZ�������������Z�������Z��Z���Z�{����{�Z�������Z�����������hDggDggZ����������tZZ���Z������Z���������Z��Z���Z���������Z��Z����Z�������Z���DggZZZZZZZZZZZZZZ����Z����Z��������Z��Z��������fZ���Z���Z���������Z��Z�������DggZZZZZZZZZZZZZZ��Z����Z����������Z��Z��Z���Z�������Z��������Z��Z�Z���ZkjqpDggZZZZZZZZZZZZZZgkssmhDggDggZ�����tDggZZZZZZZZZZZZZZ���Z\�������Z�����������\Z�������Z���Z�����fZ��������fZ���DggZZZZZZZZZZZZZZ������������Z��Z�{����{�hDggZZZZZZZZZZZZZZ���Z��������Z������������Z����������Z���Z������������Z�������DggZZZZZZZZZZZZZZ��Z���Z������������Z���������Z����Z���Z����Z��Z����Z��������DggZZZZZZZZZZZZZZ���������Z���Z������Z���������Z��Z���Z��������������Z��Z���DggZZZZZZZZZZZZZZ�{����{�Z�������Z�����������hZZ���Z�������Z��Z���Z�{����{�DggZZZZZZZZZZZZZZ�������Z����Z��Z��Z�������Z����Z���������Z���Z�������Z�DggZZZZZZZZZZZZZZ���������Z���Z���������������Z��Z������Z�����Z��������������DggZZZZZZZZZZZZZZ��Z�{����{�hZZ����Z����������Z���Z������Z��Z���������DggZZZZZZZZZZZZZZ���Z�������Z����Z��Z���Z����Z���������Z������Z���������Z��Z����hDggDggZgggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggDggZ�������ZZZZtZkhoDggZ~���ZZZZZZZtZlnZ����ZksspDggZgggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggDD�������Z����Z�{����{�Z��DDZZZZggDZZZZggZ�����Z}��������Z���Z���Z��Z���Z�������Z|���Z����DZZZZggDZZZZ��������ZZ�{�����lZtZZ�{�ZtwZqhmrsjo�pjsrs�mjpojuZZZggZ�ddlDZZZZ��������ZZ�{�����kjZtZZ�{�ZtwZlljlphnpoqs�nrjpq�kquZggZ�ddkjDZZZZ��������ZZ�{����������ZtZ�{�ZtwZlohkmlqn�kllrq�krmno�sjqqj�kkouZggrd��DZZZZ��������ZZ�{�����tZZ�����ZtwZlquZZggZ�������Z���������Z������Z���Z������DZZZZ��������ZZ�{��}����tZ�����ZtwZkojuZggZ�������Z�����Z���Z������Z��Z�����DZZZZ��������ZZ|{����tZ�{�ZtwZjhjjjjkuZZggZ������Z���Z�����������Z��������DZZZZ��������ZZ�}ZtZ�{�ZtwZphjqlolsmojjrrrknl�gjkuZggZ}�������Z���Z������DDZZZZggDZZZZggZ�����Z����Z~�����������Z���Z}�����Z����������DZZZZggDZZZZ����Z�{���}���Z��Z�����Zb�{���{�Z�����ZvxcZ��Z�{�uDZZZZ����Z�{���{���}���Z��Z�����Zb�{���{�Z�����ZvxcZ��Z�{���{�uDZZZZ�������Z�{���}�����Z��Z�{���}���ZbjZ��Z�{�����cuDZZZZ�������Z�{��{���lZ��Z�{���}���ZbjZ��ZkcuDZZZZ�������Z�{��{���mZ��Z�{���}���ZbjZ��ZlcuDZZZZ�������Z��{~�{��Z��Z�����Z�����ZjZ��ZmuDZZZZ����Z}��~�}���~����Z��Zb���{����fZ�}������cuDDZZZZggDZZZZggZ{��������Z���������Z���Z}�����Z{���������DZZZZggDZZZZ��������Z��������l�����Zb~ZtZ��Z�{���{���}���uZ�����{���{��ZtZ��Z�{�uDZZZZZZZZZZZZZZZZ���|������{���ZtZ��Z�{���{�cZ������Z�{���}���Z��DZZZZZZZZggZ~����������tDZZZZZZZZggZZZZZZZZ�������Z�����Z��Z���Z���Z�Z������Z��Z������DZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZ����DZZZZZZZZggDZZZZZZZZ��������Z�ZtZ�{���}���ZbjZ��Z���|������{���cuDZZZZZZZZ��������Z���ZtZ�{�ZtwZ�����{���{��uDZZZZZZZZ��������Z��{�ZtZ|���{�ZtwZ���uDZZZZ�����DZZZZZZZZZZZZZZ���Z�Z��ZjZ��Z���|������{���Z����DZZZZZZZZZZZZZZZZZ�b�cZtwZ���uDZZZZZZZZZZZZZZZZZ���Z�Z��Z~a�{��Z����DZZZZZZZZZZZZZZZZZZZZZZZZZZZZ��Z�ZwZ~b�cZ����DZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ��{�ZtwZ�{��uDZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ����uDZZZZZZZZZZZZZZZZZZZZZZZZZZZZ���Z��uDZZZZZZZZZZZZZZZZZ���Z����uDZZZZZZZZZZZZZZZZZ��Z��{�Z����DZZZZZZZZZZZZZZZZZZZZZZZZZZZZ���ZtwZ���ilhjuDZZZZZZZZZZZZZZZZZ���Z��uDZZZZZZZZZZZZZZZZZ��{�ZtwZ���uDZZZZZZZZZZZZZZ���Z����uDZZZZZZZZZZZZZZ������Z�uDZZZZ���Z��������l�����uDDDZZZZ��������Z����{�������ZtZ�{���}���ZtwZ��������l�����bDZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ�{���{���}���abkjjfZsjcfkhjfDZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ�{�����cuDDZZZZ��������Z������ZtZ�{���}�����ZtwZbDZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZqhromsrkpmmsqnnrlq�gjkfDZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZnhpmpnqpjsjjjrjpjp�gjkfDZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZlhnnsqrppmklprpnkm�gjkfDZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZkhlnmonssnonpqpknn�gjkfDZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZphlnkrrjsssosoqmok�gjlfDZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZmhklmsrmmnmjlprlqq�gjlfDZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZkhoplmqlrpljnqprmj�gjlfDZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZqhrklmnkjpjkjkkkkp�gjmfDZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZmhsjplmjkmksppsqkq�gjmfDZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZkhsomkllokpnqrrkrs�gjmfDZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZshqpoplkrsoosmksmq�gjnfDZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZnhrrlrklkkksnrsrls�gjnfDZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZlhnnknjpljknsmpkqo�gjnfDZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZkhlljqjmkkrsmpqjlk�gjnfDZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZphkjmokopkqnljrqpr�gjofDZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZmhjokqoqrkkoolpjsm�gjofDZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZkholorqrsjpkmkoqpj�gjofDZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZqhplsmsnomkkjkspss�gjpfDZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZmhrknpsqlpopjpnspj�gjpfDZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZkhsjqmnrpmlrkjkrqj�gjpfDZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZshompqnmkpnjospjrj�gjqfDZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZnhqprmqkorljmjrrqp�gjqfDZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZlhmrnkroqskjkoorjk�gjqfDZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZkhksljslrsoojqrjpq�gjqfDZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZohspjnpnnqqomsjoom�gjrfDZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZlhsrjlmllmrqpsomjm�gjrfDZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZkhnsjkkpkksmrnqpon�gjrfDZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZqhnojorjospslmrlrk�gjsDZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZcuDDZZZZ��������Z}��~�}ZbZ�jZtZ��Z�{�uDZZZZZZZZZZZZZZZZZZZZZZ�jZtZ��Z�{�uDZZZZZZZZZZZZZZZZZZZZZZ�jZtZ��Z�{�uDZZZZZZZZZZZZZZZZZZZZZZ�ZtZ��Z�{���{�uZZZZZZZZZZZZZZZZZggZZ���������Z������DZZZZZZZZZZZZ}��~�}���~ZtZ��Z}��~�}���~����ZZZZZZZZZggZZ��������Zb�ZgxZjcDZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZggZZ��Z���������Zb�ZgxZjcDZZZZZZZZZZZZZZZZZZZZcZ������Z�{��{���mZ��DZZZZZZZZggZ~����������tDZZZZZZZZggZZZZZZZZ}������Z������Z������DZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZZ����DZZZZZZZZZZZZZ��������Z�ZtZ�{�ZtwZ�juDZZZZZZZZZZZZZ��������Z�ZtZ�{�ZtwZ�juDZZZZZZZZZZZZZ��������Z�ZtZ�{�ZtwZ�juDZZZZZZZZZZZZZ��������Z�����ZtZ�{�uDZZZZ�����DZZZZZZZ��Z}��~�}���~ZwZ���{����Z����DZZZZZZZZZZZ���Z�Z��ZjZ��Z�Z����DZZZZZZZZZZZZZZZZZZZZZZ�����ZtwZ�uDZZZZZZZZZZZZZZZZZZZZZZ��ZbZ�ZxwZjhjcZ����DZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ�ZtwZ�ZgZ�ZdZ����{�������b�cuDZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ�ZtwZ�ZeZ�����ZdZ����{�������b�cuDZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ�ZtwZ�ZgZ������b�cuDZZZZZZZZZZZZZZZZZZZZZZ����DZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ�ZtwZ�ZeZ�ZdZ����{�������b�cuDZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ�ZtwZ�ZgZ�����ZdZ����{�������b�cuDZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ�ZtwZ�ZeZ������b�cuDZZZZZZZZZZZZZZZZZZZZZZ���Z��uDZZZZZZZZZZZZ���Z����uDZZZZZZZZ����DZZZZZZZZZZZZ���Z�Z��ZjZ��Z�Z����DZZZZZZZZZZZZZZZZZZZZ�����ZtwZ�uDZZZZZZZZZZZZZZZZZZZZ��ZbZ�ZvZjhjcZ����DZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ�ZtwZ�ZgZ�ZdZ����{�������b�cuDZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ�ZtwZ�ZeZ�����ZdZ����{�������b�cuDZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ�ZtwZ�ZgZ������b�cuDZZZZZZZZZZZZZZZZZZZZ����DZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ�ZtwZ�ZeZ�ZdZ����{�������b�cuDZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ�ZtwZ�ZgZ�����ZdZ����{�������b�cuDZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ�ZtwZ�ZeZ������b�cuDZZZZZZZZZZZZZZZZZZZZ���Z��uDZZZZZZZZZZZZ���Z����uDZZZZZZZZ���Z��uDZZZZZZZZ������Z�{��{���mab�fZ�fZ�cuDZZZZ���Z}��~�}uDDZZZZggDZZZZggZ|�����Z���Z������Z������������Z���������Z�����Z����DZZZZggDZZZZ��������Z����Zb�tZ��Z�{�ZcZ������Z�{�Z��DZZZZZZZZggZ~����������tDZZZZZZZZggZZZZZZZZ���Z��������Z�����������Z��Z�Z���ZkjqphlgksspDZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZ����DZZZZ�����DZZZZZZZZZZZ��ZZbZ�ZxZjhjZcZZ����DZZZZZZZZZZZZZZZZ������ZkhjuDZZZZZZZZZZZ�����ZbZ�ZvZjhjZcZZ����DZZZZZZZZZZZZZZZZ������ZgkhjuDZZZZZZZZZZZ����DZZZZZZZZZZZZZZZZ������ZjhjuDZZZZZZZZZZZ���Z��uDZZZZ���Z����uDDZZZZ��������Z}��Zb�ZtZ��Z�{�ZcZ������Z�{�Z��DZZZZZZZZggZ~����������tDZZZZZZZZggZZZZZZZZ���Z��������Z�����������Z��Z�Z���ZkjqphlgksspDZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZ�cZ��Z����������Z��Z��Z�����Z����Z��Z��������fZ��Z��������DZZZZZZZZggZZZZZZZZZZZ������Z��������Z���Z�����Z���������DZZZZZZZZggZZZZZZZZ�cZ���Z������Z���������Z��Z����Z��������Z��Z�ZvwZ�{��DZZZZZZZZggZZZZZZZZ�cZ�������Z�Z��Z{|�b�cZxwZ�{��DDZZZZZZZZ��������Z�{��tZ�{�ZZtwZ�{�b�����a����cuDZZZZZZZZ��������Z�~tZ�{�uDDZZZZ�����DZZZZZZZZZ��Z{|�b�cZxwZ�{��Z����DZZZZZZZZZZZZZZZ������Z�uDZZZZZZZZZ���Z��uDDZZZZZZZZZ�~ZtwZ�{�ZbZ�����b�ccuDZZZZZZZZZ��Z�~ZwZ�Z����DZZZZZZZZZZZZ������Z�uDZZZZZZZZZ���Z��uDDZZZZZZZZZZZZ��Z�ZxZjhjZ����DZZZZZZZZZZZZZZZZZZZZZZZ��Z�~ZxwZ�Z����DZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ������Z�~uDZZZZZZZZZZZZZZZZZZZZZZZ����DZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ������Z�~ZeZkhjuDZZZZZZZZZZZZZZZZZZZZZZZ���Z��uDZZZZZZZZZZZZ�����ZZ�ZwZjhjZZ����DZZZZZZZZZZZZZZZZ������ZjhjuDZZZZZZZZZZZZ����DZZZZZZZZZZZZZZZZZZZZZZZ��Z�~ZvwZ�Z����DZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ������Z�~ZeZkhjuDZZZZZZZZZZZZZZZZZZZZZZZ����DZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ������Z�~uDZZZZZZZZZZZZZZZZZZZZZZZ���Z��uDZZZZZZZZZZZZ���Z��uDZZZZ���Z}��uDDZZZZ��������Z�����Zb�ZtZ��Z�{�ZcZ������Z�{�Z��DZZZZZZZZggZ~����������tDZZZZZZZZggZZZZZZZZ���Z��������Z�����������Z��Z�Z���ZkjqphlgksspDZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZ�cZ��Z����������Z��Z��Z�����Z����Z��Z��������fZ��Z��������DZZZZZZZZggZZZZZZZZZZZ������Z��������Z���Z�����Z���������DZZZZZZZZggZZZZZZZZ�cZ���Z������Z���������Z��Z����Z��������Z��Z{|�b�cZvwZ�{��DZZZZZZZZggZZZZZZZZ�cZ�������Z�Z��Z{|�b�cZxwZ�{��DDZZZZZZZZ��������Z�{��tZ�{�ZZtwZ�{�b�����a����cuDZZZZZZZZ��������Z�~tZ�{�uDDZZZZ�����DZZZZZZZZ��Z{|�bZ�ZcZxwZ�{��Z����DZZZZZZZZZZZZZZZZZZZZ������Z�uDZZZZZZZZ���Z��uDDZZZZZZZZ�~ZtwZ�{�ZbZ�����b�ccuDZZZZZZZZ��Z�~ZwZ�Z����DZZZZZZZZZZZZZZZZ������Z�uDZZZZZZZZ���Z��uDDZZZZZZZZ��Z�ZxZjhjZ����DZZZZZZZZZZZZZZZZZZZZZZ��Z�~ZvwZ�Z����DZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ������Z�~uDZZZZZZZZZZZZZZZZZZZZZZZ����DZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ������Z�~ZgZkhjuDZZZZZZZZZZZZZZZZZZZZZZZ���Z��uDZZZZZZZZ�����ZZ�ZwZjhjZZ����DZZZZZZZZZZZZZZZZ������ZjhjuDZZZZZZZZ����DZZZZZZZZZZZZZZZZZZZ��Z�~ZxwZ�Z����DZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ������Z�~ZgZkhjuDZZZZZZZZZZZZZZZZZZZ����DZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ������Z�~uDZZZZZZZZZZZZZZZZZZZ���Z��uDZZZZZZZZ���Z��uDZZZZ���Z�����uDDZZZZ��������Z����~Zb�ZtZ��Z�{�ZcZ������Z�{�Z��DZZZZZZZZggZ~����������tDZZZZZZZZggZZZZZZZZ���Z��������Z�����������Z��Z�Z���ZkjqphlgksspDZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZZ�cZ�������ZjhjZ��Z�ZwZjhjDZZZZZZZZggZZZZZZZZZ�cZ�������Z�����b�ZeZjhocZ��Z�ZxZjDZZZZZZZZggZZZZZZZZZ�cZ�������Z}��b�ZgZjhocZ��Z�ZvZjDDZZZZ�����DZZZZZZZZZZZ��ZZ�ZxZjhjZZ����DZZZZZZZZZZZZZZZZ������Z�����b�ZeZjhocuDZZZZZZZZZZZ�����ZZ�ZvZjhjZZ����DZZZZZZZZZZZZZZZZ������Z}��bZ�ZgZjhocuDZZZZZZZZZZZ����DZZZZZZZZZZZZZZZZ������ZjhjuDZZZZZZZZZZZ���Z��uDZZZZ���Z����~uDDZZZZ��������Z����}Zb�ZtZ��Z�{�ZcZ������Z�{�Z��DZZZZZZZZggZ~����������tDZZZZZZZZggZZZZZZZZ���Z��������Z�����������Z��Z�Z���ZkjqphlgksspDZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZZ�cZ�������ZjhjZ��Z�ZwZjhjDZZZZZZZZggZZZZZZZZZ�cZ�������Z�����b�cZ��Z�ZxZjDZZZZZZZZggZZZZZZZZZ�cZ�������Z}��b�cZ��Z�ZvZjDDZZZZ�����DZZZZZZZZZZZ��ZZ�ZxZjhjZZ����DZZZZZZZZZZZZZZZZ������Z�����b�cuDZZZZZZZZZZZ�����ZZ�ZvZjhjZZ����DZZZZZZZZZZZZZZZZ������Z}��bZ�cuDZZZZZZZZZZZ����DZZZZZZZZZZZZZZZZ������ZjhjuDZZZZZZZZZZZ���Z��uDZZZZ���Z����}uDDDDDZZZZ��������Z\��~\Zb�fZ�tZ��Z�{�ZcZ������Z�{�Z��DZZZZZZZZggZ~����������tDZZZZZZZZggZZZZZZZZ���Z��������Z�����������Z��Z�Z���ZkjqphlgksspDZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZ�cZ�������ZjhjZ��Z�����DDZZZZZZZZ��������Z���{���ZtZ|���{�ZtwZ�ZvZjhjuDZZZZZZZZ��������Z���{���ZtZ|���{�ZtwZ�ZvZjhjuDZZZZZZZZ��������Z�{��ZtZ�{�uDZZZZ�����DZZZZZZZZggZ}����Z��������Z��Z�����Z���������DZZZZZZZZZZZZ��Zb�ZwZjhjcZ����DZZZZZZZZZZZZZZZZZ������Z�{��DZZZZZZZZZZZZZZZZZZZZZZZZ������Z\��~b�fZjhjcZ��Z���������\DZZZZZZZZZZZZZZZZZZZZZZZZ��������Z����uDZZZZZZZZZZZZZZZZZ������ZjhjuDZZZZZZZZZZZZZZ���Z��uDDZZZZZZZZggZ}������Z�����DZZZZZZZZ��ZbZ���{���ZcZ����DZZZZZZZZZZZZZZZZ��ZbZ���{���ZcZ����DZZZZZZZZZZZZZZZZZZZZZZZZ�{��ZtwZ�ZeZb�����b{|�b�ci{|�b�cccd{|�b�cuDZZZZZZZZZZZZZZZZ����DZZZZZZZZZZZZZZZZZZZZZZZZ�{��ZtwZ�ZeZb}��b{|�b�ci{|�b�cccd{|�b�cuDZZZZZZZZZZZZZZZZ���Z��uDZZZZZZZZ����DZZZZZZZZZZZZZZZZ��ZbZ���{���ZcZ����DZZZZZZZZZZZZZZZZZZZZZZZZ�{��ZtwZ�ZgZb}��b{|�b�ci{|�b�cccd{|�b�cuDZZZZZZZZZZZZZZZZ����DZZZZZZZZZZZZZZZZZZZZZZZZ�{��ZtwZ�ZgZb�����b{|�b�ci{|�b�cccd{|�b�cuDZZZZZZZZZZZZZZZZ���Z��uDZZZZZZZZ���Z��uDDZZZZZZZZ������Z�{��uDZZZZ���Z\��~\uDDDZZZZ��������Z�{��{�Zb�fZ�ZtZ��Z�{�ZcZ������Z�{�Z��DZZZZZZZZggZ~����������tDZZZZZZZZggZZZZZZZZ���Z��������Z�����������Z��Z�Z���ZkjqphlgksspDZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZ�cZ�{��{�b�f�cZwZ�Z����Z�ZwZ�DZZZZZZZZggDZZZZ�����DZZZZZZZZ��Z�ZxwZ�Z����DZZZZZZZZZZZ������Z�uDZZZZZZZZ����DZZZZZZZZZZZ������Z�uDZZZZZZZZ���Z��uDZZZZ���Z�{��{�uDDZZZZ��������Z�{����Zb�fZ�ZtZ��Z�{�ZcZ������Z�{�Z��DZZZZZZZZggZ~����������tDZZZZZZZZggZZZZZZZZ���Z��������Z�����������Z��Z�Z���ZkjqphlgksspDZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZ�cZ�{����b�f�cZwZ�Z����Z�ZwZ�DZZZZZZZZggDZZZZ�����DZZZZZZZZ��Z�ZvwZ�Z����DZZZZZZZZZZZ������Z�uDZZZZZZZZ����DZZZZZZZZZZZ������Z�uDZZZZZZZZ���Z��uDZZZZ���Z�{����uDDDZZZZ���������Z�������b��������Z�~kf�~lt�����Z�������u��������Z�t���Z�{�cDZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ��DZZZZZZZZggZ~����������tDZZZZZZZZggZZZZZZZZ���Z��������Z�����������Z��Z�Z���ZkjqphlgksspDZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZ�cZ�������ZjhjZ��Z�����DZZZZZZZZggDZZZZZZZZ��������Z�fZ�tZ�����uDZZZZZZZZ��������Z��~kZtZ�����ZtwZ�����ab�~kcuDZZZZZZZZ��������Z��~lZtZ�����ZtwZ�����ab�~lcuDZZZZ�����DZZZZZZZZggZ}����Z��������Z��Z���������DZZZZZZZZ��Z�~kZxZlknqnrmoplZ����DZZZZZZZZZZZZZZZZ������Z�{��DZZZZZZZZZZZZZZZZZZZZZZZZ������Z\�~kZxZlknqnrmoplZ��Z�������\DZZZZZZZZZZZZZZZZZZZZZZZZ��������Z����uDZZZZZZZZZZZZZZZZ�ZtwZjhjuDZZZZZZZZZZZZZZZZ������uDZZZZZZZZ���Z��uDDZZZZZZZZ��Z�~lZxZlknqnrmmsrZ����DZZZZZZZZZZZZZZZZ������Z�{��DZZZZZZZZZZZZZZZZZZZZZZZZ������Z\�~lZxZlknqnrmmsrZ��Z�������\DZZZZZZZZZZZZZZZZZZZZZZZZ��������Z����uDZZZZZZZZZZZZZZZZ�ZtwZjhjuDZZZZZZZZZZZZZZZZ������uDZZZZZZZZ���Z��uDDZZZZZZZZggZ}������Z���Z����Z������Z���Z������g������Z������DZZZZZZZZ�ZtwZ��~kiomppruDZZZZZZZZ��~kZtwZnjjknZdZb��~kZgZ�ZdZompprcZgZ�ZdZkllkkuDDZZZZZZZZ��Z��~kZvZjZZ����DZZZZZZZZZZZZZZZZ��~kZtwZ��~kZeZlknqnrmopmuDZZZZZZZZ���Z��uDDZZZZZZZZ�ZtwZ��~liolqqnuDZZZZZZZZ��~lZtwZnjpslZdZb��~lZgZ�ZdZolqqncZgZ�ZdZmqskuDDZZZZZZZZ��Z��~lZvZjZZ����DZZZZZZZZZZZZZZZZ��~lZtwZ��~lZeZlknqnrmmssuDZZZZZZZZ���Z��uDDZZZZZZZZ�ZtwZ��~kZgZ��~luDZZZZZZZZ��Z�ZvZkZ����DZZZZZZZZZZZZZZZZ�ZtwZ�ZeZlknqnrmopluDZZZZZZZZ���Z��uDDZZZZZZZZggZ���Z������Z������DZZZZZZZZ�~kZtwZ�������ab��~kcuDZZZZZZZZ�~lZtwZ�������ab��~lcuDZZZZZZZZ�ZtwZZ�{�b�cdnhpoppkm�gkjuDZZZZ���Z�������uDDDDZZZZ��������Z����Zb�ZtZ��Z�{�ZcZ������Z�{�Z��DZZZZZZZZggZ~����������tDZZZZZZZZggZZZZZZZZ���Z��������Z�����������Z��Z�Z���ZkjqphlgksspDZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZ�cZ����Z���Z������g�������Z�������������tDZZZZZZZZggZZZZZZZZZZZZ�b�ekcZwZjhod��b�cZeZ�i�b�c�DZZZZZZZZggZZZZZZZZ�cZ�������ZjhjZ��Z�����DZZZZZZZZggDDZZZZZZZZ��������Z��ZtZ�{�ZtwZ|{����d|{����uZggZ}����������Z������DDZZZZZZZZ��������Z����{�tZ�{�uDZZZZZZZZ��������Z��~�{�ZtZ�{�ZuDZZZZZZZZ��������Z���{�ZtZ�{�ZuDZZZZZZZZ��������Z}����ZtZ�����ZtwZkuDDZZZZ�����DZZZZZZZZggZ}����Z��������Z��Z��������DZZZZZZZZ��ZbZ�ZvZjhjZcZ����DZZZZZZZZZZZZZZZZ������Z�{��DZZZZZZZZZZZZZZZZZZZZZZZZ������Z\�ZvZjhjZ��Z����b�c\DZZZZZZZZZZZZZZZZZZZZZZZZ��������Z����uDZZZZZZZZZZZZZZZZ������ZjhjuDZZZZZZZZ���Z��uDDZZZZZZZZggZ���Z���Z������Z����Z���Z�������Z�����DZZZZZZZZ��Z�ZwZjhjZ����DZZZZZZZZZZZZZZZZZZ������ZjhjuDZZZZZZZZ����DZZZZZZZZZZZZZZZZ��ZbZ�ZwZkhjZcZ����DZZZZZZZZZZZZZZZZZZZZZZZZ������ZkhjuDZZZZZZZZZZZZZZZZ���Z��uDZZZZZZZZ���Z��uDDZZZZZZZZggZ���Z���Z������Z����Z���Z�������Z�����DZZZZZZZZ����{�ZtwZ��b���b�cdbjhoccuZggZ��������������Z�������Z���Z���������DZZZZZZZZ��~�{�ZtwZ����{�uDZZZZZZZZ���{�ZtwZb�i��~�{�ZeZ��~�{�cdjhouDDZZZZZZZZggZ}����Z���ZZ��������Z���Z��������Z�����Z���Z���Z�����DZZZZZZZZ�����ZZbZbZb{|�bb���{�Zg��~�{�ci���{�cZxZ��cZ��DZZZZZZZZZZZZZZZZZZZb{|�b���{�ZgZ��~�{�cZxZ��cZcZ{�~DZZZZZZZZZZZZZZZZZZZb}����ZvZ�{��}����cZcZZ����DZZZZZZZZZZZZZZZZ��~�{�ZtwZ���{�uDZZZZZZZZZZZZZZZZ���{�ZtwZb�i��~�{�ZeZ��~�{�cdjhouDZZZZZZZZZZZZZZZZ}����ZtwZ}����ZeZkuDZZZZZZZZ���Z����uDZZZZZZZZ������Z���{�uDZZZZ���Z����uDDZZZZ��������Z}|��Zb�ZtZ��Z�{�ZcZ������Z�{�Z��DZZZZZZZZggZ~����������tDZZZZZZZZggZZZZZZZZ���Z��������Z�����������Z��Z�Z���ZkjqphlgksspDZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZ�cZ����Z���Z������g�������Z�������������tDZZZZZZZZggZZZZZZZZZZZZ�b�ekcZwZbkimcd�ld�b�cZeZ�i�b�cddl�uDZZZZZZZZggDZZZZZZZZ��������Z��ZtZ�{�ZtwZ|{����d|{����uDDZZZZZZZZ��������Z����{�tZ�{�uDZZZZZZZZ��������Z���}{�ZtZ�{�ZtwZ�uDZZZZZZZZ��������Z��{���ZtZ|���{�ZtwZ�ZvZjhjuDZZZZZZZZ��������Z��~�{�ZtZ�{�ZuDZZZZZZZZ��������Z���{�ZtZ�{�ZuDZZZZZZZZ��������Z}����ZtZ�����ZtwZkuDDZZZZ�����DDZZZZZZZZggZ}������Z����Z���Z�������Z�����DZZZZZZZZ��Z�ZwZjhjZ����DZZZZZZZZZZZZZZZZ������ZjhjuDZZZZZZZZ�����ZbZ�ZwZkhjZcZ����DZZZZZZZZZZZZZZZZ������ZkhjuDZZZZZZZZ����DZZZZZZZZZZZZZZZZ��Z�ZwZgkhjZ����DZZZZZZZZZZZZZZZZZZZZZZZZ������ZgkhjuDZZZZZZZZZZZZZZZZ���Z��uDZZZZZZZZ���Z��uDDZZZZZZZZggZ}������Z����Z���Z�������Z�����DZZZZZZZZ��Z��{���Z����DZZZZZZZZZZZZZZZZ���}{�ZtwZg�uDZZZZZZZZ���Z��uDDZZZZZZZZ����{�ZtwZ��b���b���}{�cibmhjccuZggZ��������������Z�������Z���DZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZggZ���������DZZZZZZZZ��~�{�ZtwZ����{�uDZZZZZZZZ���{�ZtwZb���}{�ib��~�{�d��~�{�cZeZlhjd��~�{�cimhjuDDZZZZZZZZggZ}����Z���Z��������Z���Z��������Z������Z���Z���Z�����DZZZZZZZZ�����ZbZbZZb{|�bb���{�Zg��~�{�ci���{�cZxZ��ZcZ��DZZZZZZZZZZZZZZZZZZZb{|�b���{�ZgZ��~�{�cZxZ��ZcZcZZ{�~DZZZZZZZZZZZZZZZZZZZbZ}����ZvZ�{��}����ZcZcZ����DZZZZZZZZZZZZZZZZ��~�{�ZtwZ���{�uDZZZZZZZZZZZZZZZZ���{�Ztwb���}{�ib��~�{�d��~�{�cZeZlhjd��~�{�cimhjuDZZZZZZZZZZZZZZZZ}����ZtwZ}����ZeZkuDZZZZZZZZ���Z����uDDZZZZZZZZ��Z��{���Z����DZZZZZZZZZZZZZZZZ���{�ZtwZg���{�uDZZZZZZZZ���Z��uDDZZZZZZZZ������Z���{�uDZZZZ���Z}|��uDDZZZZ��������Z\dd\Zb�ZtZ��Z�����uZ�ZtZ��Z�{�cZ������Z�{�Z��DZZZZZZZZggZ~����������tDZZZZZZZZggZZZZZZZZ���Z��������Z�����������Z��Z�Z���ZkjqphlgksspDZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZ�cZ�������ZjhjZ��Z�����Z���������DDZZZZ�����DZZZZZZZZggZ}����Z��������Z��Z��������DZZZZZZZZ��ZbZbZ�ZvZjZZcZ���ZbZ�ZiwZjhjZcZcZ����DZZZZZZZZZZZZZZZZ������Z�{��DZZZZZZZZZZZZZZZZZZZZZZZZ������Z\�ZvZjZ���Z�ZiwZjhjZ��Z�dd�\DZZZZZZZZZZZZZZZZZZZZZZZZ��������Z����uDZZZZZZZZZZZZZZZZ������ZjhjuDZZZZZZZZ���Z��uDDZZZZZZZZ��ZbZbZ�ZwZjZZcZ���ZbZ�ZvwZjhjZcZcZ����DZZZZZZZZZZZZZZZZ������Z�{��DZZZZZZZZZZZZZZZZZZZZZZZZ������Z\�ZwZjZ���Z�ZvwZjhjZ��Z�dd�\DZZZZZZZZZZZZZZZZZZZZZZZZ��������Z����uDZZZZZZZZZZZZZZZZ������ZjhjuDZZZZZZZZ���Z��uDDZZZZZZZZggZ���Z�����Z���Z�������Z�����DZZZZZZZZ��ZbZ�ZwZjZZ���ZZ�ZxZjhjZcZ����DZZZZZZZZZZZZZZZZ������ZjhjuDZZZZZZZZ���Z��uDDZZZZZZZZ��ZbZ�ZwZkZcZ����DZZZZZZZZZZZZZZZZ������ZkhjuDZZZZZZZZ���Z��uDDZZZZZZZZ��ZbZ�ZwZjhjZ���Z�ZiwZjZcZ����DZZZZZZZZZZZZZZZZ������ZkhjuDZZZZZZZZ���Z��uDDZZZZZZZZ��ZbZ�ZwZkhjcZ����DZZZZZZZZZZZZZZZZ������Zb�{�b�ccuDZZZZZZZZ���Z��uDDZZZZZZZZggZ���Z�����Z���Z�������Z����DZZZZZZZZ������Z��Zb�ZdZ���Zb�{�b�cccuDZZZZ���Z\dd\uDDZZZZ��������Z\dd\Zb�ZtZ��Z�{�uZ�ZtZ��Z�{�cZ������Z�{�Z��DZZZZZZZZggZ~����������tDZZZZZZZZggZZZZZZZZ���Z��������Z�����������Z��Z�Z���ZkjqphlgksspDZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZ�cZ�������ZjhjZ��Z�����Z���������DDZZZZ�����DZZZZZZZZggZ}����Z��������Z��Z��������DZZZZZZZZ��ZbZbZ�ZvZjhjZZcZ���ZbZ�ZiwZjhjZcZcZ����DZZZZZZZZZZZZZZZZ������Z�{��DZZZZZZZZZZZZZZZZZZZZZZZZ������Z\�ZvZjhjZ���Z�ZiwZjhjZ��Z�dd�\DZZZZZZZZZZZZZZZZZZZZZZZZ��������Z����uDZZZZZZZZZZZZZZZZ������ZjhjuDZZZZZZZZ���Z��uDDZZZZZZZZ��ZbZbZ�ZwZjhjZZcZ���ZbZ�ZvwZjhjZcZcZ����DZZZZZZZZZZZZZZZZ������Z�{��DZZZZZZZZZZZZZZZZZZZZZZZZ������Z\�ZwZjhjZ���Z�ZvwZjhjZ��Z�dd�\DZZZZZZZZZZZZZZZZZZZZZZZZ��������Z����uDZZZZZZZZZZZZZZZZ������ZjhjuDZZZZZZZZ���Z��uDDZZZZZZZZggZ���Z�����Z���Z�������Z�����DZZZZZZZZ��ZbZ�ZwZjhjZZ���ZZ�ZxZjhjZcZ����DZZZZZZZZZZZZZZZZ������ZjhjuDZZZZZZZZ���Z��uDDZZZZZZZZ��ZbZ�ZwZkhjZcZ����DZZZZZZZZZZZZZZZZ������ZkhjuDZZZZZZZZ���Z��uDDZZZZZZZZ��ZbZ�ZwZjhjZ���Z�ZiwZjhjZcZ����DZZZZZZZZZZZZZZZZ������ZkhjuDZZZZZZZZ���Z��uDDZZZZZZZZ��ZbZ�ZwZkhjcZ����DZZZZZZZZZZZZZZZZ������Zb�cuDZZZZZZZZ���Z��uDDZZZZZZZZggZ���Z�����Z���Z�������Z����DZZZZZZZZ������Z��Zb�ZdZ���Zb�ccuDZZZZ���Z\dd\uDDZZZZ��������Z��ZZb�ZtZ��Z�{�ZcZ������Z�{�Z��DZZZZZZZZggZ~����������tDZZZZZZZZggZZZZZZZZ���Z��������Z�����������Z��Z�Z���ZkjqphlgksspDZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZ�cZ����Z��������Z��������Z���Z�����������Z�����Z���Z���������DZZZZZZZZggZZZZZZZZZZZ������tDZZZZZZZZggZZZZZZZZZZZZZZZZ���b�cZwZkZeZ�ZeZ�ddlil[ZeZ�ddmim[ZeZhhhZuZ���ZvZkhjDZZZZZZZZggZZZZZZZZZZZ���Z�������Z��������Z�Z��Z����Z���������Z��Z���b�e�cZwDZZZZZZZZggZZZZZZZZZZZ���b�cd���b�cDZZZZZZZZggDZZZZZZZZggZZZZZZZZ�cZ����Z��������������Z������Z�Z��Z��Z����Z����Z���b�{�a����cDZZZZZZZZggZZZZZZZZZZZ��Z�����Z��������hZZ�������Z�{�a����Z����Z�Z�������Z����DZZZZZZZZggZZZZZZZZZZZ�����DZZZZZZZZggDZZZZZZZZ��������Z��ZtZ�{�ZtwZ|{����d|{����d|{����uggZ���������Z��������DDZZZZZZZZZZZZ��������Z�}����}{�tZ|���{�ZtwZ�ZvZjhjuggZ}����Z����Z��Z��������DZZZZZZZZZZZZ��������Z���}{�ZtZ�{�ZtwZ{|�b�cuZZZZZZZggZ���Z��������Z�����DZZZZZZZZZZZZ��������Z��~�{�tZ�{�ZuDZZZZZZZZZZZZ��������Z}����tZ�����ZuDZZZZZZZZZZZZ��������Z���{�tZ�{�ZuDZZZZZZZZZZZZ��������Z�{������tZ�{�ZuDZZZZZZZZ��������Z�{}���ZtZ�{�ZtwZkhjuDDZZZZZ�����DZZZZZZZZZZZZggZ}������Z�����Z���Z�������Z�����DZZZZZZZZ��Z�ZwZjhjZ����DZZZZZZZZZZZZZZZZ������ZkhjuDZZZZZZZZ���Z��uDDZZZZZZZZ��ZZ���}{�ZwZkhjZZ����DZZZZZZZZZZZZZZZZ��Z�}����}{�Z����DZZZZZZZZZZZZZZZZZZZZZZZZ������Z�{���k�����uDZZZZZZZZZZZZZZZZ����DZZZZZZZZZZZZZZZZZZZZZZZZ������Z�{���uDZZZZZZZZZZZZZZZZ���Z��uDZZZZZZZZ���Z��uDDZZZZZZZZ��ZZ���}{�ZwZlhjZZ����DZZZZZZZZZZZZZZZZ��Z�}����}{�Z����DZZZZZZZZZZZZZZZZZZZZZZZZ������Zkhji�{�����luDZZZZZZZZZZZZZZZZ����DZZZZZZZZZZZZZZZZZZZZZZZZ������Z�{�����luDZZZZZZZZZZZZZZZZ���Z��uDZZZZZZZZ���Z��uDDZZZZZZZZ��ZZ���}{�ZwZkjhjZZ����DZZZZZZZZZZZZZZZZ��Z�}����}{�Z����DZZZZZZZZZZZZZZZZZZZZZZZZ������Zkhji�{�����kjuDZZZZZZZZZZZZZZZZ����DZZZZZZZZZZZZZZZZZZZZZZZZ������Z�{�����kjuDZZZZZZZZZZZZZZZZ���Z��uDZZZZZZZZ���Z��uDDZZZZZZZZ��Z���}{�ZxZ���b�{�a����cZ����DZZZZZZZZZZZZZZZZ��Z�}����}{�Z����DZZZZZZZZZZZZZZZZZZZZZZZZ������ZjhjuDZZZZZZZZZZZZZZZZ����DZZZZZZZZZZZZZZZZZZZZZZZZ������Z�{��DZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ������Z\�ZxZ���b�{�a����cZ��Z��b�c\DZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ��������Z���uDZZZZZZZZZZZZZZZZZZZZZZZZ������Z�{�a����uDZZZZZZZZZZZZZZZZ���Z��uDZZZZZZZZ���Z��uDDZZZZZZZZggZ������Z��������Z��Z{|�b�cZvZkhjDZZZZZZZZ�����Z���}{�ZxZkjhjZ����DZZZZZZZZZZZZZZZZ���}{�ZtwZ���}{�ZgZkjhjuDZZZZZZZZZZZZZZZZ�{}���ZtwZ�{}���d�{�����kjuDZZZZZZZZ���Z����uDDZZZZZZZZ�����Z���}{�ZxZkhjZ����DZZZZZZZZZZZZZZZZ���}{�ZtwZ���}{�ZgZkhjuDZZZZZZZZZZZZZZZZ�{}���ZtwZ�{}���d�{���uDZZZZZZZZ���Z����uDDZZZZZZZZggZ}������Z�����Z���Z����ZjZvZ���}{�ZvZkDZZZZZZZZ��~�{�ZtwZkhjuDZZZZZZZZ�{������ZtwZ���}{�uDZZZZZZZZ���{�twZ��~�{�ZeZ�{������uDZZZZZZZZ}����ZtwZluDDZZZZZZZZggZ}����Z���Z��������Z���Z��������Z������Z���Z���Z�����DZZZZZZZZ�����ZbZbZb{|�bb���{�ZgZ��~�{�ci���{�cZxZ��cZ��DZZZZZZZZZZZZZZZZZZb{|�b���{�ZgZ��~�{�cZxZ��cZcZ{�~DZZZZZZZZZZZZZZZZZZb}����ZvZ�{��}����ZcZcZ����DZZZZZZZZZZZZZZZZ��~�{�ZtwZ���{�uDZZZZZZZZZZZZZZZZ�{������ZtwZ�{������db���}{�ZiZb�{�b}����cccuDZZZZZZZZZZZZZZZZ���{�ZtwZ��~�{�ZeZ�{������uDZZZZZZZZZZZZZZZZ}����ZtwZ}����ZeZkuDZZZZZZZZ���Z����uDDZZZZZZZZggZ}������Z�����Z�����Z�����Z���b�e�cZwZ���b�cd���b�cDZZZZZZZZ���{�ZtwZ���{�d�{}���uDDZZZZZZZZ��Z�}����}{�Z����DZZZZZZZZZZZZZZZZ���{�ZtwZkhji���{�uDZZZZZZZZ���Z��uDDZZZZZZZZ������Z���{�uDZZZZZ���Z��uDDDZZZZggDZZZZggZ{��������Z���������Z��Z}������Z���DZZZZggDZZZZ��������Z����|b�tZ��Z�{�cZ������Z�����Z��DZZZZZZZZggZ~����������tDZZZZZZZZggZZZZZZZZ�������Z�Z����Z����ZgkZvwZ{|�b�cil��ZvZlDZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZ����DDZZZZZZZZ��������Z�tZ�����ZtwZjuDZZZZZZZZ��������Z�tZ�{�ZtwZ{|�b�cuDDZZZZ�����DZZZZZZZZ��b�ZwZkhjZ��Z�ZwZjhjcZ����DZZZZZZZZZZZZZZZZ������ZjuDZZZZZZZZ���Z��uDDZZZZZZZZ��bZ�ZxZkhjcZ����DZZZZZZZZZZZZZZZZ�����Z�ZxwZlhjZ����DZZZZZZZZZZZZZZZZZZZZZZZZ�ZtwZ�ilhjuDZZZZZZZZZZZZZZZZZZZZZZZZ�ZtwZ�ekuDZZZZZZZZZZZZZZZZ���Z����uDZZZZZZZZZZZZZZZZ������Z�uDZZZZZZZZ���Z��uDDZZZZZZZZggZ�ZvZ�ZvZkDZZZZZZZZ�����Z�ZvZkhjZ����DZZZZZZZZZZZZZZZZ�ZtwZ�dlhjuDZZZZZZZZZZZZZZZZ�ZtwZ�ZgkuDZZZZZZZZ���Z����uDZZZZZZZZ������Z�uDZZZZ���Z����|uDDZZZZ��������Z�~��b�tZ��Z�{�uZ�tZ��Z�����cZ�����Z�{�Z��DZZZZZZZZggZ~����������tDZZZZZZZZggZZZZZZZZ�������Z�dl��DZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZZ����DZZZZ�����DZZZZZZZZ������Z�dblhjZddZ�cuDZZZZ���Z�~��uDDZZZZ��������Z���Zb�ZtZ��Z�{�ZcZ������Z�{�Z��DZZZZZZZZggZ~����������tDZZZZZZZZggZZZZZZZZ���Z��������Z�����������Z��Z�Z���ZkjqphlgksspDZZZZZZZZggDZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZ�cZ�������Z�{�a���Z��Z�����DZZZZZZZZggDZZZZZZZZggZ}��������Zb�cZksslZ�������Z��Z���Z����������Z��Z}���������hDZZZZZZZZggZ{��Z������Z��������hDZZZZZZZZggDZZZZZZZZggZ��������������Z���Z���Z��Z������Z���Z������Z�����fZ����Z��Z�������DZZZZZZZZggZ������������fZ���Z���������Z��������Z����Z���Z���������Z����������DZZZZZZZZggZ���Z���tDZZZZZZZZggZkhZ���������������Z��Z������Z����Z����Z������Z���Z�����Z���������DZZZZZZZZggZ������fZ����Z����Z��Z����������Z���Z���Z���������Z����������hDZZZZZZZZggZlhZ���������������Z��Z������Z����Z����Z���������Z���Z�����Z���������DZZZZZZZZggZ������fZ����Z����Z��Z����������Z���Z���Z���������Z����������Z��Z���DZZZZZZZZggZ�������������Z���i��Z�����Z���������Z��������Z����Z���Z������������hDZZZZZZZZggZmhZ{��Z�����������Z���������Z����������Z��������Z��Z���Z��Z����DZZZZZZZZggZ��������Z����Z�������Z���Z���������Z���������������tDZZZZZZZZggZ����Z�������Z��������Z��������Z���������Z��Z���Z����������Z��DZZZZZZZZggZ}���������fZ|�������Z���Z���Z������������hDZZZZZZZZggZnhZ�������Z���Z����Z��Z���Z����������Z���Z���Z�����Z��Z���DZZZZZZZZggZ������������Z���Z��Z����Z��Z�������Z��Z�������Z��������Z�������DZZZZZZZZggZ����Z����Z��������Z�������Z��������Z�����Z�������Z����������hDZZZZZZZZggDZZZZZZZZggZ����Z�����{�Z��Z�����~~Z|�Z��Z�����Z{�~Z}�����|�����Z��{�Z��aaDZZZZZZZZggZ{�~Z{��Z�����Z��Z�����~Z�{��{����fZ��}��~���fZ|��Z���Z�����~Z��fDZZZZZZZZggZ��Z�����~Z�{��{����Z��Z��}�{��{|�����Z{�~Z������Z���Z{DZZZZZZZZggZ�{���}��{�Z������Z{�Z~��}�{��~hZ��Z��Z���Z��{��Z��Z�����Z��DZZZZZZZZggZ}�����|�����Z|Z��{|�Z���Z{��Z~��}�fZ��~��}�fZ��}�~��{�fZ��}�{�fDZZZZZZZZggZ����{��fZ��Z}��������{�Z~{�{��Zb��}��~���fZ|��Z���Z�����~Z��fDZZZZZZZZggZ���}�����Z��Z��|������Z���~�Z��Z����}�uZ����Z��Z��fZ~{�{fZ��DZZZZZZZZggZ�������uZ��Z|������Z�����������cZ�����Z}{��~Z{�~Z��Z{��Z�����DZZZZZZZZggZ��Z��{|�����fZ�����Z��Z}����{}�fZ����}�Z��{|�����fZ��Z����DZZZZZZZZggZb��}��~���Z������}Z��Z�������cZ{������Z��Z{��Z�{�Z���Z��Z��DZZZZZZZZggZ��Z��Z����Z�����{�fZ��Z��Z{~���~Z��Z��Z�����|�����Z��Z��}�DZZZZZZZZggZ~{�{�hDZZZZZZZZggDZZZZZZZZggZ���tZ����Z��~�Z�������Z���Z���������Z�����Z���Z}Z�������Z��Z���DZZZZZZZZggZZZZZZZZZ��������Z��������Z��Z���Z�Z��~�Z������������Z�������DZZZZZZZZggZZZZZZZZZ�������Z�����Zb}�i��cDDZZZZZZZZ��������Z�tZ�����ZtwZklruDDZZZZZZZZggZ�����Z��Z���b��cZwZ������������ZeZ������������fZ���Z��ZwZke�iklrhDZZZZZZZZggZ����Z���Z����������Z��Z������Z���������Z����������hDZZZZZZZZggZ���Z��������ZmokrnmqljrrrmlZ��Zl�nofZ��Z���Z������Z��Z�����hDZZZZZZZZggZ��Z�������Z�������Z�������Z��Z���������fZ����Z���Z����������DZZZZZZZZggZ�������g��g������Z����������Z��������hZb��������Z����Z���DZZZZZZZZggZ�����Z������Z���Z������Z����Z����Zl�omhcDZZZZZZZZggZ������Z���Z���b�cZ����Z���������Z�����Z�����ZvZkj�goqZ��������DZZZZZZZZggZ����Z���Z��Zg�Z�������hDDZZZZZZZZ����Z�{���}���Z��Z�����Zb�{���{�Z�����ZvxcZ��Z�{�uDDZZZZZZZZ��������Z{kt�{�ZtwZjhjrmmmmmmmmmmmmkqrrlquDZZZZZZZZ��������Z{lt�{�ZtwZjhjklojjjjjjjmqqkqnslmuDZZZZZZZZ��������Z{mt�{�ZtwZjhjjllmlkmssrqsksnnqrjsuDZZZZZZZZ��������Z{nt�{�ZtwZjhjjjnmnrrqqqqqjqpknoqnluDDZZZZZZZZ��������Z������{~tZ�{���}���bjZ��Z�cZtwZbDZZZZZZZZZZZZZZZZjhjfDZZZZZZZZZZZZZZZZjhjjqqrlknjnnljpjmrklnpfDZZZZZZZZZZZZZZZZjhjkoojnkrpomospmolppsnfDZZZZZZZZZZZZZZZZjhjlmkpqjoslrkonqpjrnjpfDZZZZZZZZZZZZZZZZjhjmjqqkporpppqpolmmpnqfDZZZZZZZZZZZZZZZZjhjmrmkrrpnmjlknklpnnrrfDZZZZZZZZZZZZZZZZjhjnorjsompjmklnlqknpqjfDZZZZZZZZZZZZZZZZjhjomlnnoknokrrmqpjnooofDZZZZZZZZZZZZZZZZjhjpjplnplkrkpnrpsqrqrpfDZZZZZZZZZZZZZZZZjhjpqsojppksjrolosnnnonfDZZZZZZZZZZZZZZZZjhjqollmnlklmqolnlmojmsfDZZZZZZZZZZZZZZZZjhjrlnnmppslkjsrrnnpkmrfDZZZZZZZZZZZZZZZZjhjrspklkorprsqpjpsjmllfDZZZZZZZZZZZZZZZZjhjspqlsplpnornonqmkpkrfDZZZZZZZZZZZZZZZZjhkjmqspqsmprkopqoqrnpjfDZZZZZZZZZZZZZZZZjhkkjrknmppmnjlpnmknljmfDZZZZZZZZZZZZZZZZjhkkqqrmjmopopnmjjjkrmpfDZZZZZZZZZZZZZZZZjhklnqjmnqrojkjmlrjojqjfDZZZZZZZZZZZZZZZZjhkmkoqpmoqqrrpkqmkolmpfDZZZZZZZZZZZZZZZZjhkmrnjlmllroslslmlpjlsfDZZZZZZZZZZZZZZZZjhknokrljjsrnnoqojqqlsofDZZZZZZZZZZZZZZZZjhkokskpjnljloqmlkpqomjfDZZZZZZZZZZZZZZZZjhkorpjojmjkqpposjopnokfDZZZZZZZZZZZZZZZZjhkpolnsoqlrsomsjrrmqrpfDZZZZZZZZZZZZZZZZjhkqkrojlopslpokrmnkjpjfDZZZZZZZZZZZZZZZZjhkqrnjqpoqnqlprspjpsnqfDZZZZZZZZZZZZZZZZjhkrnsllmmrnsmrmnkjnkopfDZZZZZZZZZZZZZZZZjhkskmsnrolsssopojnpjnqfDZZZZZZZZZZZZZZZZjhksqrloqnmmlsqoroolkmofDZZZZZZZZZZZZZZZZjhljnlkoonknlrqppmjjpprfDZZZZZZZZZZZZZZZZjhlkjopnqpskjqmojjjlqnkfDZZZZZZZZZZZZZZZZjhlkprqmsmrmjjolmkojlnpfDZZZZZZZZZZZZZZZZjhllmknmookmknjlnjrjjopfDZZZZZZZZZZZZZZZZjhllsmqnkjkjpnrqqmllpnlfDZZZZZZZZZZZZZZZZjhlmooppjqkmklrpjjjmpqlfDZZZZZZZZZZZZZZZZjhlnkqkssmprrpsppjlnqorfDZZZZZZZZZZZZZZZZjhlnqrmpkpmsjnosnlrpoqqfDZZZZZZZZZZZZZZZZjhlomskoljssrjqmlnqjlrofDZZZZZZZZZZZZZZZZjhlossoqolnnmpprpjqkopqfDZZZZZZZZZZZZZZZZjhlpospmonrnspsrnjjmoqqfDZZZZZZZZZZZZZZZZjhlqksmmqkonrnjkjnpmkknfDZZZZZZZZZZZZZZZZjhlqqrprnokjjmjrqkjlnmofDZZZZZZZZZZZZZZZZjhlrmqprkqmkmjqmrnmloksfDZZZZZZZZZZZZZZZZjhlrspmmlslorlsnrmnlrspfDZZZZZZZZZZZZZZZZjhlsonpnlklrsmnlkjpmkssfDZZZZZZZZZZZZZZZZjhmjklpkmmjoqrkssqjnkqqfDZZZZZZZZZZZZZZZZjhmjqjlojmolsnrlqrmjoklfDZZZZZZZZZZZZZZZZjhmklqooqkjjjnlmsokqqlsfDZZZZZZZZZZZZZZZZjhmkrnomqmkkkrjsqnsmrsjfDZZZZZZZZZZZZZZZZjhmlnkksnprponmkpqmmoskfDZZZZZZZZZZZZZZZZjhmlsqomlrpmqloqskprolrfDZZZZZZZZZZZZZZZZjhmmomooonksljqplmmnnrnfDZZZZZZZZZZZZZZZZjhmnjslporpsqjnonjrkrslfDZZZZZZZZZZZZZZZZjhmnpnppqpqmnpkjjrlmnrrfDZZZZZZZZZZZZZZZZjhmoksqpnlmkoprrnlppjpmfDZZZZZZZZZZZZZZZZjhmoqnoorrrslllmkpqsmkpfDZZZZZZZZZZZZZZZZjhmplsjonsmprsknjqklmqpfDZZZZZZZZZZZZZZZZjhmprmloopkkorosskoqmolfDZZZZZZZZZZZZZZZZjhmqmqkpnjsqsmrknrkrrnjfDZZZZZZZZZZZZZZZZjhmqsjqrmolsmnrkkrnpmomfDZZZZZZZZZZZZZZZZjhmrnnkkpsrskjlsrorlpmlfDZZZZZZZZZZZZZZZZjhmrsqkpqokknjnnjnpnsokfDZZZZZZZZZZZZZZZZjhmsnssmrjrlnjonlnlkkkqfDZZZZZZZZZZZZZZZZjhnjjlnmkpnklqnosqnsoqsfDZZZZZZZZZZZZZZZZjhnjonpokjrkjqrkskjonsrfDZZZZZZZZZZZZZZZZjhnkjposslnsrommrrqooorfDZZZZZZZZZZZZZZZZjhnkorlqrsoknmosmksorlofDZZZZZZZZZZZZZZZZjhnljspslsnpnnlmqmqsonmfDZZZZZZZZZZZZZZZZjhnlpjrnmsomkjprknlspskfDZZZZZZZZZZZZZZZZjhnmkkqmnpnrkrkmjjknnpnfDZZZZZZZZZZZZZZZZjhnmplmpqppqqnolqnsoqlpfDZZZZZZZZZZZZZZZZjhnnklqnopjrjoknjsmplrkfDZZZZZZZZZZZZZZZZjhnnplrqkjlplrjnrkpjkkmfDZZZZZZZZZZZZZZZZjhnoklqnpnnkmspmjlonmorfDZZZZZZZZZZZZZZZZjhnoplmqnmmnrkrqnkqqlmlfDZZZZZZZZZZZZZZZZjhnpkkqoqkokllnjrlskqsjfDZZZZZZZZZZZZZZZZjhnppjrsqlsslnommnoqspjfDZZZZZZZZZZZZZZZZjhnqjsqsqkolksjqmkkmsrofDZZZZZZZZZZZZZZZZjhnqornosjnrpsroprsnsnqfDZZZZZZZZZZZZZZZZjhnrjprrolsmnooqjqknlklfDZZZZZZZZZZZZZZZZjhnroojqrkoqrkpjlnjmknsfDZZZZZZZZZZZZZZZZjhnsjmjmsrrjnoolomlspomfDZZZZZZZZZZZZZZZZjhnsojqqlppqsrjmnonmkqkfDZZZZZZZZZZZZZZZZjhnssrlqrpsooppkknjmrllfDZZZZZZZZZZZZZZZZjhojnoopjkjqokskllomsjrfDZZZZZZZZZZZZZZZZjhojslpksjkqsjolmoolmmofDZZZZZZZZZZZZZZZZjhokmsnoqokkjkmnpkjnnjofDZZZZZZZZZZZZZZZZjhokrpjqqpnljrmonpmqsorfDZZZZZZZZZZZZZZZZjholmlnrknmqpokorpjljmpfDZZZZZZZZZZZZZZZZjholqrpqjrspljnroqronkqfDZZZZZZZZZZZZZZZZjhomlnpnqsrrpskknjkssjrfDZZZZZZZZZZZZZZZZjhomqjnknporsqmnoskonmpfDZZZZZZZZZZZZZZZZjhonkosqlrlnmlklkoqmsnqfDZZZZZZZZZZZZZZZZjhonpkmlnmqosqnjqlpjsjsfDZZZZZZZZZZZZZZZZjhoojpnqkkqsolmsnkrlqsmfDZZZZZZZZZZZZZZZZjhoooknkojqonjpkkljjspofDZZZZZZZZZZZZZZZZjhoospkoqrqsmomssoppqqqfDZZZZZZZZZZZZZZZZjhopnjqjkmrlromrqpoppokfDZZZZZZZZZZZZZZZZjhoprojnqmomolprsqnsopkfDZZZZZZZZZZZZZZZZjhoqlsksqomopljkrqnjsllfDZZZZZZZZZZZZZZZZjhoqqmkompojmolnpsnklpjfDZZZZZZZZZZZZZZZZjhorkpskqmspmojpkrlksjjfDZZZZZZZZZZZZZZZZjhorpjnsjnojjmkpnqslnmmfDZZZZZZZZZZZZZZZZjhosjmrqnnppjlkjqsoqjjofDZZZZZZZZZZZZZZZZjhosnqjqkjqqnplkpsmnkqnfDZZZZZZZZZZZZZZZZjhossjjrkrspnolnppjlosnfDZZZZZZZZZZZZZZZZjhpjmlsjroknmrsnkrssprqfDZZZZZZZZZZZZZZZZjhpjqooolojllnmllpplprrfDZZZZZZZZZZZZZZZZjhpkkrjkonkkjppkommksoofDZZZZZZZZZZZZZZZZjhpkpjlsrqqlkoplmrooosjfDZZZZZZZZZZZZZZZZjhpljlnjnjsqokljnnlnomqfDZZZZZZZZZZZZZZZZjhplnnmmlrrjklmpsmjmjmlfDZZZZZZZZZZZZZZZZjhplrpjrposnllqolprjlopfDZZZZZZZZZZZZZZZZjhpmlqppppsoqjplrnmqlkmfDZZZZZZZZZZZZZZZZjhpmpsjqnpllmpksnsrqqrkfDZZZZZZZZZZZZZZZZjhpnkjmkkqsnljpqskjskqkfDZZZZZZZZZZZZZZZZjhpnokmqspkmqmpljqrlsqrfDZZZZZZZZZZZZZZZZjhpnsllqsnpplopkojjnnojfDZZZZZZZZZZZZZZZZjhpommjklqljkksorpnnqlofDZZZZZZZZZZZZZZZZjhpoqmorjqlqjsjmjlmrskkfDZZZZZZZZZZZZZZZZjhppkmsrnrllnoljmsllojlfDZZZZZZZZZZZZZZZZjhpponllpmlonnojokqqjpofDZZZZZZZZZZZZZZZZjhppsnmjpomsnlsrkqmnrqkfDZZZZZZZZZZZZZZZZjhpqmnllpqolklmojnnkknlfDZZZZZZZZZZZZZZZZjhpqqmsrrlmosjsljjqmskkfDZZZZZZZZZZZZZZZZjhprkmosllnrjqlmrljplpqfDZZZZZZZZZZZZZZZZjhpromjnjjmjsrlrkkjjmslfDZZZZZZZZZZZZZZZZjhprslmmlrklmrooqomrjkqfDZZZZZZZZZZZZZZZZjhpsmknqkrjopjkkqqjmrplcuDDZZZZZZZZ��������Z������{��tZ�{���}���bjZ��Z�cZtwZbDZZZZZZZZZZZZZZZZjhjfDZZZZZZZZZZZZZZZZgjhjjjjjjjjjjjjjjonmllssmrnljjnsfDZZZZZZZZZZZZZZZZjhjjjjjjjjjjjjjjkqlqnopqnssqjpkfDZZZZZZZZZZZZZZZZgjhjjjjjjjjjjjjjkmlmjkqrkrllslmmfDZZZZZZZZZZZZZZZZgjhjjjjjjjjjjjjjkkonolqplrlrsrqlfDZZZZZZZZZZZZZZZZgjhjjjjjjjjjjjjjjnppolsnpssormjjfDZZZZZZZZZZZZZZZZjhjjjjjjjjjjjjjoknrrnsoqlprorkjfDZZZZZZZZZZZZZZZZgjhjjjjjjjjjjjjjlomlkprsnmkkqnnofDZZZZZZZZZZZZZZZZgjhjjjjjjjjjjjjjolkmpljpmskmpojnfDZZZZZZZZZZZZZZZZgjhjjjjjjjjjjjjjkrksojpjjmjkprrkfDZZZZZZZZZZZZZZZZjhjjjjjjjjjjjjjpmlsjposorqlnonnfDZZZZZZZZZZZZZZZZjhjjjjjjjjjjjjjrpknoklsmpjrqrknfDZZZZZZZZZZZZZZZZgjhjjjjjjjjjjjjjqmooqqjlksnmojlrfDZZZZZZZZZZZZZZZZjhjjjjjjjjjjjjjspmrjpqporoollqqfDZZZZZZZZZZZZZZZZjhjjjjjjjjjjjjjqosrpmposqksnknkfDZZZZZZZZZZZZZZZZjhjjjjjjjjjjjjjloqssssklrmjpssjfDZZZZZZZZZZZZZZZZgjhjjjjjjjjjjjjjnponqlsqnqosrnnnfDZZZZZZZZZZZZZZZZgjhjjjjjjjjjjjjjqoopsljprqnokmmpfDZZZZZZZZZZZZZZZZjhjjjjjjjjjjjjkjksoqmollmqjrnqlfDZZZZZZZZZZZZZZZZgjhjjjjjjjjjjjjkqmksjmnnjpnllmjpfDZZZZZZZZZZZZZZZZgjhjjjjjjjjjjjjjqqkrjjkmmprlrjsrfDZZZZZZZZZZZZZZZZjhjjjjjjjjjjjjkjsrjqonjssroolmrfDZZZZZZZZZZZZZZZZgjhjjjjjjjjjjjjjljnqlmoqrjjnpksofDZZZZZZZZZZZZZZZZgjhjjjjjjjjjjjjjrmqljskjsslmosklfDZZZZZZZZZZZZZZZZjhjjjjjjjjjjjjknjrrklqsmqkkkkmofDZZZZZZZZZZZZZZZZjhjjjjjjjjjjjjklrpsjkqkoqorrloqfDZZZZZZZZZZZZZZZZjhjjjjjjjjjjjjkqqrrrojqqrksrkjpfDZZZZZZZZZZZZZZZZjhjjjjjjjjjjjjjpnnjropkojpsprskfDZZZZZZZZZZZZZZZZjhjjjjjjjjjjjjkpkmlrllppqlnjrllfDZZZZZZZZZZZZZZZZgjhjjjjjjjjjjjjjqonjskpokksopkrrfDZZZZZZZZZZZZZZZZgjhjjjjjjjjjjjjjjjmpojqkrrrmkqsjfDZZZZZZZZZZZZZZZZjhjjjjjjjjjjjjjskljsmqlnssknsrnfDZZZZZZZZZZZZZZZZjhjjjjjjjjjjjjkropqoqjsosqspjkjfDZZZZZZZZZZZZZZZZgjhjjjjjjjjjjjjjmknslpojpoksknrmfDZZZZZZZZZZZZZZZZgjhjjjjjjjjjjjjjsmjsnosnsoksprrsfDZZZZZZZZZZZZZZZZjhjjjjjjjjjjjjkqsknmmrpjkmlskkqfDZZZZZZZZZZZZZZZZgjhjjjjjjjjjjjjjkmjlsqsqkqmmjrppfDZZZZZZZZZZZZZZZZjhjjjjjjjjjjjjlmjsqmrolkqorpsmsfDZZZZZZZZZZZZZZZZjhjjjjjjjjjjjjlmsssonjnrnlkkqmqfDZZZZZZZZZZZZZZZZjhjjjjjjjjjjjjkomsmqqpkqnnoonjrfDZZZZZZZZZZZZZZZZgjhjjjjjjjjjjjjmprqjnlrmkormqpqrfDZZZZZZZZZZZZZZZZjhjjjjjjjjjjjjmpsljmqojrljrjjrsfDZZZZZZZZZZZZZZZZgjhjjjjjjjjjjjjjsmrmnkqllmppmpssfDZZZZZZZZZZZZZZZZjhjjjjjjjjjjjjjsnmmmsrkrsoklpsjfDZZZZZZZZZZZZZZZZjhjjjjjjjjjjjjnknrkmkrqjnloroprfDZZZZZZZZZZZZZZZZgjhjjjjjjjjjjjjjmqslmkpnrjljsmknfDZZZZZZZZZZZZZZZZjhjjjjjjjjjjjjjrnjmkopmjnqslnlnfDZZZZZZZZZZZZZZZZgjhjjjjjjjjjjjjmnlplsmnmnrlronlsfDZZZZZZZZZZZZZZZZjhjjjjjjjjjjjjnmqklksksoqnlsknofDZZZZZZZZZZZZZZZZgjhjjjjjjjjjjjjkjnqoqojjorqqponkfDZZZZZZZZZZZZZZZZgjhjjjjjjjjjjjjkkkkrpqkmrsoosmlmfDZZZZZZZZZZZZZZZZjhjjjjjjjjjjjjmqonsoqqloqlosromfDZZZZZZZZZZZZZZZZjhjjjjjjjjjjjjkmsklrnklklksqopofDZZZZZZZZZZZZZZZZjhjjjjjjjjjjjjkjqqoqnmjmqoqlpnjfDZZZZZZZZZZZZZZZZjhjjjjjjjjjjjjlsmskroskrqpnrjjjfDZZZZZZZZZZZZZZZZgjhjjjjjjjjjjjjnlqsjojsjpjjpjqqnfDZZZZZZZZZZZZZZZZjhjjjjjjjjjjjjllqqnjqpkknjmsooofDZZZZZZZZZZZZZZZZjhjjjjjjjjjjjjkjrnsopspllspqsklfDZZZZZZZZZZZZZZZZgjhjjjjjjjjjjjjlmjqmrjksnoqjoqorfDZZZZZZZZZZZZZZZZjhjjjjjjjjjjjjkoqpkljmqqmspsnmofDZZZZZZZZZZZZZZZZjhjjjjjjjjjjjjjmmnoqkjlpsonnjrlfDZZZZZZZZZZZZZZZZgjhjjjjjjjjjjjjnkolokorjpmnmpklmfDZZZZZZZZZZZZZZZZjhjjjjjjjjjjjjmlpoopsrrspsjqknpfDZZZZZZZZZZZZZZZZgjhjjjjjjjjjjjjnnqjnlpojkjnolnnpfDZZZZZZZZZZZZZZZZjhjjjjjjjjjjjjmnolqpnqsoljmsqqlfDZZZZZZZZZZZZZZZZgjhjjjjjjjjjjjjjqjnrsplmslkjsqnpfDZZZZZZZZZZZZZZZZjhjjjjjjjjjjjjkkqqpsqrqokmpslknfDZZZZZZZZZZZZZZZZgjhjjjjjjjjjjjjkjqqnmnknpkpjsoqrfDZZZZZZZZZZZZZZZZjhjjjjjjjjjjjjlkrpmmnmlsmlkoskjfDZZZZZZZZZZZZZZZZjhjjjjjjjjjjjjlnkmlpmsnskmmmkmkfDZZZZZZZZZZZZZZZZjhjjjjjjjjjjjjmsjoqnplljsrmjqjjfDZZZZZZZZZZZZZZZZgjhjjjjjjjjjjjjlpoqjpqsljmopjqokfDZZZZZZZZZZZZZZZZjhjjjjjjjjjjjjmqkmoknksksosljlkfDZZZZZZZZZZZZZZZZgjhjjjjjjjjjjjjkqkppslkmmpjrlnmkfDZZZZZZZZZZZZZZZZgjhjjjjjjjjjjjjlrporlrokoqsknmomfDZZZZZZZZZZZZZZZZgjhjjjjjjjjjjjjlmrklonllpmnnprjsfDZZZZZZZZZZZZZZZZjhjjjjjjjjjjjjjpoqpposqprorjjplfDZZZZZZZZZZZZZZZZgjhjjjjjjjjjjjjlrlkjknmrnpkrklpqfDZZZZZZZZZZZZZZZZjhjjjjjjjjjjjjkjqjksmkqplkknlonfDZZZZZZZZZZZZZZZZjhjjjjjjjjjjjjkrkksmnpmppnnkkkjfDZZZZZZZZZZZZZZZZjhjjjjjjjjjjjjjsrnjnpolqrlmlplqfDZZZZZZZZZZZZZZZZgjhjjjjjjjjjjjjmmknskojlrlqolonlfDZZZZZZZZZZZZZZZZgjhjjjjjjjjjjjjkrmjlroqmopjnkpprfDZZZZZZZZZZZZZZZZgjhjjjjjjjjjjjjkpljqnjjkopqnnsnsfDZZZZZZZZZZZZZZZZjhjjjjjjjjjjjjnrmjmmknsnsoomljkfDZZZZZZZZZZZZZZZZgjhjjjjjjjjjjjjqkopjoomkqlmrlkkofDZZZZZZZZZZZZZZZZjhjjjjjjjjjjjjrrrlklmsokroqkroofDZZZZZZZZZZZZZZZZgjhjjjjjjjjjjjjmjsjjorjokmlmrlnnfDZZZZZZZZZZZZZZZZgjhjjjjjjjjjjjjpkjqpooksqlroknspfDZZZZZZZZZZZZZZZZjhjjjjjjjjjjjjmoposspsppmmnqrmjfDZZZZZZZZZZZZZZZZjhjjjjjjjjjjjjmoqrlmsposklqpmrmfDZZZZZZZZZZZZZZZZgjhjjjjjjjjjjjjnpllpjrqjjkonnoqrfDZZZZZZZZZZZZZZZZjhjjjjjjjjjjjjpllqsqplskqllokopfDZZZZZZZZZZZZZZZZjhjjjjjjjjjjjjqlrmrsnqlqljpoqnkfDZZZZZZZZZZZZZZZZjhjjjjjjjjjjjjlprjspnppkolkkpqmfDZZZZZZZZZZZZZZZZgjhjjjjjjjjjjjjkjspjrlojnpjoslqrfDZZZZZZZZZZZZZZZZjhjjjjjjjjjjjjjlmkksnsmrmrjjomqfDZZZZZZZZZZZZZZZZgjhjjjjjjjjjjjjornpsjorjjolsslnqfDZZZZZZZZZZZZZZZZgjhjjjjjjjjjjjjjlkjmqnrlokknnnsnfDZZZZZZZZZZZZZZZZgjhjjjjjjjjjjjjlmmlmkrlsnoorqnjrfDZZZZZZZZZZZZZZZZgjhjjjjjjjjjjjjnlmmmpsnlrrknkskpfDZZZZZZZZZZZZZZZZgjhjjjjjjjjjjjjnmsmmsmqspsqmqrnnfDZZZZZZZZZZZZZZZZjhjjjjjjjjjjjjnkmnkpnqjqmrmoopofDZZZZZZZZZZZZZZZZjhjjjjjjjjjjjjjprnkqpmpnkosknppfDZZZZZZZZZZZZZZZZjhjjjjjjjjjjjjnqoroomnjjnnmjpnkfDZZZZZZZZZZZZZZZZjhjjjjjjjjjjjjrmpqspqrpqnqoqpsofDZZZZZZZZZZZZZZZZgjhjjjjjjjjjjjjroqpmqmnpnpporpnjfDZZZZZZZZZZZZZZZZjhjjjjjjjjjjjjlkskmlrkllsmnjjslfDZZZZZZZZZZZZZZZZgjhjjjjjjjjjjjjpllnlrnlompnmkknrfDZZZZZZZZZZZZZZZZgjhjjjjjjjjjjjjkjsrmosnmlonmrnmjfDZZZZZZZZZZZZZZZZjhjjjjjjjjjjjjpomkjnmkmqqpmmpokfDZZZZZZZZZZZZZZZZgjhjjjjjjjjjjjjnqorjkssjlkqkjqpsfDZZZZZZZZZZZZZZZZgjhjjjjjjjjjjjjmqronloklponoqjnjfDZZZZZZZZZZZZZZZZjhjjjjjjjjjjjjnjsmslmmlkrpqrppnfDZZZZZZZZZZZZZZZZjhjjjjjjjjjjjjrqnlnmrmsknrorlskfDZZZZZZZZZZZZZZZZjhjjjjjjjjjjjjlolkrkrrnoprnlrrlfDZZZZZZZZZZZZZZZZgjhjjjjjjjjjjjjjmpjrkmkmpjnllooqfDZZZZZZZZZZZZZZZZgjhjjjjjjjjjjjjojokroooslnlrjsjlfDZZZZZZZZZZZZZZZZjhjjjjjjjjjjjjqrpssnjmmlmmoomkqfDZZZZZZZZZZZZZZZZgjhjjjjjjjjjjjjpqjljrqpspksnsjpjfDZZZZZZZZZZZZZZZZjhjjjjjjjjjjjjkpkjroqoqomsmlnorfDZZZZZZZZZZZZZZZZjhjjjjjjjjjjjjorolqkrrnmplokojsfDZZZZZZZZZZZZZZZZgjhjjjjjjjjjjjjmolnpqoqlsqsjnqskfDZZZZZZZZZZZZZZZZgjhjjjjjjjjjjjjkrmqljrnnsoplsjorfDZZZZZZZZZZZZZZZZjhjjjjjjjjjjjjrrpjpprsrkmnsnskpfDZZZZZZZZZZZZZZZZjhjjjjjjjjjjjjppnrplprjqknprqjjfDZZZZZZZZZZZZZZZZjhjjjjjjjjjjjjpmrmkpkokqjpnpoksfDZZZZZZZZZZZZZZZZjhjjjjjjjjjjjjloknnlmjqlrmqpjqlfDZZZZZZZZZZZZZZZZgjhjjjjjjjjjjjjkqlmsnnnolopknrmncuDDZZZZZZZZ��������Z�fZ�t�����uDZZZZZZZZ��������Z�kfZ�lfZ�fZ�fZ�fZ�lfZ�tZ�{�uDZZZZZZZZ��������Z���tZ�{�ZtwZjhjugg����Z��������Z��Z��Z��������Z�������Z������DZZZZZZZZ��������Z��tZ�{�ZtwZkhjuZgg����Z��������Z��Z��Z��������Z�������Z������DDZZZZZZZZggZ������Z����bcfZ�����bcuDDZZZZZZZZ��������Z�kt�{�uDDZZZZZ�����DDZZZZZZZZggZ}����Z��������Z��Z��������DZZZZZZZZ��ZbZ�ZvwZjhjZcZ����DZZZZZZZZZZZZZZZZ������Z�{��DZZZZZZZZZZZZZZZZZZZZZZZZ������Z\�ZvwZjhjZ��Z���b�c\DZZZZZZZZZZZZZZZZZZZZZZZZ��������Z����uDZZZZZZZZZZZZZZZZ������b�{�a���cuDZZZZZZZZ���Z��uDDZZZZZZZZggZ}������Z�����Z���Z�������Z�����DZZZZZZZZ��ZbZ�ZwZkhjZcZ����DZZZZZZZZZZZZZZZZ������ZjhjuDZZZZZZZZ���Z��uDDZZZZZZZZ��ZbZ�ZwZ�{���ZcZ����DZZZZZZZZZZZZZZZZ������ZkhjuDZZZZZZZZ���Z��uDDZZZZZZZZggZ{�������Z���������tZkZvwZ�ZvZluZ�il��ZwZ�uDZZZZZZZZggZ�ZwZ�dbkZeZ�i�cZ���Z���ZvwZl�grDDZZZZZZZZ�ZtwZ����|b�cuDZZZZZZZZ�ZtwZ�~��b�fZg�cuDZZZZZZZZ�ZtwZ�����b�{�b�cdb�gkhjccuZggZ}Z����Z����ZjhoZ���Z��������DZZZZZZZZ�kZtwZbkhji�{�b�ccZdZ�{�b�cZeZkhjuZgg�kdklrZ��Z��Z�����Z��Z�klrfokl�DZZZZZZZZ�lZtwZ�ZgZ�kuDDZZZZZZZZggZ{����������Z���������Z���Z���bke�li�kcZ�wZ�ZeZ�DZZZZZZZZ�ZtwZkhjiblhjd�ke�lcuDZZZZZZZZ�ZtwZlhjd�ld�uDZZZZZZZZ�ZtwZ�d�uDZZZZZZZZ�ZtwZ�d�db{kZeZ�db{lZeZ�db{mZeZ�d{ncccuDDZZZZZZZZggZ}���ZktZ�kZwZ�Z�������Z��Zl�gnmZ��������hZ�����Z�ZvZl�grfDZZZZZZZZggZZZZZZZ�kZ���Z��Z����ZmoZ����fZ���Z�kd�kZ��Z�����fZ��Z�kZ���ZvZrZ����hDZZZZZZZZggZZZZZZZ��Z����Z����Z�������Z��Z��d���l���ZeZ�������������Z�ZvZqojhDZZZZZZZZggDZZZZZZZZ��ZbZ�ZiwZjZ��Z�ZiwZjcZ����DZZZZZZZZZZZZZZZZ�kZtwZ�ZeZokmhjuDZZZZZZZZZZZZZZZZ�kZtwZ�kZgZokmhjuDDZZZZZZZZZZZZZZZZggZ}���ZltZ�kg��ZvZkilophZ���Z�gZ���Z�gZ���������Z�����Z���Z����DZZZZZZZZZZZZZZZZggZZZZZZZZ�kZwZ�Z��ZlnZ����hDZZZZZZZZZZZZZZZZggDZZZZZZZZ����DZZZZZZZZZZZZZZZZ�kZtwZ�uDZZZZZZZZZZZZZZZZgg����}b�kcuZgg��Z�Z����Z��Z�kZwZb������cZb�����cZb�kcDZZZZZZZZ���Z��uDDZZZZZZZZ�lZtwZblhjdb�lZgZ�kd�kcZgZ�kd�lcZdZ�uDZZZZZZZZggZ�kZeZ�lZwZl�ibl�e�cZ��Z�����Z���������hDDZZZZZZZZggZ���b�cZwZ���bl��d�kdbke�li�kccZwDZZZZZZZZggZb�d���l���e������{~b�ce�kcZeZb�d���l���e������{��b�ce�cuDZZZZZZZZggZb�����cZeZb����cDDZZZZZZZZ�kZtwZ�kZeZ�{�b�cd������{~b�cZeZ������{~b�cuZZZZZZZZggZ����DZZZZZZZZ�lZtwZb�lZeZ������{��b�ccZeZ�uZZZZZZZZggZ����DZZZZZZZZ�lZtwZ�lZeZ������{��b�cd�{�b�cuDZZZZZZZZ������Zb�kZeZ�lcuDZZZZ���Z���uDDDZZZZ��������Z���lZb�tZ��Z�{�cZ������Z�{�Z��DZZZZZZZZggZ~����������tDZZZZZZZZggZZZZZZZZ���Z��������Z�����������Z��Z�Z���ZkjqphlgksspDZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZ�cZ�������Z�{�a���Z��Z�����DZZZZ�����DZZZZZZZZggZ}����Z��������Z��Z���������DZZZZZZZZ��ZbZ�ZvwZjhjZcZZ����DZZZZZZZZZZZZZZZZ������Z�{��DZZZZZZZZZZZZZZZZZZZZZZZZ������Z\�ZvwZjhjZ��Z���lb�c\DZZZZZZZZZZZZZZZZZZZZZZZZ��������Z����uDZZZZZZZZZZZZZZZZ������b�{�a���cuDZZZZZZZZ���Z��uDDZZZZZZZZggZ}������Z�����Z���Z�������Z�����DZZZZZZZZ��ZbZ�ZwZkhjZcZ����DZZZZZZZZZZZZZZZZ������ZjhjuDZZZZZZZZ���Z��uDDZZZZZZZZ��ZbZ�ZwZlhjZcZ����DZZZZZZZZZZZZZZZZ������ZkhjuDZZZZZZZZ���Z��uDDZZZZZZZZggZ}������Z�����Z���Z�������Z����DZZZZZZZZ������ZbZ�{������l����d���b�cZcuDZZZZ���Z���luDDDZZZZ��������Z���kjZb�tZ��Z�{�cZ������Z�{�Z��DZZZZZZZZggZ~����������tDZZZZZZZZggZZZZZZZZ���Z��������Z�����������Z��Z�Z���ZkjqphlgksspDZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZ�cZ�������Z�{�a���Z��Z�����DZZZZ�����DZZZZZZZZggZ}����Z��������Z��Z���������DZZZZZZZZ��ZbZ�ZvwZjhjZcZZ����DZZZZZZZZZZZZZZZZZZZ������Z�{��DZZZZZZZZZZZZZZZZZZZZZZZZ������Z\�ZvwZjhjZ��Z���kjb�c\DZZZZZZZZZZZZZZZZZZZZZZZZ��������Z����uDZZZZZZZZZZZZZZZZZZZ������b�{�a���cuDZZZZZZZZ���Z��uDDZZZZZZZZggZ}������Z�����Z���Z�������Z�����DZZZZZZZZ��ZbZ�ZwZkhjZcZ����DZZZZZZZZZZZZZZZZ������ZjhjuDZZZZZZZZ���Z��uDDZZZZZZZZ��ZbZ�ZwZkjhjZcZ����DZZZZZZZZZZZZZZZZ������ZkhjuDZZZZZZZZ���Z��uDDZZZZZZZZggZ}������Z�����Z���Z�������Z����DZZZZZZZZ������ZbZ�{������kj����d���b�cZcuDZZZZ���Z���kjuDDDZZZZ��������Z���Zb�tZ��Z�{�uZ|{�tZ��Z�{�cZ������Z�{�Z��DZZZZZZZZggZ~����������tDZZZZZZZZggZZZZZZZZ���Z��������Z�����������Z��Z�Z���ZkjqphlgksspDZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZ�cZ�������Z�{�a���Z��Z�����DZZZZ�����DZZZZZZZZggZ}����Z��������Z��Z���������DZZZZZZZZ��ZbZ�ZvwZjhjZcZZ����DZZZZZZZZZZZZZZZZZ������Z�{��DZZZZZZZZZZZZZZZZZZZZZZZZ������Z\�ZvwZjhjZ��Z���b�fZ|{�c\DZZZZZZZZZZZZZZZZZZZZZZZZ��������Z����uDZZZZZZZZZZZZZZZZZ������b�{�a���cuDZZZZZZZZ���Z��uDDZZZZZZZZ��ZbZ|{�ZvwZjhjZ��Z|{�ZwZkhjZcZZ����DZZZZZZZZZZZZZZZZZ������Z�{��DZZZZZZZZZZZZZZZZZZZZZZZZ������Z\|{�ZvwZjhjZ��Z|{�ZwZkhjZ��Z���b�fZ|{�c\DZZZZZZZZZZZZZZZZZZZZZZZZ��������Z����uDZZZZZZZZZZZZZZZZZ������b�{�a���cuDZZZZZZZZ���Z��uDDZZZZZZZZggZ}������Z�����Z���Z�������Z�����DZZZZZZZZ��ZbZ�ZwZkhjZcZ����DZZZZZZZZZZZZZZZZ������ZjhjuDZZZZZZZZ���Z��uDDZZZZZZZZ��ZbZ�ZwZ|{�ZcZ����DZZZZZZZZZZZZZZZZ������ZkhjuDZZZZZZZZ���Z��uDDZZZZZZZZggZ}������Z�����Z���Z�������Z����DZZZZZZZZ������ZbZ���b�ci���b|{�ccuDZZZZ���Z���uDDDZZZZ��������ZZ���Zb�ZtZ��Z�{�ZcZ������Z�{�Z��DZZZZZZZZggZ~����������tDZZZZZZZZggZZZZZZZZZ���Z��������Z�����������Z��Z�Z���ZkjqphlgksspDZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZZ�cZ���bg�cZwZg���b�cDZZZZZZZZggZZZZZZZZZ�cZ���b�cZwZ�Z��Z{|�b�cZvZ��DZZZZZZZZggZZZZZZZZZ�cZ���b�cZwZ�ZgZ�ddmim[Z��Z��ZvZ{|�b�cZvZ|{����DZZZZZZZZggZZZZZZZZZ�cZ���b�{����������lZgZ�cZwZ}��b�cDZZZZZZZZggZZZZZZZZZ�cZ}��b�cZwZkhjZgZjhod�ddlZ��Z{|�b�cZvZ��DZZZZZZZZggZZZZZZZZZ�cZ}��b�cZwZkhjZgZjhod�ddlZeZb�ddncin[Z��DZZZZZZZZggZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ��vZ{|�b�cZv|{����DDZZZZZZZZ��������Z��ZtZ�{�ZtwZ|{����d|{����uZggZ}����������Z��������DDZZZZZZZZ��������Z�ZtZ�����uDZZZZZZZZ��������Z��{���ZtZ|���{�ZtwZ�ZvZjhjuDZZZZZZZZ��������Z���}{�ZtZ�{�ZtwZ{|�b�cZuDZZZZZZZZ��������Z�{��tZ�{�uDZZZZZZZZ��������Z���ZtZ�{�uDDZZZZ�����DZZZZZZZZggZ����Z���}{�ZvZ�{���l���DZZZZZZZZ��Z���}{�ZxZ�{���l���Z����DZZZZZZZZZZZZZZZZ���ZtwZ�����b���}{�i�{���l���cuDZZZZZZZZZZZZZZZZ���}{�ZtwZ���}{�ZgZ���d�{���l���uDZZZZZZZZ���Z��uDDZZZZZZZZ��Z���}{�ZvZjhjZ����DZZZZZZZZZZZZZZZZ������Z�{��DZZZZZZZZZZZZZZZZZZZZZZZZ������Z\���}{�ZvwZjhjZ�����Z���������Z��Z���b�c\DZZZZZZZZZZZZZZZZZZZZZZZZ��������Z����uDZZZZZZZZZZZZZZZZ���}{�ZtwZg���}{�uDZZZZZZZZ���Z��uDDZZZZZZZZggZ}������Z�����Z���Z�������Z�����DZZZZZZZZ��Z���}{�ZwZjhjZZ��Z���}{�ZwZ�{���l���Z��Z���}{�ZwZ�{�����ZZ����DZZZZZZZZZZZZZZZZ������ZjhjuDZZZZZZZZ���Z��uDDZZZZZZZZ��ZZ���}{�ZwZ�{����������lZ����DZZZZZZZZZZZZZZZZ��Z��{���Z����DZZZZZZZZZZZZZZZZZZZZZZZZ������ZgkhjuDZZZZZZZZZZZZZZZZ����DZZZZZZZZZZZZZZZZZZZZZZZZ������ZkhjuDZZZZZZZZZZZZZZZZ���Z��uDZZZZZZZZ���Z��uDDZZZZZZZZ��ZZ���}{�ZwZ�{���m��������lZ����DZZZZZZZZZZZZZZZZ��Z��{���Z����DZZZZZZZZZZZZZZZZZZZZZZZZ������ZkhjuDZZZZZZZZZZZZZZZZ����DZZZZZZZZZZZZZZZZZZZZZZZZ������ZgkhjuDZZZZZZZZZZZZZZZZ���Z��uDZZZZZZZZ���Z��uDDZZZZZZZZ��Z���}{�ZvZ��Z����DZZZZZZZZZZZZZZZZ��Z��{���Z����DZZZZZZZZZZZZZZZZZZZZZZZZ������Zg���}{�uDZZZZZZZZZZZZZZZZ����DZZZZZZZZZZZZZZZZZZZZZZZZ������Z���}{�uDZZZZZZZZZZZZZZZZ���Z��uDZZZZZZZZ����DZZZZZZZZZZZZZZZZ��Z���}{�ZvZ|{����Z����DZZZZZZZZZZZZZZZZZZZZZZZZ���ZtwZ���}{�ZgZb���}{�d���}{�d���}{�ciphjuDZZZZZZZZZZZZZZZZZZZZZZZZ��Z��{���Z����DZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ������Zg���uDZZZZZZZZZZZZZZZZZZZZZZZZ����DZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ������Z���uDZZZZZZZZZZZZZZZZZZZZZZZZ���Z��uDZZZZZZZZZZZZZZZZ���Z��uDZZZZZZZZ���Z��uDDZZZZZZZZ���ZtwZ�{�����ZgZ���}{�uDZZZZZZZZ��Z{|�b���cZvZ��Z����DZZZZZZZZZZZZZZZZ��Z��{���Z����DZZZZZZZZZZZZZZZZZZZZZZZZ������Zg���uDZZZZZZZZZZZZZZZZ����DZZZZZZZZZZZZZZZZZZZZZZZZ������Z���uDZZZZZZZZZZZZZZZZ���Z��uDZZZZZZZZ����DZZZZZZZZZZZZZZZZ��Z{|�b���cZvZ|{����Z����DZZZZZZZZZZZZZZZZZZZZZZZZ���ZtwZ���ZgZb���d���d���ciphjuDZZZZZZZZZZZZZZZZZZZZZZZZ��Z��{���Z����DZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ������Zg���uDZZZZZZZZZZZZZZZZZZZZZZZZ����DZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ������Z���uDZZZZZZZZZZZZZZZZZZZZZZZZ���Z��uDZZZZZZZZZZZZZZZZ���Z��uDZZZZZZZZ���Z��uDDZZZZZZZZ���ZtwZ�{���l���ZgZ���}{�uDZZZZZZZZ��Z{|�b���cZvZ��Z����DZZZZZZZZZZZZZZZZ��Z��{���Z����DZZZZZZZZZZZZZZZZZZZZZZZZ������Z���uDZZZZZZZZZZZZZZZZ����DZZZZZZZZZZZZZZZZZZZZZZZZ������Zg���uDZZZZZZZZZZZZZZZZ���Z��uDZZZZZZZZ����DZZZZZZZZZZZZZZZZ��Z{|�b���cZvZ|{����Z����DZZZZZZZZZZZZZZZZZZZZZZZZ���ZtwZ���ZgZb���d���d���ciphjuDZZZZZZZZZZZZZZZZZZZZZZZZ��Z��{���Z����DZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ������Z���uDZZZZZZZZZZZZZZZZZZZZZZZZ����DZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ������Zg���uDZZZZZZZZZZZZZZZZZZZZZZZZ���Z��uDZZZZZZZZZZZZZZZZ���Z��uDZZZZZZZZ���Z��uDDZZZZZZZZ���ZtwZ{|�b�{����������lZgZ���}{�cuDZZZZZZZZ��Z���ZvZ��Z����DZZZZZZZZZZZZZZZZ���ZtwZkhjZgZ���d���djhouDZZZZZZZZZZZZZZZZ��Z��{���Z����DZZZZZZZZZZZZZZZZZZZZZZZZ������Zg���uDZZZZZZZZZZZZZZZZ����DZZZZZZZZZZZZZZZZZZZZZZZZ������Z���uDZZZZZZZZZZZZZZZZ���Z��uDZZZZZZZZ����DZZZZZZZZZZZZZZZZ��Z���ZvZ|{����Z����DZZZZZZZZZZZZZZZZZZZZZZZZ���ZtwZkhjZg���d���djhoZeZ���d���d���d���ilnhjuDZZZZZZZZZZZZZZZZZZZZZZZZ��Z��{���Z����DZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ������Zg���uDZZZZZZZZZZZZZZZZZZZZZZZZ����DZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ������Z���uDZZZZZZZZZZZZZZZZZZZZZZZZ���Z��uDZZZZZZZZZZZZZZZZ���Z��uDZZZZZZZZ���Z��uDDZZZZZZZZ���ZtwZ{|�b�{���m��������lZgZ���}{�cuDZZZZZZZZ��Z���ZvZ��Z����DZZZZZZZZZZZZZZZZ���ZtwZkhjZgZ���d���djhouDZZZZZZZZZZZZZZZZ��Z��{���Z����DZZZZZZZZZZZZZZZZZZZZZZZZ������Z���uDZZZZZZZZZZZZZZZZ����DZZZZZZZZZZZZZZZZZZZZZZZZ������Zg���uDZZZZZZZZZZZZZZZZ���Z��uDZZZZZZZZ����DZZZZZZZZZZZZZZZZ��Z���ZvZ|{����Z����DZZZZZZZZZZZZZZZZZZZZZZZZ���ZtwZkhjZg���d���djhoZeZ���d���d���d���ilnhjuDZZZZZZZZZZZZZZZZZZZZZZZZ��Z��{���Z����DZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ������Z���uDZZZZZZZZZZZZZZZZZZZZZZZZ����DZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ������Zg���uDZZZZZZZZZZZZZZZZZZZZZZZZ���Z��uDZZZZZZZZZZZZZZZZ���Z��uDZZZZZZZZ���Z��uDDZZZZZZZZggZ}������Z�����Z���Z�������Z�����DZZZZZZZZ��Zbb���}{�ZvZ�{����������lZcZ���Zb���}{�ZxZjhjccZ����DZZZZZZZZZZZZZZZZZ�{��twZZ}��~�}bZ�}fZjhjfZ�fZlqfZ���{����cbkcuDZZZZZZZZ���Z��uDDZZZZZZZZ�ZtwZ�����ZbZ�����b���}{�i�{����������lccuDZZZZZZZZ����Z��{~�{��bZ�Z���ZncZ��DZZZZZZZZZZZ����ZjZwxDZZZZZZZZZZZZZZZZ�{��ZtwZ}��~�}bZ�}fZjhjfZ���}{�fZlqfZ���{����cbkcuDZZZZZZZZZZZ����ZkZwxDZZZZZZZZZZZZZZZZ�{��ZtwZ}��~�}bZ�}fZjhjfZ���}{�ZgZ�{����������lfZlqfDZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ���{����cbjcuDZZZZZZZZZZZ����ZlZwxDZZZZZZZZZZZZZZZZ�{��ZtwZg}��~�}bZ�}fZjhjfZ���}{�ZgZ�{�����fZlqfZ���{����cbkcuDZZZZZZZZZZZ����ZmZwxDZZZZZZZZZZZZZZZZ�{��ZtwZg}��~�}bZ�}fZjhjfZ���}{�ZgZ�{���m��������lfZlqfDZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ���{����cbjcuDZZZZZZZZ���Z����uDDZZZZZZZZ��Z��{���Z����DZZZZZZZZZZZZZZZZ������Zg�{��uDZZZZZZZZ����DZZZZZZZZZZZZZZZZ������Z�{��uDZZZZZZZZ���Z��uDZZZZ���Z���uDDDZZZ��������Z}��Zb�ZtZ��Z�{�cZ������Z�{�Z��DZZZZZZZZggZ~����������tDZZZZZZZZggZZZZZZZZ���Z��������Z�����������Z��Z�Z���ZkjqphlgksspDZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZ�cZ}��bg�cZwZ}��b�cDZZZZZZZZggZZZZZZZZ�cZ}��b�cZwZ���b�{����������lZgZ�cDZZZZZZZZggZZZZZZZZ�cZ}��b�{�����ZeZ�cZZwZg}��b�cDZZZZZZZZggZZZZZZZZ�cZ}��b�cZwZkhjZgZ�d�ilhjZ��Z{|�b�cZvZ��DZZZZZZZZggZZZZZZZZ�cZ}��b�cZwZkhjZgZjhod�ddlZeZb�ddncin[Z��DZZZZZZZZggZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ��vZ{|�b�cZv|{����DZZZZZZZZggDZZZZZZZZ��������Z��ZtZ�{�ZtwZ|{����d|{����uDDZZZZZZZZ��������Z���}{�ZtZ�{�ZtwZ{|�b�cuDZZZZZZZZ��������Z�{��tZ�{�uDZZZZZZZZ��������Z���ZtZ�{�uDDZZZZ�����DZZZZZZZZggZ����Z���}{�ZvZ�{���l���DZZZZZZZZ��Z���}{�ZxZ�{���l���Z����DZZZZZZZZZZZZZZZZ���ZtwZ�����b���}{�i�{���l���cuDZZZZZZZZZZZZZZZZ���}{�ZtwZ���}{�ZgZ���d�{���l���uDZZZZZZZZ���Z��uDDZZZZZZZZ��Z���}{�ZvZjhjZ����DZZZZZZZZZZZZZZZZ������Z�{��DZZZZZZZZZZZZZZZZZZZZZZZZ������Z\���}{�ZvwZjhjZ�����Z���������Z��Z}��b�c\DZZZZZZZZZZZZZZZZZZZZZZZZ��������Z����uDZZZZZZZZZZZZZZZZ���}{�ZtwZg���}{�uDZZZZZZZZ���Z��uDDZZZZZZZZggZ}������Z�����Z���Z�������Z�����DZZZZZZZZ��Z���}{�ZwZjhjZZ��Z���}{�ZwZ�{���l���Z����DZZZZZZZZZZZZZZZZ������ZkhjuDZZZZZZZZ���Z��uDDZZZZZZZZ��ZZ���}{�ZwZ�{�����Z����DZZZZZZZZZZZZZZZZ������ZgkhjuDZZZZZZZZ���Z��uDDZZZZZZZZ��Z���}{�ZwZ�{����������lZ��Z���}{�ZwZ�{���m��������lZ����DZZZZZZZZZZZZZZZZ������ZjhjuDZZZZZZZZ���Z��uDDZZZZZZZZ���ZtwZ{|�b���}{�cuDZZZZZZZZ��ZbZ���ZvZ��cZ����DZZZZZZZZZZZZZZZZ������ZbkhjZgZjhod���d���cuDZZZZZZZZ����DZZZZZZZZZZZZZZZZ��Zb���ZvZ|{����cZ����DZZZZZZZZZZZZZZZZZZZZZZZZ������ZbkhjZgjhod���d���ZeZ���d���d���d���ilnhjcuDZZZZZZZZZZZZZZZZ���Z��uDZZZZZZZZ���Z��uDDZZZZZZZZ���ZtwZ{|�b���}{�Zg�{���l���cuDZZZZZZZZ��ZbZ���ZvZ��cZ����DZZZZZZZZZZZZZZZZ������ZbkhjZgZjhod���d���cuDZZZZZZZZ����DZZZZZZZZZZZZZZZZ��Zb���ZvZ|{����cZ����DZZZZZZZZZZZZZZZZZZZZZZZZ������ZbkhjZgjhod���d���ZeZ���d���d���d���ilnhjcuDZZZZZZZZZZZZZZZZ���Z��uDZZZZZZZZ���Z��uDDZZZZZZZZ���ZtwZ{|�Zb���}{�ZgZ�{�����cuDZZZZZZZZ��Z���ZvZ��Z����DZZZZZZZZZZZZZZZZ������ZbgkhjZeZjhod���d���cuDZZZZZZZZ����DZZZZZZZZZZZZZZZZ��Zb���ZvZ|{����cZ����DZZZZZZZZZZZZZZZZZZZZZZZZ������ZbgkhjZejhod���d���ZgZ���d���d���d���ilnhjcuDZZZZZZZZZZZZZZZZ���Z��uDZZZZZZZZ���Z��uDDZZZZZZZZggZ}������Z�����Z���Z�������Z�����DZZZZZZZZ������Z���b�{����������lZgZ���}{�cuDZZZ���Z}��uDDZZZ��������Z�{�Zb�ZtZ��Z�{�cZ������Z�{�Z��DZZZZZZZZggZ~����������tDZZZZZZZZggZZZZZZZZ���Z��������Z�����������Z��Z�Z���ZkjqphlgksspDZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZ�cZ�{�bjhjcZwZjhjDZZZZZZZZggZZZZZZZZ�cZ�{�bg�cZwZg�{�b�cDZZZZZZZZggZZZZZZZZ�cZ�������Z�{�a���Z��Z�����Z��Z�ZvZjhjDZZZZZZZZggZZZZZZZZ�cZ�������Z�{�a����Z��Z�����Z��Z�ZxZjhjDDZZZZZZZZ��������Z��{���ZtZ|���{�ZtwZ�ZvZjhjuDZZZZZZZZ��������Z���}{�ZtZ�{�ZtwZ{|�b�cZuDZZZZZZZZ��������Z�{��tZ�{�uDZZZZZZZZ��������Z���ZtZ�{�uDDZZZZ�����DZZZZZZZZggZ����ZjhjZvwZ���}{�ZvwZ�{���l���DZZZZZZZZ��Z���}{�ZxZ�{���l���Z����DZZZZZZZZZZZZZZZZ���ZtwZ�����b���}{�i�{���l���cuDZZZZZZZZZZZZZZZZ���}{�ZtwZ���}{�ZgZ���d�{���l���uDZZZZZZZZ���Z��uDDZZZZZZZZ��Z���}{�ZvZjhjZ����DZZZZZZZZZZZZZZZZ������Z�{��DZZZZZZZZZZZZZZZZZZZZZZZZ������Z\���}{�ZvwZjhjZ�����Z���������Z��Z�{�b�c\DZZZZZZZZZZZZZZZZZZZZZZZZ��������Z����uDZZZZZZZZZZZZZZZZ���}{�ZtwZg���}{�uDZZZZZZZZ���Z��uDDZZZZZZZZggZ}����Z��������Z��Z��������DZZZZZZZZ��Z���}{�ZwZ�{����������lZ����DZZZZZZZZZZZZZZZZ������Z�{��DZZZZZZZZZZZZZZZZZZZZZZZZ������Z\�Z��Z�Z��������Z��Z�{����������lZ��Z�{�b�c\DZZZZZZZZZZZZZZZZZZZZZZZZ��������Z����uDZZZZZZZZZZZZZZZZ��Z��{���Z����DZZZZZZZZZZZZZZZZZZZZZZZZ������b�{�a���cuDZZZZZZZZZZZZZZZZ����DZZZZZZZZZZZZZZZZZZZZZZZZ������b�{�a����cuDZZZZZZZZZZZZZZZZ���Z��uDZZZZZZZZ���Z��uDDZZZZZZZZ��Z���}{�ZwZ�{���m��������lZ����DZZZZZZZZZZZZZZZZ������Z�{��DZZZZZZZZZZZZZZZZZZZZZZZZ������Z\�Z��Z�Z��������Z��Z�{���m��������lZ��Z�{�b�c\DZZZZZZZZZZZZZZZZZZZZZZZZ��������Z����uDZZZZZZZZZZZZZZZZ��Z��{���Z����DZZZZZZZZZZZZZZZZZZZZZZZZ������b�{�a����cuDZZZZZZZZZZZZZZZZ����DZZZZZZZZZZZZZZZZZZZZZZZZ������b�{�a���cuDZZZZZZZZZZZZZZZZ���Z��uDZZZZZZZZ���Z��uDDZZZZZZZZggZ}������Z�����Z���Z�������Z�����DZZZZZZZZ��Z���}{�ZwZjhjZ��Z���}{�ZwZ�{�����Z����DZZZZZZZZZZZZZZZZ������ZjhjuDZZZZZZZZ���Z��uDDZZZZZZZZggZ}������Z�����Z���Z�������Z�����DZZZZZZZZ�{��ZtwZ���b���}{�ci}��b���}{�cuDZZZZZZZZ��Z��{���Z����DZZZZZZZZZZZZZZZZ������Zg�{��uDZZZZZZZZ����DZZZZZZZZZZZZZZZZ������Z�{��uDZZZZZZZZ���Z��uDZZZ���Z�{�uDDZZZ��������Z{�}���Zb�ZtZ��Z�{�ZcZ������Z�{�Z��DZZZZZZZZggZ~����������tDZZZZZZZZggZZZZZZZZ���Z��������Z�����������Z��Z�Z���ZkjqphlgksspDZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZ�cZ{�}���bg�cZwZg{�}���b�cDZZZZZZZZggZZZZZZZZ�cZ�������Z�Z��Z�����DDZZZZZZZZ��������Z��{���ZtZ|���{�ZtwZ�ZvZjhjuDZZZZZZZZ��������Z���}{�ZtZ�{�ZtwZ{|�b�cuDZZZZZZZZ��������Z�{��ZtZ�{�uDDZZZ�����DZZZZZZggZ}����Z��������Z��Z���������DZZZZZZ��Z���}{�ZxZkhjZ����DZZZZZZZZZ������Z�{��DZZZZZZZZZZZZZZZZ������Z\{|�b�cZxZkhjZ��Z{�}���b�c\DZZZZZZZZZZZZZZZZ��������Z����uDZZZZZZZZZ������Z�uDZZZZZZ���Z��uDDZZZZZZggZ}������Z�����Z���Z�������Z�����DZZZZZZ��Z���}{�ZwZjhjZ����DZZZZZZZZZ������ZjhjuDZZZZZZ�����Z���}{�ZwZkhjZ����DZZZZZZZZZ��Z��{���Z����DZZZZZZZZZZZZZZZZ������Zg�{����������luDZZZZZZZZZ����DZZZZZZZZZZZZZZZZ������Z�{����������luDZZZZZZZZZ���Z��uDZZZZZZ���Z��uDDZZZZZZggZ}������Z�����Z���Z�������Z�����DZZZZZZ��Z���}{�ZvZjhsZ����DZZZZZZZZZ�{��ZtwZ{�}�{�b���}{�ib����bkhjZgZ���}{�d���}{�cccuDZZZZZZ����DZZZZZZZZZ�{��ZtwZ�{����������lZgZ{�}�{�b����bkhjZgZ���}{�d���}{�ci���}{�cuDZZZZZZ���Z��uDDZZZZZZ��Z��{���Z����DZZZZZZZZZ�{��ZtwZg�{��uDZZZZZZ���Z��uDDZZZZZZ������Z�{��uDZZZ���Z{�}���uDDZZZ��������Z{�}}��Zb�ZtZ��Z�{�cZ������Z�{�Z��DZZZZZZZZggZ~����������tDZZZZZZZZggZZZZZZZZ���Z��������Z�����������Z��Z�Z���ZkjqphlgksspDZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZ�cZ{�}}��bg�cZwZ�{�����ZgZ{�}}��b�cDZZZZZZZZggZZZZZZZZ�cZ�������Z�Z��Z�����DDZZZZZZZZ��������Z��{���ZtZ|���{�ZtwZ�ZvZjhjuDZZZZZZZZ��������Z���}{�ZtZ�{�ZtwZ{|�b�cuDZZZZZZZZ��������Z�{��ZtZ�{�uDDZZZ�����DZZZZZZggZ}����Z��������Z��Z��������DZZZZZZ��Z���}{�ZxZkhjZ����DZZZZZZZZZ������Z�{��DZZZZZZZZZZZZZZZZ������Z\{|�b�cZxZkhjZ��Z{�}}��b�c\DZZZZZZZZZZZZZZZZ��������Z����uDZZZZZZZZZ������Z�uDZZZZZZ���Z��uDDZZZZZZggZ}������Z�����Z���Z�������Z�����DZZZZZZ��Z�ZwZkhjZ����DZZZZZZZZZ������ZjhjuDZZZZZZ�����Z�ZwZjhjZ����DZZZZZZZZZ������Z�{����������luDZZZZZZ�����Z�ZwZgkhjZ����DZZZZZZZZZ������Z�{�����uDZZZZZZ���Z��uDDZZZZZZggZ}������Z�����Z���Z�������Z�����DZZZZZZ��Z���}{�ZxZjhsZ����DZZZZZZZZZ�{��ZtwZ{�}�{�b����bkhjZgZ���}{�d���}{�ci���}{�cuDZZZZZZ����DZZZZZZZZZ�{��ZtwZ�{����������lZgZ{�}�{�b���}{�i����bkhjZgZ���}{�d���}{�ccuDZZZZZZ���Z��uDDDZZZZZZ��Z��{���Z����DZZZZZZZZZ�{��ZtwZ�{�����ZgZ�{��uDZZZZZZ���Z��uDDZZZZZZ������Z�{��uDZZZ���Z{�}}��uDDDZZZ��������Z{�}�{�Zb�ZtZ��Z�{�cZ������Z�{�Z��DZZZZZZZZggZ~����������tDZZZZZZZZggZZZZZZZZ���Z��������Z�����������Z��Z�Z���ZkjqphlgksspDZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZ�cZ{�}�{�bg�cZwZg{�}�{�b�cDZZZZZZZZggZZZZZZZZ�cZ{�}�{�b�cZwZg{�}�{�bkhji�cZeZ�{����������lZ���Z���ZxZkhjDZZZZZZZZggZZZZZZZZ�cZ{�}�{�b�cZwZ�Z���Z���ZvZ��DDZZZZZZZZ��������Z��ZtZ�{�ZtwZ|{����d|{����d|{����uDDZZZZZZZZ��������Z��{���ZtZ|���{�ZtwZ�ZvZjhjuDZZZZZZZZ��������Z�}����}{�ZtZ|���{�uDZZZZZZZZ��������Z���}{�ZtZ�{�ZtwZ{|�b�cuDZZZZZZZZ��������Z�{��ZtZ�{�uDDZZZ�����DZZZZZZggZ����Z��������Z���ZvwkhjDZZZZZZ��Z���}{�ZxZkhjZ����DZZZZZZZZZZZZZZZZ���}{�ZtwZkhji���}{�uDZZZZZZZZZZZZZZZZ�}����}{�ZtwZ���uDZZZZZZ����DZZZZZZZZZZZZZZZZ�}����}{�ZtwZ�{��uDZZZZZZ���Z��uDDZZZZZZggZ}������Z�����Z���Z�������Z�����DZZZZZZ��Z���}{�ZwZjhjZ����DZZZZZZZZZ��Z�}����}{�Z����DZZZZZZZZZZZZZZZZ��Z��{���Z����DZZZZZZZZZZZZZZZZZZZZZZZZ������Zbg�{����������lcuDZZZZZZZZZZZZZZZZ����DZZZZZZZZZZZZZZZZZZZZZZZZ������Zb�{����������lcuDZZZZZZZZZZZZZZZZ���Z��uDZZZZZZZZZ����DZZZZZZZZZZZZZZZZ������ZjhjuDZZZZZZZZZ���Z��uDZZZZZZ���Z��uDDZZZZZZ��Z���}{�ZvZ��Z����DZZZZZZZZZ��Z��{���Z����DZZZZZZZZZZZZZZZZ��Z�}����}{�Z����DZZZZZZZZZZZZZZZZZZZZZZZZ������Zbg�{����������lZeZ���}{�cuDZZZZZZZZZZZZZZZZ����DZZZZZZZZZZZZZZZZZZZZZZZZ������Zg���}{�uDZZZZZZZZZZZZZZZZ���Z��uDZZZZZZZZZ����DZZZZZZZZZZZZZZZZ��Z�}����}{�Z����DZZZZZZZZZZZZZZZZZZZZZZZZ������Zb�{����������lZgZ���}{�cuDZZZZZZZZZZZZZZZZ����DZZZZZZZZZZZZZZZZZZZZZZZZ������Z���}{�uDZZZZZZZZZZZZZZZZ���Z��uDZZZZZZZZZ���Z��uDZZZZZZ���Z��uDDZZZZZZggZ}������Z�����Z���Z�������Z�����DZZZZZZ�{��ZtwZZ}��~�}bZkhjfZ���}{�fZjhjfZlqfZ�}������ZcblcuDDZZZZZZ��Z�}����}{�Z����DZZZZZZZZZ�{��ZtwZ�{����������lZgZ�{��uDZZZZZZ���Z��uDDZZZZZZ��Z��{���Z����DZZZZZZZZ�{��ZtwZg�{��uDZZZZZZ���Z��uDDZZZZZZ������Z�{��uDZZZ���Z{�}�{�uDDDZZZ��������Z{�}�{�Zb�ZtZ��Z�{�uZ�ZtZ��Z�{�cZ������Z�{�Z��DZZZZZZZZggZ~����������tDZZZZZZZZggZZZZZZZZ���Z��������Z�����������Z��Z�Z���ZkjqphlgksspDZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZZ�cZ�������ZjhjZ��Z�����DDZZZZZZZZ��������Z���}{�ZtZ�{�uDZZZZZZZZ��������Z�{��ZtZ�{�uDZZZ�����DDZZZZZggZ}����Z��������Z��Z���������DZZZZZ��Zb�ZwZjhjZ���Z�ZwZjhjZcZ����DZZZZZZZZZZZ������Z�{��Z������DZZZZZZZZZZZZZZZZ\{�}�{�bjhjfZjhjcZ��Z������������\DZZZZZZZZZZZZZZZZ��������Z����uDZZZZZZZZZZZ������ZjhjuDZZZZZ���Z��uDDZZZZZggZ}������Z�����Z���Z�������Z�����DZZZZZ��Z�ZwZjhjZ����DZZZZZZZZ��Z�ZxZjhjZ����DZZZZZZZZZZZ������ZjhjuDZZZZZZZZ����DZZZZZZZZZZZ������Z�{�����uDZZZZZZZZ���Z��uDZZZZZ���Z��uDDZZZZZ��Z�ZwZjhjZ����DZZZZZZZZ��Z�ZxZjhjZ����DZZZZZZZZZZZ������Z�{����������luDZZZZZZZZ����DZZZZZZZZZZZ������Zg�{����������luDZZZZZZZZ���Z��uDZZZZZ���Z��uDDDZZZZZggZ}������Z�����Z���Z�������Z�����DZZZZZ���}{�ZtwZ{|�b�i�cuDDZZZZZ�{��ZtwZ{�}�{�b���}{�cuDDZZZZZ��Z�ZvZjhjZ����DZZZZZZZZZ�{��ZtwZ�{�����ZgZ�{��uDZZZZZ���Z��uDDZZZZZ��Z�ZvZjhjZ����DZZZZZZZZZ�{��ZtwZg�{��uDZZZZZ���Z��uDDZZZZZ������Z�{��uDZZZ���Z{�}�{�uDDDZZZZ��������Z����Zb�ZtZ��Z�{�cZ������Z�{�Z��DZZZZZZZZggZ~����������tDZZZZZZZZggZZZZZZZZ���Z��������Z�����������Z��Z�Z���ZkjqphlgksspDZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZ�cZ�������Zb��b�cZgZ��bg�ccilhjDZZZZZZZZggZZZZZZZZ�cZ����bg�cZwZ����b�cDDZZZZZZZZ��������Z��{���ZtZ|���{�ZtwZ�ZvZjhjuDZZZZZZZZ��������Z���}{�ZtZ�{�ZtwZ{|�b�cuDZZZZZZZZ��������Z���ZtZ�{�uDZZZZZZZZ��������Z�{��ZtZ�{�uDDZZZZ�����DZZZZZZZZggZ}������Z�����Z���Z�������Z�����DZZZZZZZZ��Z���}{�ZwZjhjZ����DZZZZZZZZZZZZZZZZ������ZjhjuDZZZZZZZZ���Z��uDDZZZZZZZZggZ}������Z�����Z���Z�������Z�����DZZZZZZZZ���ZtwZ��b���}{�cuDZZZZZZZZ�{��ZtwZb���ZgZkhji���cdjhouDDZZZZZZZZZ��Z��{���Z����DZZZZZZZZZZZZZZZZ�{��ZtwZg�{��uDZZZZZZZZ���Z��uDDZZZZZZZZ������Z�{��uDZZZZ���Z����uDDZZZZ��������ZZ}���Zb�ZtZ��Z�{�cZ������Z�{�Z��DZZZZZZZZggZ~����������tDZZZZZZZZggZZZZZZZZ���Z��������Z�����������Z��Z�Z���ZkjqphlgksspDZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZ�cZ�������Zb��b�cZeZ��bg�ccilhjDZZZZZZZZggZZZZZZZZ�cZ}���bg�cZwZ}���b�cDDZZZZZZZZ��������Z���}{�ZtZ�{�ZtwZ{|�b�cuDZZZZZZZZ��������Z���ZtZ�{�uDZZZZZZZZ��������Z�{��ZtZ�{�uDZZZZ�����DZZZZZZZZggZ}������Z�����Z���Z�������Z�����DZZZZZZZZ��Z���}{�ZwZjhjZ����DZZZZZZZZZZZZZZZZ������ZkhjuDZZZZZZZZ���Z��uDDDZZZZZZZZggZ}������Z�����Z���Z�������Z�����DZZZZZZZZ���ZtwZ��b���}{�cuDZZZZZZZZ�{��ZtwZb���ZeZkhji���cdjhouDDZZZZZZZZ������Z�{��uDZZZZ���Z}���uDDZZZZ��������ZZ�{��Zb�ZtZ��Z�{�cZ������Z�{�Z��DZZZZZZZZggZ~����������tDZZZZZZZZggZZZZZZZZ���Z��������Z�����������Z��Z�Z���ZkjqphlgksspDZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZ�cZ�������Zb��b�cZgZ��bg�ccib��b�cZeZ��bg�ccDZZZZZZZZggZZZZZZZZ�cZ�{��bg�cZwZg�{��b�cDDZZZZZZZZ��������Z��{���ZtZ|���{�ZtwZ�ZvZjhjuDZZZZZZZZ��������Z���}{�ZtZ�{�ZtwZ{|�b�cuDZZZZZZZZ��������Z���ZtZ�{�uDZZZZZZZZ��������Z�{��ZtZ�{�uDDZZZZ�����DZZZZZZZZggZ}������Z�����Z���Z�������Z�����DZZZZZZZZ��Z���}{�ZwZjhjZ����DZZZZZZZZZZZZZZZZ������ZjhjuDZZZZZZZZ���Z��uDDZZZZZZZZggZ}������Z�����Z���Z�������Z�����DZZZZZZZZ���ZtwZ��b���}{�cuDZZZZZZZZ�{��ZtwZb���ZgZkhji���cib���ZeZkhji���cuDDZZZZZZZZ��Z��{���Z����DZZZZZZZZZZZZ������Zg�{��uDZZZZZZZZ����DZZZZZZZZZZZZ������Z�{��uDZZZZZZZZ���Z��uDZZZZ���Z�{��uDDZZZZ��������Z{�}����Zb�ZtZ��Z�{�cZ������Z�{�Z��DZZZZZZZZggZ~����������tDZZZZZZZZggZZZZZZZZ���Z��������Z�����������Z��Z�Z���ZkjqphlgksspDZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZ�cZ�������Z���bZ�ZeZ����bZ�d�ZeZkhjccDDZZZZ�����DZZZZZZZZggZ}������Z�����Z���Z�������Z�����DZZZZZZZZ��Z�ZwZjhjZ����DZZZZZZZZZZZZZZZZ������ZjhjuDZZZZZZZZ���Z��uDDZZZZZZZZggZ}������Z�����Z���Z�������Z�����DZZZZZZZZ������ZbZ���bZ�ZeZ����bZ�d�ZeZkhjccZcuDZZZZ���Z{�}����uDDDDZZZ��������Z{�}}���Zb�ZtZ��Z�{�cZ������Z�{�Z��DZZZZZZZZggZ~����������tDZZZZZZZZggZZZZZZZZ���Z��������Z�����������Z��Z�Z���ZkjqphlgksspDZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZ�cZ�������Z���bZ�ZeZ����bZ�d�ZgZkhjccuZZZ�ZxwZkhjDZZZZZZZZggZZZZZZZZ�cZ�������Z�Z��Z�����DDZZZZ�����DZZZZZZZZggZ}����Z��������Z��Z���������DZZZZZZZZ��Z�ZvZkhjZ����DZZZZZZZZZZZZZZZZZ������Z�{��DZZZZZZZZZZZZZZZZZZZZZZZZ������Z\�ZvZkhjZ��Z{�}}���b�c\DZZZZZZZZZZZZZZZZZZZZZZZZ��������Z����uDZZZZZZZZZZZZZZZZZ������Z�uDZZZZZZZZ���Z��uDDZZZZZZZZggZ}������Z�����Z���Z�������Z�����DZZZZZZZZ��Z�ZwZkhjZ����DZZZZZZZZZZZZZZZZ������ZjhjuDZZZZZZZZ���Z��uDDZZZZZZZZggZ}������Z�����Z���Z�������Z�����DZZZZZZZZ������ZbZ���bZ�ZeZ����bZ�d�ZgZkhjcccuDZZZZ���Z{�}}���uDDZZZZ��������Z{�}�{��Zb�ZtZ��Z�{�cZ������Z�{�Z��DZZZZZZZZggZ~����������tDZZZZZZZZggZZZZZZZZ���Z��������Z�����������Z��Z�Z���ZkjqphlgksspDZZZZZZZZggZ�����tDZZZZZZZZggZZZZZZZZ�cZ�������Zb���bZbkhjZeZ�cibkhjZgZ�cccilhjZuZ�Z�Z�ZvZkhjDZZZZZZZZggZZZZZZZZ�cZ�������Z�Z��Z�����DZZZZ�����DZZZZZZZZggZ}����Z��������Z��Z���������DZZZZZZZZ��Z{|�b�cZxwZkhjZ����DZZZZZZZZZZZZZZZZ������Z�{��DZZZZZZZZZZZZZZZZZZZZZZZZ������Z\{|�b�cZxwZkhjZ��Z{�}�{��b�c\DZZZZZZZZZZZZZZZZZZZZZZZZ��������Z����uDZZZZZZZZZZZZZZZZ������Z�uDZZZZZZZZ���Z��uDDZZZZZZZZggZ}������Z�����Z���Z�������Z�����DZZZZZZZZ��Z�ZwZjhjZ����DZZZZZZZZZZZZZZZZ������ZjhjuDZZZZZZZZ���Z��uDDZZZZZZZZggZ}������Z�����Z���Z�������Z�����DZZZZZZZZ������bZjhod���bZbkhje�cibkhjg�cZcZcuDZZZZ���Z{�}�{��uDD���ZZ�{����{�uD