--
@ER--B$FbsEHo0OR52gR4g-cRRj.jd$R1MHbDO$H0ROQM
R--fN]C8:CsR#//$DMbH0OH$N/lb0DN.Uj4J4.b/blNb#Cs/0N0/LDH/MoC_OFsN/6ol0kD38PEyf4R

--
-
-R****************************************************************-RR--
-R#zMHCoM8kRvDb0HDsHC
R--aoNsC:0RR0pN0CHOROmsN
R6-N-RsDOEHR#0=FRDoRHOLODF	k_lD-0
-3R4RoDFH-ORRsNsNl$RkHD0bCDHsHRI0bERHLbCkRV#5RHMOCN#RRFVbCHbDHHMM
o2---
-3R.RFLDO-	RRHk#MmoRsRON6DRAFRO	v0kDHHbDC5sRvazp44UXU-2
--
-RFRBbH$soRE05RO2.jjj,jR.j14R$DMbH0OH$Q,RM
O3-R-RqRDDsEHo0s#RCs#CP3C8
R--****************************************************************R-R-
-
-R****************************************************************-RR--
-RswH#s0uFO8k0q#5,,RAR2qA

---W-RHE80qRR-I0H8EVRFRHqRM0bk
R--W0H8E-ARR8IH0FERVRRAHkMb0-
-R-
-RRqA-HRL0HIN#qCRhF7RVDRNDMRHb#k0
R--
R--****************************************************************R-R-
H
DLssN$CRHCRC;
Ck#RCHCC03#8F_Do_HO4c4n3DND;D

HNLss#$R$DMbH;V$
Ck#RM#$bVDH$03N0LsHk#0C3DND;D

HNLssF$RsdON;#
kCsRFO3NdFNsOObFl3DND;D

HNLss#$R$DMbH;V$
Ck#RM#$bVDH$03N0LsHk#0C3DND;C

M00H$HRwsu#0skF8OR0#HR#
RCRoMHCsOR5
RRRRR8IH0REq:MRH0CCosR;
RRRRR8IH0REA:MRH0CCosR
RR
2;RbRRFRs05R
RRRRRq:RRRRHMR8#0_oDFHPO_CFO0sH5I8q0E-84RF0IMF2Rj;R
RRRRRA:RRRRHMR8#0_oDFHPO_CFO0sH5I8A0E-84RF0IMF2Rj;R
RRRRRq:ARR0FkR8#0_oDFHPO_CFO0sH5I8A0E*8IH0-Eq4FR8IFM0R
j2RRRRR-R-R*ARRRq
R;R2
8CMRswH#s0uFO8k0
#;
ONsECH0Os0kCsRNORE4FwVRH0s#u8sFk#O0R
H#
RRR#MHoNNDR_GNkR#:R0D8_FOoH_OPC05FsI0H8E4q-RI8FMR0Fj
2;R#RRHNoMD_RLNRkG:0R#8F_Do_HOP0COFIs5HE80AR-48MFI0jFR2
;
LHCoMR
RRsVFqqM8:FRVsNRHRRHMjFR0R8IH0-Eq4CRoMNCs0RC
RRRRRsVFqAM8:FRVsLRHRRHMjFR0R8IH0-EA4CRoMNCs0RC
RRRRRRRRqIA5HE80AN*HRH+RL<2R=5RqHRN2qRh7AL5H2R;
RRRRR8CMRMoCC0sNCFRVs8qMAR;
RMRC8CRoMNCs0VCRFMsq8
q;CRM8NEsO4
;
-*-R*************************************************************R**R
---N-R8C8so,5qRRA,)2C#

---v-RF#PCRosCHC#0s0#RFCRsbODNCHRbbkCLV
'#-
-R-*-R*************************************************************R**R
--
LDHs$NsRCHCC
;RkR#CHCCC38#0_oDFH4O_43ncN;DD
Ck#RCHCC03#8F_Do_HOkHM#o8MC3DND;D

HNLss#$R$DMbH;V$
Ck#RM#$bVDH$03N0LsHk#0C3DND;D

HNLssF$RsdON;#
kCsRFO3NdFNsOObFl3DND;C

M00H$8RN8osCR
H#RoRRCsMCH
O5RRRRRHRI8R0E:MRH0CCosR;
RRRRRosCR:RRR0HMCsoCRR--hCNlRRFV0RECDCCPDR
RR
2;RbRRFRs05R
RRRRRqRRR:MRHR8#0_oDFHPO_CFO0sH5I8-0E4FR8IFM0R;j2
RRRRARRR:RRRRHM#_08DHFoOC_POs0F58IH04E-RI8FMR0Fj
2;RRRRRCR)#RR:FRk0#_08DHFoOC_POs0F58IH04E-RI8FMR0FjR2
R;R2
RRRNs00H0LkC3R\s	NM\RR:HCM0o;Cs
RRRNs00H0LkC3R\sFClPMC_FN_IsRM\:MRH0CCosC;
MN8R8C8so
;
NEsOHO0C0CksRONsEF4RV8RN8osCR
H#
RRR#MHoN)DRCD#k0RR:#_08DHFoOC_POs0F58IH04E-RI8FMR0Fj
2;
oLCHRM
RCR)#0kDRR<=qRR+AR;
RFRVsFDFbR.:VRFsHMRHR0jRFHRI8-0E4CRoMNCs0RC
RRRRR0N0skHL0\CR3MsN	F\RVCRso:#RRLDNCHDR#CRsoS;
S0N0skHL0\CR3lsCF_PCMIF_N\sMRRFVs#CoRD:RNDLCRRH#4R;
RCRLo
HMRRRRRCRsoR#:bCHbL
kVRRRRRFRbsl0RN
b5RRRRRRRRR=QR>CR)#0kD5,H2
RRRRRRRRRRm=)>RCH#52R
RRRRR2R;
RMRC8CRoMNCs0VCRFFsDF;b.
8CMRONsE
4;
R--****************************************************************R-R-

---V-RDsFF5bQMkR0,mbk0k
02---
-*R**************************************************************R*R-
-
DsHLNRs$HCCC;kR
#HCRC3CC#_08DHFoO4_4nNc3D
D;
LDHs$NsROFsN
d;kR#CFNsOds3FOFNOlNb3D
D;
M
C0$H0RFVDFHsR#R
RRMoCCOsHRR5
RRRRR8IH0hEQRRR:HCM0oRCs:d=RcR;
RRRRR8IH0zEmaRR:HCM0oRCs:d=RcR;
RRRRRlMkLRCsRRR:HCM0oRCs:4=R;R
RRRRRHCM8GRRRRH:RMo0CC:sR=R4
R;R2
RRRb0FsRR5
RRRRRbQMkR0R:HRRM0R#8F_Do_HOP0COFIs5HE80Q4h-RI8FMR0Fj
2;RRRRRkRm00bkRF:Rk#0R0D8_FOoH_OPC05FsI0H8Eamz-84RF0IMF2Rj
RRR2R;
R0RN0LsHkR0C\N3sMR	\:MRH0CCosR;
R0RN0LsHkR0C\C3slCFP__MFIMNs\RR:HCM0o;Cs
8CMRFVDF
s;
ONsECH0Os0kCsRNORE4FVVRDsFFRRH#
R
RRR--)HCo#s0CRlBFbCFMMR0
RFROlMbFCRM0Ns88CRo
RRRRRMoCCOsHRR5
RRRRRRRRI0H8ERR:HCM0o;Cs
RRRRRRRRCRsoRRR:MRH0CCos-R-RlhNCVRFRC0ERPDCCRD
RRRRR
2;RRRRRFRbs50R
RRRRRRRRRRqRRR:H#MR0D8_FOoH_OPC05FsR8IH04E-RI8FMR0Fj
2;RRRRRRRRRRARRH:RM0R#8F_Do_HOP0COFRs5I0H8ER-48MFI0jFR2R;
RRRRRRRR)RC#:kRF00R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj
RRRR2RR;R
RR8CMRlOFbCFMM
0;
RRR#MHoN)DRCD#k0RR:#_08DHFoOC_POs0F58IH0hEQ-84RF0IMF2Rj;R

R-R-RMVkOF0HMsROCCN0#RRNl0kDHHbDC0sRFER#HRV0NNRPDRkCD0CVRRL$HCM8GHRL0
#
RVRRk0MOHRFM#VEH0sxCFM5H8RCG:MRH0CCoss2RCs0kMMRH0CCos#RH
RRRRPRRNNsHLRDC#b0CRH:RMo0CC
s;RLRRCMoH
RRRR#RR0RCb:4=R;R
RRRRRVRFsHMRHR04RFMRH8-CG4FRDFRb
RRRRRRRR#b0CRR:=#b0CR.*R;R
RRRRRCRM8DbFF;R
RRRRRskC0s#MR0;Cb
RRRCRM8#VEH0sxCF
;
RORRF0M#NRM0#VEH08N8C:sRR0HMCsoCRR:=#VEH0sxCFM5H82CG;R
RRMOF#M0N0CRDMEo0RRRRRH:RMo0CC:sR=HRI8Q0EMk/MlsLC;-

--R
-sRNO0EHCkO0sFCRVDRVFRFs-MRFCHRbbHCDMRC8#o0NC-
-RL

CMoHRR
RRsVFDbFF_R4:VRFs[MRHR04RFkRMlsLC/o.RCsMCN
0CRLRRCMoH
RRRRsRRCqo#:8RN8osC
RRRRoRRCsMCHlORN5bR
RRRRRRRRHRI8R0E=D>RC0MoEE-#HNV08s8C,R
RRRRRRsRRCRoRRR=>HCM8GR
RRRRR2R
RRRRRb0FsRblN5R
RRRRRRqRRRR=>QkMb0C5DMEo0**5.[2-4-84RF0IMFCRDMEo0*5.*[2-4+H#EV80N82Cs,R
RRRRRRARRRR=>QkMb0C5DMEo0*[.*-84RF0IMFCRDMEo0**5.[2-4+H#EV80N82Cs,R
RRRRRR)RRC=#R>kRm00bk5MDCo*0E[R-48MFI0DFRC0MoE[*5-+42#VEH08N8C
s2RRRRR;R2
RRRRVRRFFsDF.b_:FRVsRR	HjMRRR0F#VEH08N8C4s-RMoCC0sNCR
RRRRRRNRR0H0sLCk0Rs\3N\M	RRFVs#CoRD:RNDLCRRH#HCM8GS;
S0SN0LsHkR0C\C3slCFP__MFIMNs\VRFRosC#RR:DCNLD#RHR
4;RRRRRCRLo
HMRRRRRRRRRR--mbk0kD05C0MoE[*5-+42#VEH08N8C4s-RI8FMR0FDoCM05E*[2-42=R<RR
RRRRRR-RR-RRRRbQMkD05C0MoE**.54[-2E+#HNV08s8C-84RF0IMFCRDMEo0*5.*[2-42R;
RRRRRRRRs#Co:bRRHLbCkRV
RRRRRRRRb0FsRblN5R
RRRRRRRRRRRRQ=Q>RM0bk5MDCo*0E.[*5-+42	
2,RRRRRRRRRRRRm>R=R0mkb5k0DoCM05E*[2-4+
	2RRRRRRRRR
2;RRRRRMRC8CRoMNCs0VCRFFsDF.b_;R
RR8CMRMoCC0sNCFRVsFDFb;_4
R
RR_HV##FkNH:RVMR5kClLsFRl8RR.=2R4RMoCC0sNCR
RRoLCHRM
RRRRRV--FFsDFdb_:FRVsRRHH4MRRR0FDoCM0#E-E0HVNC88sCRoMNCs0RC
RRRRRsVFDbFF_Rd:VRFsHMRHR04RFCRDMEo0RMoCC0sNCS
SS0N0skHL0\CR3MsN	F\RVCRso:#RRLDNCHDR#MRH8;CG
SSSNs00H0LkC3R\sFClPMC_FN_IsRM\FsVRCRo#:NRDLRCDH4#R;R
RRRRRLHCoMR
RRRRRRsRRC:o#RHRbbkCLVR
RRRRRRbRRFRs0l5Nb
RRRRRRRRRRRR=QR>MRQb5k0I0H8E-QhH
2,RRRRRRRRRRRRm>R=R0mkb5k0I0H8Eamz-
H2RRRRRRRRR
2;RRRRRMRC8CRoMNCs0VCRFFsDFdb_;R
RRRRR-m-Rkk0b0H5I8m0Ez#a-E0HVNC88sR-48MFI0IFRHE80m-zaDoCM0RE2
RRRR-RR-RRRRR<=QkMb0H5I8Q0EhE-#HNV08s8C-84RF0IMFHRI8Q0EhC-DMEo02R;
RMRC8CRoMNCs0HCRVF_#k;#N
8CMRONsE
4;
R--****************************************************************R-R-
R--
R--NC88sCasCW5RHE80qW,RHE80A-2
--R
-*R**************************************************************R*R-
-
DsHLNRs$HCCC;kR
#HCRC3CC#_08DHFoO4_4nNc3D
D;kR#CHCCC38#0_oDFHNO_sEH03DND;#
kCCRHC#C30D8_FOoH_#kMHCoM8D3ND
;
CHM00N$R8s8CaCsCR
H#RoRRCsMCH
O5RRRRRHRI8q0ERH:RMo0CC
s;RRRRRHRI8A0ERH:RMo0CCRs
R;R2
RRRb0FsRR5
RRRRRRqARRRRRH:RM0R#8F_Do_HOP0COFIs5HE80AH*I8q0E-84RF0IMF2Rj;R
RRRRRb8sFkRO0:kRF00R#8F_Do_HOP0COFIs5HE80AH+I8q0E-84RF0IMF2Rj
RRRR-RR-RRA*
RqR2RR;M
C88RN8aCss;CC
NR
sHOE00COkRsCNEsO4VRFR8N8CssaCHCR#R

RFROMN#0M00REHCEo:ERR8#0_oDFHPO_CFO0s654RI8FMR0Fj:2R=mRBh1e_ap7_mBtQ_Be a5m)I0H8E4q-,nR42
;
RORRFFlbM0CMRFVDFRs
RRRRRMoCCOsHRR5
RRRRRRRRI0H8ERQhRH:RMo0CC;sR
RRRRRRRRHRI8m0Ez:aRR0HMCsoCRR;
RRRRRRRRMLklCRsRRH:RMo0CC;sR
RRRRRRRRMRH8RCGR:RRR0HMCsoC
RRRR2RR;R
RRRRRb0FsRR5
RRRRRRRRQkMb0:RRRRHM#_08DHFoOC_POs0F58IH0hEQ-84RF0IMF2Rj;R
RRRRRRmRRkk0b0RR:FRk0#_08DHFoOC_POs0F58IH0zEmaR-48MFI0jFR2R
RRRRR2R;
RMRC8FROlMbFC;M0
-
-RMVH8ER0CFRDOHN0FFMRVER0CHREo#EC04R''MRHRE"0CoEHE
"
RVRRk0MOHRFM80CbE8WH0sERCs0kMMRH0CCos#RH
RRRLHCoMR
RRRRRVRFsHMRHRR468MFI0jFRRFDFbR
RRRRRRHRRV0R5EHCEoHE52RR='24'RC0EMR
RRRRRRRRRRsRRCs0kM+RH4R;
RRRRRRRRCRM8H
V;RRRRRMRC8FRDF
b;RRRRRCRs0MksR
j;RCRRM88RCEb0W0H8E
;
RORRF0M#NRM080CbE:RRR0HMCsoCRR:=80CbE8WH0
E;RORRF0M#NRM0I0H8ERR:HCM0oRCs:I=RHE80AH+I8q0E+
4;R0RR$RbCD#HlRRH#NNss$8R5CEb0+84RF0IMF2RjRRFVHCM0o;Cs
-R
-HRVM08REsCRCHJksRC8MLklCRs#5C0E_lMkL#CsRRHMNNMRs$sNRRFVHCM0o#Cs2R

RkRVMHO0FOMRNhDOkClLss#RCs0kMHRDlH#R#R
RRRRRPHNsNCLDRC0E_lMkL#CsRD:RH;l#
RRRLHCoMR
RRRRR0_ECMLklC5s#j:2R=HRI8q0E;R
RRRRRVRFsHMRHR04RFCR8b+0E4FRDFRb
RRRRRRRR0_ECMLklC5s#H:2R=ER0Ck_MlsLC#-5H4.2/R5+R0_ECMLklC5s#H2-4R8lFR;.2
RRRRCRRMD8RF;Fb
RRRRsRRCs0kMER0Ck_MlsLC#R;
RCRRMO8RNhDOkClLs
#;RR
RRMOF#M0N0kRMlsLC#RR:D#HlRR:=OONDhLklC;s#
-R
-NRODDOkNR0C0_ECD#Hl
R
RRMVkOF0HMNRODHOplCRs0MksRlDH##RH
RRRRPRRNNsHLRDC0_ECD#HlRD:RH;l#
RRRRPRRNNsHLRDCMLklRRRRRH:RMo0CC
s;RLRRCMoH
RRRR0RREDC_H5l#j:2R=;Rj
RRRRMRRkRlL:I=RHE80qR;
RRRRRsVFRHHRMRR408FRCEb0+D4RF
FbRRRRRRRRRC0E_lDH#25HRR:=0_ECD#Hl54H-2RR+MLkl*8IH0
E;RRRRRRRRRlMkL=R:RlMkLR/.+MR5kRlLlRF8.
2;RRRRRMRC8FRDF
b;RRRRRCRs0MksRC0E_lDH#R;
RMRC8NRODHOplR;

RRRO#FM00NMROPCDRHl:HRDl:#R=NRODHOplR;
RHR#oDMNRHRLoC0sCRR:#_08DHFoOC_POs0F5OPCD5Hl80CbE2+4-84RF0IMF2Rj;-

-sROCCN0RC0ERONsECH0Os0kCVRFRC0ER8N8C0sRs
CC
oLCH
MRRVRRFMsN8Rq:VRFsHHNRMRRj0IFRHE80qR-4oCCMsCN0
RRRRLRRHso0C5C5H4N+2H*I8-0E4FR8IFM0R*HNI0H8E<2R=BRRm_he1_a7pQmtB _eB)am5Rj,I0H8EHq-N2+4
RRRRRRRRRR&qIA5HE80AH*5N2+4-84RF0IMFHRI8A0E*2HN
RRRRRRRRRR&Bemh_71a_tpmQeB_ mBa),5jR2HN;R
RR8CMRMoCC0sNCFRVs8NMq
;
RVRRFFsDF:b.VRFs[MRHR04RFCR8bR0EoCCMsCN0
RRRlR4:RFVDFRs
RRRRRMoCCOsHRblNRR5
RRRRRRRRI0H8ERQhRR=>PDCOH[l52RR-PDCOH[l5-,42
RRRRRRRRHRI8m0Ez=aR>CRPOlDH54[+2RR-PDCOH[l52R,
RRRRRRRRMLklCRsRRR=>MLklC5s#[2-4,R
RRRRRRHRRMG8CRRRR=[>R
RRRRRRRR
R2RRRRRFRbsl0RN5bR
RRRRRRRRMRQbRk0R=RR>HRLoC0sCC5POlDH5-[24FR8IFM0ROPCD5Hl[2-42R,
RRRRRRRRmbk0kR0RRR=>L0Hos5CCPDCOH[l5+-424FR8IFM0ROPCD5Hl[
22RRRRR;R2
RRRCRM8RMoCC0sNCFRVsFDFb
.;
RRRb8sFkRO0<L=RHso0CPC5CHODlC58b+0E4.2-RI8FMR0FPDCOH8l5CEb02R2;
M
C8sRNO;E4
-
-R****************************************************************-
-RCaER#kMHCoM8kRlDb0HDk$R#RC#vazp44(G(-
-R****************************************************************D

HNLssQ$R ;  
Ck#RCHCC03#8F_Do_HO4c4n3DND;#
kCCRHC#C30D8_FOoH_HNs0NE3D
D;kR#CHCCC38#0_oDFH#O_HCoM8D3ND
;
CHM00v$Rz4pa((X4R
H#SR
RRsbF0
R5RRRRRRRq:MRHR0R#8F_Do_HOP0COF4s5nFR8IFM0R;j2
RRRRARRRH:RM#RR0D8_FOoH_OPC05Fs48nRF0IMF2Rj;R
RRRRRuRR:FRk0#_08DHFoOC_POs0F5Rdd8MFI0jFR2S
S2
;
RNRR0H0sLCk0RH\3Ms0CM_NDH0M#NHM0N80C\RR:HCM0o;Cs
8CMRpvzaX4(4
(;
R--#0$MEHC##sR0NDM#N_0CF
VV-D-RHNLss#$RHslbH
l;-k-R##CRHslbHel3b	NON3oCN;DD
R--#0$MEHC##sR0NDM#N_0CF
M
NEsOHO0C0CksRs#0kRO0FvVRz4pa((X4R
H#
RRRObFlFMMC0zRvpUa4X_4U Rv
RRRRRsbF0
R5S4Sq(q,R4Rn,q,46Rcq4,4Rqdq,R4R.,q,44Rjq4,gRqRRRRRRRRRH:RM0R#8F_DoRHO;S
SqRU,qR(,qRn,qR6,qRc,qRd,qR.,qR4,qSjSSRSRRH:RM0R#8F_DoRHO;S
SA,4(RnA4,4RA6A,R4Rc,A,4dR.A4,4RA4A,R4Rj,ARgRRRRRR:RRRRHM#_08DHFoO
R;SUSA,(RA,nRA,6RA,cRA,dRA,.RA,4RA,jRASSSSR:RRRRHM#_08DHFoO
R;
RSRRdRu6u,RdRc,u,ddR.ud,dRu4u,RdRj,u,.gRUu.,.Ru(RRRRRRRRF:Rk#0R0D8_FOoHRS;
Snu.,.Ru6u,R.Rc,u,.dR.u.,.Ru4u,R.Rj,u,4gRUu4SRSRRF:Rk#0R0D8_FOoHRS;
S(u4,4Runu,R4R6,u,4cRdu4,4Ru.u,R4R4,u,4jRRugRRRRRRRR:kRF00R#8F_DoRHO;S
SuRU,uR(,uRn,uR6,uRc,uRd,uR.,uR4,uSjSSRSRRF:Rk#0R0D8_FOoHRS
S2S;
CRM8ObFlFMMC0
;
RNRR0H0sLCk0RM#$_NLDOL	_F:GRRFLFDMCN;R
RR0N0skHL0#CR$LM_D	NO_GLFRRFVvazp44UXUv_ RO:RFFlbM0CMRRH#a )z;S

#MHoNqDRQ:hRR8#0_oDFHPO_CFO0s4R5(FR8IFM0R;j2
HS#oDMNRhAQR#:R0D8_FOoH_OPC0RFs5R4(8MFI0jFR2
;
So#HMRNDu7)mR#:R0D8_FOoH_OPC0RFs5Rd68MFI0jFR2
;
S0N0skHL0\CR30HMCNsMDM_H#M0N00HNCR8\FlVRkRD0:NRDLRCDH4#R;C
Lo
HM
RRRqRQh<"=Rj&"RRSq;RR--bRk0NCRxsHFRMsRVF
M0RARRQ<hR=jR""RR&A
;
SDlk0RR:vazp44UXUv_ 
RRRRbRRFRs0lRNb5R
RRRRRRRRRR(q4RR=>q5Qh4,(2
RRRRRRRR4Rqn>R=RhqQ524n,R
RRRRRRqRR4=6R>QRqh6542R,
RRRRRRRRqR4c=q>RQ4h5c
2,RRRRRRRRRdq4RR=>q5Qh4,d2
RRRRRRRR4Rq.>R=RhqQ524.,R
RRRRRRqRR4=4R>QRqh4542R,
RRRRRRRRqR4j=q>RQ4h5j
2,RRRRRRRRRRqg=q>RQgh52R,
RRRRRRRRq=UR>QRqh25U,R
RRRRRRqRR(>R=RhqQ5,(2
RRRRRRRRnRqRR=>q5Qhn
2,RRRRRRRRRRq6=q>RQ6h52R,
RRRRRRRRq=cR>QRqh25c,R
RRRRRRqRRd>R=RhqQ5,d2
RRRRRRRR.RqRR=>q5Qh.
2,RRRRRRRRRRq4=q>RQ4h52R,
RRRRRRRRq=jR>QRqh25j,R
RRRRRRARR4=(R>QRAh(542R,
RRRRRRRRAR4n=A>RQ4h5n
2,RRRRRRRRR6A4RR=>A5Qh4,62
RRRRRRRR4RAc>R=RhAQ524c,R
RRRRRRARR4=dR>QRAhd542R,
RRRRRRRRAR4.=A>RQ4h5.
2,RRRRRRRRR4A4RR=>A5Qh4,42
RRRRRRRR4RAj>R=RhAQ524j,R
RRRRRRARRg>R=RhAQ5,g2
RRRRRRRRURARR=>A5QhU
2,RRRRRRRRRRA(=A>RQ(h52R,
RRRRRRRRA=nR>QRAh25n,R
RRRRRRARR6>R=RhAQ5,62
RRRRRRRRcRARR=>A5Qhc
2,RRRRRRRRRRAd=A>RQdh52R,
RRRRRRRRA=.R>QRAh25.,R
RRRRRRARR4>R=RhAQ5,42
RRRRRRRRjRARR=>A5Qhj
2,RRRRRRRRR6udRR=>u7)m52d6,R
RRRRRRuRRd=cR>)Rumd75c
2,RRRRRRRRRdudRR=>u7)m52dd,R
RRRRRRuRRd=.R>)Rumd75.
2,RRRRRRRRR4udRR=>u7)m52d4,R
RRRRRRuRRd=jR>)Rumd75j
2,RRRRRRRRRgu.RR=>u7)m52.g,R
RRRRRRuRR.=UR>)Rum.75U
2,RRRRRRRRR(u.RR=>u7)m52.(,R
RRRRRRuRR.=nR>)Rum.75n
2,RRRRRRRRR6u.RR=>u7)m52.6,R
RRRRRRuRR.=cR>)Rum.75c
2,RRRRRRRRRdu.RR=>u7)m52.d,R
RRRRRRuRR.=.R>)Rum.75.
2,RRRRRRRRR4u.RR=>u7)m52.4,R
RRRRRRuRR.=jR>)Rum.75j
2,RRRRRRRRRgu4RR=>u7)m524g,R
RRRRRRuRR4=UR>)Rum475U
2,RRRRRRRRR(u4RR=>u7)m524(,R
RRRRRRuRR4=nR>)Rum475n
2,RRRRRRRRR6u4RR=>u7)m5246,R
RRRRRRuRR4=cR>)Rum475c
2,RRRRRRRRRdu4RR=>u7)m524d,R
RRRRRRuRR4=.R>)Rum475.
2,RRRRRRRRR4u4RR=>u7)m5244,R
RRRRRRuRR4=jR>)Rum475j
2,RRRRRRRRRRug=u>R)5m7g
2,RRRRRRRRRRuU=u>R)5m7U
2,RRRRRRRRRRu(=u>R)5m7(
2,RRRRRRRRRRun=u>R)5m7n
2,RRRRRRRRRRu6=u>R)5m76
2,RRRRRRRRRRuc=u>R)5m7c
2,RRRRRRRRRRud=u>R)5m7d
2,RRRRRRRRRRu.=u>R)5m7.
2,RRRRRRRRRRu4=u>R)5m74
2,RRRRRRRRRRuj=u>R)5m7jS2
S
2;SRS
RRRu<u=R)5m7d8dRF0IMF2Rj;-SR-NR0	FCRMRD$dLcRH
0#
8CMRs#0k;O0
-
-R****************************************************************-RR--
-RAe.pimB5Rq,Au,R)2m7

---N-RI0H8ERR-I0H8EVRFRHqRM0bk
R--L8IH0-ERR8IH0FERVRRAHkMb0-
-R-
-Rmu)7RR-aRECVDkDRFbs80kORI5NHE80RL+RI0H8EHRI8RC2VlsFRFLDOl	RkHD0bCDHsR#3
R--
R--****************************************************************R-R-
H
DLssN$CRHC
C;kR#CHCCC38#0_oDFH4O_43ncN;DD
Ck#RCHCC03#8F_Do_HON0sHED3NDk;
#HCRC3CC#_08DHFoOM_k#MHoCN83D
D;
LDHs$NsROFsN
d;kR#CFNsOds3FOFNOlNb3D
D;
0CMHR0$ep.AmRBiHS#
oCCMsRHO5S
SN8IH0:ERR0HMCsoC;S
SL8IH0:ERR0HMCsoC;S
SM8CC_bbHCMDHCRR:HCM0o
CsS
2;SsbF0
R5SRSqR:RRRRHMR8#0_oDFHPO_CFO0sI5NHE80-84RF0IMF2Rj;S
SARRRRH:RM#RR0D8_FOoH_OPC05FsL8IH04E-RI8FMR0Fj
2;S)Sum:7RR0FkR8#0_oDFHPO_CFO0sI5NHE80+HLI8-0E4FR8IFM0R
j2S
2;S0N0skHL0\CR3MsN	:\RR0HMCsoC;N
S0H0sLCk0RL\3CMoH_C0sC:\RR0HMCsoC;N
S0H0sLCk0Rs\3CPlFCF_M_sINM:\RR0HMCsoC;M
C8.ReABpmi
;
NEsOHO0C0CksRFLDOR	#FeVR.mApBHiR#S

-q-RRGlNHllkRMVkOF0HMCRMC88CRCIEMIRNHE80RRH#MRF0CNJkDFR0RHLI8
0ESR--bbksF:#CRMVH8ER0CJR#kCNsRsNsNI$RHE80RFVslER0CMRHbRk0LRk##CHx#R
RRMVkOF0HM$RllRNG5DPNk,CNRDPNkRCL:MRH0CCosS2
S0sCkRsMHCM0oRCsHS#
LHCoM-RR-$Rll
NGSVSHRDPNkRCN>NRPDLkCRC0EMS
SS0sCkRsMPkNDC
N;SDSC#SC
SCSs0MksRDPNk;CL
CSSMH8RVS;
CRM8lN$lG
;
RORRFFlbM0CMRpvzaX4(4R(
RRRRRsbF0
R5RRRRRRRRR:qRRRHMR8#0_oDFHPO_CFO0s4R5nFR8IFM0R;j2
RRRRRRRRRRA:MRHR0R#8F_Do_HOP0COF5sR48nRF0IMF2Rj;R
RRRRRRuRRRF:Rk#0R0D8_FOoH_OPC0RFs5Rdd8MFI0jFR2S
S2R;
RMRC8FROlMbFC;M0
R
RRMOF#M0N0zRWvRRRRH:RMo0CC:sR=(R4;R

RFROMN#0MZ0R 4)m(RR:#_08DHFoOC_POs0FRR:="jjjjjjjjjjjjjjjj;j"
O
SF0M#NRM0INH8R:RRR0HMCsoCRR:=5I5NHE80+vWz-/42W2zv;R
RRMOF#M0N0HRI8RLRRH:RMo0CC:sR=5R5L8IH0WE+z4v-2z/Wv
2;RORRF0M#NRM0I8bsR:RRR0HMCsoCRR:=INH8RI+RH;8L
FSOMN#0MI0RNRssRRR:HCM0oRCs:I=RHR8N*HRI8
L;RORRF0M#NRM0IGlNR:RRR0HMCsoCRR:=lN$lGH5I8RN,ILH82
;
SR--aRECHkMb0N#Rs#CRb0DHR0HMF(R4-0LHRkOEM
	#R0RR$RbCqb0$C#RHRsNsN5$RjFR0R8IHN2-4RRFV#_08DHFoOC_POs0F5WRRz4v-RI8FMR0Fj
2;R0RR$RbCAb0$C#RHRsNsN5$RjFR0R8IHL2-4RRFV#_08DHFoOC_POs0F5WRRz4v-RI8FMR0Fj
2;
-S-RC0ERCCDl0CM#VRFRC0ERsuN0DHNRl1kRI)F#sRNC(R4-0LH#HRI8SC
0C$bR$10bHCR#sRNsRN$50jRFbRIs48-2VRFR8#0_oDFHPO_CFO0sR5RW-zv4FR8IFM0R;j2
-
S-ER0CNRbsN0HDsRbFO8k0N#RsdCRcH-L0I#RHR8C5W.*z
v2Sb0$C0Ru$RbCHN#Rs$sNRR5j0IFRN-ss4F2RV0R#8F_Do_HOP0COF.s5*vWz-84RF0IMF2Rj;S

-a-REHCRM0bk#MRHRINRHR8NNNss$VRFR-4ULRH0OMEk	S#
#MHoNqDRNNss$RRRRq:R0C$b;#
SHNoMDNRAs$sNRRRR:0RA$;bC
-
S-ER0CNRusN0HDsRuFO8k0sRNsRN$NN#RRsINssRNsRN$FdVRnH-L0EROk#M	
RRR#MHoNuDRLRkVRRRRRu:R0C$b;R
RRo#HMRNDu8sFqNss$RR:ub0$CS;

oLCHRMR-L-RD	FO_Dlk0S

-a-RECC#RF0IRFbsO#C#CO#REoNMCER0CNRPsLHNDICRHE80RbHMkR0#HFM0RGVHCI8RHE80RbHMk30#
-S-RCaER8IH0FERVER0CMRHb#k0RCNsRRHMWRzvoksFbV#RFLsRF30E
RRRsHC#xNC_:sRbF#OC#qR5,NRqs$sN2L
SCMoHR-R-RFbsO#C#R#sCH_xCNS
SqsNsNI$5H-8N4<2R=XR a55qN8IH04E-RI8FMR0FW*zv58IHN2-42W,Rz;v2
VSSFHsR8HGRMRRj0IFRH-8N.FRDFSb
SNSqs$sN5GH82=R<RWq5z5v*H+8G442-RI8FMR0FW*zvH28G;R
RRRRRCRM8DbFF;C
SMb8RsCFO#s#RCx#HC;_N
R
RR#sCH_xCLb:RsCFO#5#RAA,RNNss$R2
RCRLoRHMRR--bOsFCR##sHC#xLC_
ASSNNss$H5I84L-2=R<Ra X5LA5I0H8ER-48MFI0WFRz5v*ILH8-242,zRWv
2;RRRRRFRVs8RHGMRHR0jRFHRI8.L-RFDFbS
SSsANs5N$H28GRR<=Az5WvH*584G+2R-48MFI0WFRzHv*8;G2
CSSMD8RF;FbR-R-RGH8
RRRCRM8bOsFCR##sHC#xLC_;S

-o-RCsMCNR0C0RECu0NsHRNDu8sFkRO0NNss$$RLRDlk0DHb$oHMRC0ER-4ULRH0OMEk	F#RV-
S-ER0CMRHb#k0RR0FVlFsR-dnLRH0u0NsHRNDu8sFk#O03
RR
RRRolCMkND0:FRVsGRNRRHMjFR0R8IHNR-4oCCMsCN0
oSSCkMlD:0LRsVFRRLGHjMRRR0FILH8-o4RCsMCN
0CSlSSkGD0Rv:Rz4pa((X4
SSSSsbF0NRlb
R5SSSSS=qR>NRqs$sN52NG,S
SSASSRR=>AsNsNL$5G
2,SSSSS=uR>LRuk5V5NIG*H28L+2LG
SSSS;S2
SSSHbV_H4bN:VRHRC5MCb8_HDbCHRMC=2R4RMoCC0sNCS
SSkSLVHbb:FRVsRRHHjMRRR0F.z*WvR-4oCCMsCN0
SSSS0SN0LsHkR0C\N3sMR	\FsVRCRo#:NRDLRCDH4#R;S
SSNSS0H0sLCk0RL\3CMoH_C0sCF\RVCRso:#RRLDNCHDR#;R4
SSSS0SN0LsHkR0C\C3slCFP__MFIMNs\VRFRosC#RR:DCNLD#RHR
4;SSSSLHCoMSR
SSSSs#Co:bRRHLbCkSV
SSSSSsbF0NRlbS5
SSSSSRSQ=u>RL5kV5*NGILH82G+L225H,S
SSSSSS=mR>sRuFs8qs5N$5*NGILH82G+L225H
SSSS2SS;S
SSMSC8CRoMNCs0LCRkbVbHS;
SMSC8CRoMNCs0HCRVH_bb;N4
SSSHbV_HjbN:VRHRC5MCb8_HDbCHRMC=2RjRMoCC0sNCS
SSsSuFs8qs5N$5*NGILH82G+L2=R<RkuLVN55GH*I8+L2L;G2
SSSCRM8oCCMsCN0R_HVbNHbjS;
S8CMRMoCC0sNCCRoMDlk0
L;S8CMRMoCC0sNCCRoMDlk0
N;
-S-R	aNCER0CNRusN0HDsRuFO8k0sRNsRN$NRM8LDkH8ER0C8RN8RCs0CsC3qRRRMskMoHMRl#k
-S-RRH#H0MHNxDHCR8,0MECREF0CssRFRI#F0VREbCRNHs0NbDRskF8ON0RsNCR888C3-
S-FRwsGRCNDlbCH,RVRRqH6#RUH-L0I#RHR8CNRM8A#RHR-.cL#H0R8IHC0,RERCMqHRV0H#RM
RcSR--4L(-HO0RE	kM#MRN8RRAV#H0RRHM.(R4-0LHRkOEM3	#RERaCsRNsRN$IDHDROHMDCk8R.c*=-
S-RRUl0kDHHbDCRs#VlFsHRMoUnRd-0LHRsuN0DHNRFus80kO#R3RaRECVDkDRFbs80kORDIHDCRLR-
S-+Rc.R=n4L(-HO0RE	kM#HRI8RC3RswFRH0E#GRCNDlbCER0CkR)Ml1kRRH#H0MHHHNDxRC80
F:SR--RjRR'R#,RRRRR'Rj#R,RRRRRR5uu42,4ERH,u4u5,D42Fu,Ru,5jjH2E,uRu5jj,2
DFSR--aMECREF0CssRFRI#NRsCVlFsCL8RN8#CRRFM0RECI0H8EVRFRHqRM(R4-0LHRkOEMR	#N
M8SR--0RECI0H8EVRFRHARM(R4-0LHRkOEM3	#RFRwsER0CGRCNDlbCS:
-a-RE'CRqD'RFRFb504RF2Rd
-S-RRRRj,'#RRRRRuRRu,5.4H2E,uRu54.,2,DFR5uu42,jERH,u4u5,Dj2Fj,R'S#
-R-RRuRu54d,2,EHR5uud2,4DRF,u.u5,Ej2Hu,Ru,5.jF2D,'Rj#R,RRRRRR#j'
-S-RRRRj,'#RRRRRuRRu,5djH2E,uRu5jd,2,DFR#j',RRRRRRRj,'#RRRRRjRR'S#
-a-RE'CRAD'RFRFb504RF2R4
-S-RRRRj,'#RRRRRjRR'R#,RRRRR'Rj#R,RRRRRR5uuj2,4ERH,uju5,D42Fj,R'
#
RNRR8s8bFR8:bOsFCR##5Fus8sqsN
$2SNSPsLHND)CRkkM1lRRRR#:R0D8_FOoH_OPC05FsI8bs*vWz-84RF0IMF2RjRR:=5EF0CRs#='>Rj;'2
RRRRPRRNNsHLRDC1)klFCIeORR:#_08DHFoOC_POs0F5sIb8z*WvR-48MFI0jFR2R;
RRRRRsPNHDNLCkR1lI)FRRRR:0R1$;bC
RRRRPRRNNsHLRDCNGH8RRRRRRR:HCM0o;Cs
RRRRPRRNNsHLRDCLGH8RRRRRRR:HCM0o;Cs
RRRRPRRNNsHLRDC[RRRRRRRRRR:HCM0o;Cs
RRRRPRRNNsHLRDC	RRRRRRRRRR:HCM0o;Cs
CSLoRHMRR--bOsFCR##Nb88s
F8S-S-RHQM0DHNHRxC0RECsMkMHRMo#Rkl5M)k12kl
RRRRVRRFNsRGMRHR0jRFlRIN4G-RFDFbS
SS8LHG=R:R;NG
SSS[RRRRR:=.G*N;S
SSR	RR=R:R+[RR
4;SHSSVGRNRI>RH-8N4sRFR8LHGRR>ILH8-04RE
CMSSSSH[VRRI<RbRs80MECRSRSRR--xFCsR0CGC
M8SSSSSl1k)5FI[:2R= RZ)(m4;S
SSMSC8VRH;S
SSVSHR<	RRsIb8ER0CRMRS-SR-CRxsCFRGM0C8S
SS1SSkFl)I25	RR:=Zm )4
(;SSSSCRM8H
V;SCSSD
#CSSSS1)klF[I52=R:RFus8sqsNN$5GH*I8LL+H28G5WRRz4v-RI8FMR0FR2Rj;R
RRRRRRRRRRVRHR<	RRsIb8ER0CSM
SSSS1)klF	I52=R:RFus8sqsNN$5GH*I8LL+H28G5W.*z4v-RI8FMR0FW2zv;S
SSMSC8VRH;S
SS8CMR;HV
SSS-O-RFCMPs00RENCRs$sNRRFVOMEk	H#RMR0FNNMRs$sNRRFVL#H0
SSSVRFsHRLGHjMRRR0FI8bs-D4RF
FbSSSSVRFsDHGRMRRj0WFRz4v-RFDFbS
SS)SSkkM1lL5HGz*WvG+D2=R:Rl1k)5FIH2LG52DG;S
SSMSC8FRDFRb;RR--DSG
SMSC8FRDFRb;RR--H
LGSMSC8FRDFRb;RR--NSG
SR--pbFFRRFM0RECqMRH8
CGSFSVs8RHGMRHR04RFHRI84N-RFDFbR
RRRRRRVRRFNsRGMRHR0jRFlRIN4G-RFDFbS
SSHSL8:GR=GRNRH-R8
G;SSSS[RRRRR:=N+GRR8LHGS;
S	SSRRRR:[=RR4+R;S
SSVSHRRNG>HRI84N-RRFsLGH8RI>RH-8L4ER0CRM
RRRRRRRRRRRRRVRHR<[RRsIb8ER0CRMRS-SR-CRxsCFRGM0C8S
SSSSS1)klF[I52=R:R)Z m;4(
SSSSMSC8VRH;S
SSHSSVRR	<bRIs08RERCMRRSS-x-RCRsFCCG0MS8
SSSSSl1k)5FI	:2R= RZ)(m4;S
SSCSSMH8RVS;
SCSSDV#HR8LHGRR<jER0CSM
SSSSH[VRRj<RRC0EMS
SSSSS[=R:R+[RRI.*l;NG
RRRRRRRRRRRRRRRCRM8H
V;RRRRRRRRRRRRRHRRVRR	<RRj0MEC
SSSS	SSRR:=	RR+.l*IN
G;SSSSS8CMR;HV
SSSSVSHR<[RRRNG0MEC
SSSS1SSkFl)I25[RR:=Zm )4
(;SSSSS#CDH[VRRI<RbRs80MEC
SSSS1SSkFl)I25[RR:=Zm )4R(;RR--xFCsR0CGC
M8SSSSS8CMR;HV
SSSS-S-REF0CHsI#RC,0RECHCM8G#RHR0MFRRHM0REC1)klFRI,8MFRFH0EMSo
SSSSH	VRRR<=N0GRE
CMSSSSSkS1lI)F5R	2:Z=R 4)m(R;
RRRRRRRRRRRRRDRC#RHV	RR<I8bsRC0EMS
SSSSS1)klF	I52=R:R)Z m;4(R-R-RsxCFGRC08CM
SSSS-S-REF0CHsI#RC,0RECHCM8G#RHR0MFRRHM0REC1)klFRI,8MFRFH0EMSo
SSSSCRM8H
V;SSSSCCD#
SSSSkS1lI)F5R[2:u=RsqF8s$sN5*NGILH8+8LHGR25RvWz-84RF0IMFRRRj
2;RRRRRRRRRRRRRHRRVRR	<bRIs08RE
CMSSSSSkS1lI)F5R	2:u=RsqF8s$sN5*NGILH8+8LHG.25*vWz-84RF0IMFzRWv
2;SSSSS8CMR;HV
SSSS8CMR;HV
SSSCRM8DbFF;-RR-GRN
SSS-O-RFCMPs00RENCRs$sNRRFVOMEk	H#RMR0FNNMRs$sNRRFVL#H0
RRRRRRRRFRVsLRHGMRHR0jRFbRIs48-RFDFbS
SSFSVsGRDRRHMjFR0RvWz-D4RF
FbSSSSSl1k)eFICHO5LWG*zDv+G:2R=kR1lI)F5GHL2G5D2S;
SCSSMD8RF;FbR-R-R
DGSCSSMD8RF;FbR-R-RGHL
SSS-q-R808REsCRF[IRkR#0ONsC0RC800FREsCRkHMMM#oRkRl
RRRRRRRR)1kMk:lR=kR)Ml1kR1+RkFl)IOeC;S
SCRM8DbFF;-RR-8RHGS
S-p-RFRFbF0MREACRR8HMCSG
SsVFRGHxRRHM4FR0R8IHLR-4DbFF
RRRRRRRRFRVsGRLRRHMjFR0RNIlGR-4DbFF
SSSS8NHG=R:RRLG-xRHGS;
S[SSRRRR:N=RHR8G+GRL;S
SSRS	R:RR=RR[+;R4
SSSSRHVL>GRR8IHLR-4FNsRHR8G>HRI84N-RC0EMR
RRRRRRRRRRRRRRRHV[RR<I8bsRC0EMSRRS-R-RsxCFGRC08CM
SSSS1SSkFl)I25[RR:=Zm )4
(;SSSSS8CMR;HV
SSSSVSHR<	RRsIb8ER0CRMRS-SR-CRxsCFRGM0C8S
SSSSS1)klF	I52=R:R)Z m;4(
SSSSMSC8VRH;S
SSDSC#RHVNGH8Rj<RRC0EMS
SSHSSVRR[<RRj0MECRSRSS-R-R[N8kR#00RECHOM8HRC#lkF8DIFRl
NGSSSSSRS[:[=RR.+R*NIlGS;
SSSSCRM8H
V;SSSSSRHV	RR<jER0CSM
SSSSS:	R=RR	+*R.IGlN;S
SSCSSMH8RVS;
SSSSH[VRRL<RGER0CSM
SSSSSl1k)5FI[:2R= RZ)(m4;R
RRRRRRRRRRRRRR#CDH[VRRI<RbRs80MECRRRRRR--xFCsR0CGC
M8SSSSSkS1lI)F5R[2:Z=R 4)m(S;
SSSSCRM8H
V;SSSSSRHV	=R<RRLG0MEC
SSSS1SSkFl)I25	RR:=Zm )4
(;RRRRRRRRRRRRRCRRDV#HR<	RRsIb8ER0CRMRR-RR-CRxsCFRGM0C8S
SSSSS1)klF	I52=R:R)Z m;4(
SSSSMSC8VRH;S
SSDSC#SC
SSSS1)klF[I52=R:RFus8sqsNN$5H*8GILH8+2LG5WRRz4v-RI8FMR0FR2Rj;R
RRRRRRRRRRRRRRRHV	RR<I8bsRC0EMS
SSSSS1)klF	I52=R:RFus8sqsNN$5H*8GILH8+2LG5W.*z4v-RI8FMR0FW2zv;S
SSCSSMH8RVS;
SCSSMH8RVS;
SMSC8FRDFRb;RR--LSG
S-S-RMOFP0CsRC0ERsNsNF$RVEROk#M	R0HMFMRNRsNsNF$RVHRL0R#
RRRRRRRRVRFsHRNGHjMRRR0FI8bs-D4RF
FbSSSSVRFsDHGRMRRj0WFRz4v-RFDFbS
SS1SSkFl)IOeC5GHN*vWz+2DGRR:=1)klFHI5N5G2D;G2
SSSS8CMRFDFbR;R-D-RGS
SS8CMRFDFbR;R-H-RNSG
S-S-R8q8RC0ERIsFR#[k0sROCCN08FR0RC0ERMskMoHMRl#k
RRRRRRRRkR)Ml1kRR:=)1kMk+lRRl1k)eFIC
O;SMSC8FRDFRb;RR--H
xGS-S-RCaER0FkbRk0b8sFkRO0H8#RCHsPCV8RsRFl0RECsMkMHRMo#
klRRRRR)Rum<7R=kR)Ml1k5HNI8+0EL8IH04E-RI8FMR0Fj
2;S8CMRFbsO#C#R8N8b8sF;C

ML8RD	FO#
;
-*-R*************************************************************R**R
---
-R- -RM00H$CR7OsDNNF0HMFRVsMRk#MHoCl8RkHD0bCDHs-
-R-
-RHaE##RHRC0ERHlNMMRC0$H0RsVFRC0ER#kMHCoM8kRlDb0HDsHC3aRRE0CRINFRsHOE00COk#sC
R--8HCVMRC8LFCDI#RkCER0CMRC0HH0CN#RLCFP,MRN8kRl#L0RCNRD#H0RMER0HV#RH3DCRERaC-
-RF0IRONsECH0Os0kCN#Rs0CREDCRFOoHRsPC#MHFR8NMRC0ERFLDOP	RCHs#F
M3-
-R-*-R*************************************************************R**R
--
LDHs$NsRCHCCk;
#HCRC3CC#_08DHFoO4_4nNc3D
D;kR#CHCCC38#0_oDFHNO_sEH03DND;#
kCCRHC#C30D8_FOoH_#kMHCoM8D3ND
;
DsHLNRs$#b$MD$HV;#
kC$R#MHbDVN$30H0sLCk0#D3ND
;
DsHLNRs$FNsOdk;
#FCRsdON3OFsNlOFbD3ND
;
CHM00v$RzRpaHR#
RoRRCsMCH
O5RRRRRIRRHE80RRR:HCM0oRCs:.=RcR;
RRRRRIRNHE80RH:RMo0CC:sR=.R4;R
RRRRRRHLI8R0E:MRH0CCos=R:R
4.S2SR;R
RRFRbs
05SqSRRRRR:MRHR8#0_oDFHPO_CFO0sI5NHE80RR-48MFI0jFR2S;
SRRAR:RRRRHM#_08DHFoOC_POs0F5HLI8R0E-84RF0IMF2Rj;S
SRmu)7RR:FRk0#_08DHFoOC_POs0F58IH0-ER4FR8IFM0R
j2RRRRR2RR;R
RR0N0skHL0\CR3MsN	:\RR0HMCsoC;R
RR0N0skHL0\CR38lFk\DCR#:R0MsHoR;
R0RN0LsHkR0C\F3b8\ClRH:RMo0CC
s;RNRR0H0sLCk0Rb\3Fl8CL\k#R#:R0MsHoR;
R0RN0LsHkR0C\M3C8s_0CRC\:MRH0CCosR;
R0RN0LsHkR0C\C3Lo_HM0CsC\RR:HCM0o;Cs
RRRNs00H0LkC3R\sFClPMC_FN_IsRM\:MRH0CCosC;
Mv8Rz;pa
-
-R****************************************************************-RR--
-R-
-RoDFHNORsHOE00COk#sCRsVFROmsN
R6-
-R-*-R*************************************************************R**R
--
ONsECH0Os0kCFRDoRHOFvVRzRpaH
#
-V-RHRM80RECDoNsCIsRHE80RH5I8N0ERRFsI0H8E
L2
RRRVOkM0MHFRb#k58IH0,ENR8IH0REL:MRH0CCoss2RCs0kMMRH0CCos#RH
RRRLHCoMR
RRRRRH5VRI0H8E>NRR8IH02ELRC0EMR
RRRRRRsRRCs0kMHRI8N0E;R
RRRRRCCD#
RRRRRRRRCRs0MksR8IH0;EL
RRRRCRRMH8RVR;
RMRC8kR#b
;
-V-RHRM80REC#DlNDRCsI0H8EIR5HE80NsRFR8IH02EL
R
RRMVkOF0HMMRHVH5I8N0E,HRI8L0ERH:RMo0CCRs2skC0sHMRMo0CCHsR#R
RRoLCHRM
RRRRRRHV58IH0REN<HRI8L0E2ER0CRM
RRRRRRRRskC0sIMRHE80NR;
RRRRR#CDCR
RRRRRRsRRCs0kMHRI8L0E;R
RRRRRCRM8H
V;RCRRMH8RM
V;
R--0RECVDFDFMIHoMRC#Cks#ER0NI0RHE80A#RHRINDNR$#oNsC0RCs0MENRRFsCNJkDFR0R8IH0
Eq-k-R#oHMRk'#bN'RM'8RH'MV3R

RFROMN#0MI0RHE80qRR:HCM0oRCs:H=RMNV5I0H8EL,RI0H8E
2;RORRF0M#NRM0I0H8E:ARR0HMCsoCRR:=#5kbN8IH0RE,L8IH0;E2
-
-RC0ERlOFbCFMMw0RH0s#u8sFk#O0RC5#CLRNF2PC
R
RRlOFbCFMMw0RH0s#u8sFk#O0
RRRoCCMs5HO
RRRRIRRHE80qRR:HCM0o;Cs
RRRRIRRHE80ARR:HCM0o
CsR2RR;R
RRsbF0
R5RRRRRRRqRH:RM#RR0D8_FOoH_OPC05FsN8IH04E-RI8FMR0Fj
2;RRRRRRRARH:RM#RR0D8_FOoH_OPC05FsL8IH04E-RI8FMR0Fj
2;RRRRRARqRF:Rk#0R0D8_FOoH_OPC05FsL8IH0NE*I0H8ER-48MFI0jFR2R
RRRRR-A-RRq*R
RRR2R;
RMRC8FROlMbFC;M0
-
-RC0ERlOFbCFMMN0R8s8CaCsCRC5#CLRNF2PC
R
RRlOFbCFMMN0R8s8CaCsC
RRRoCCMs5HO
RRRRIRRHE80qRR:HCM0o;Cs
RRRRIRRHE80ARR:HCM0o
CsR2RR;R
RRsbF0
R5RRRRRARqRRRRRRR:H#MR0D8_FOoH_OPC05FsL8IH0NE*I0H8ER-48MFI0jFR2R;
RRRRRFbs80kORF:Rk#0R0D8_FOoH_OPC05FsL8IH0NE+I0H8ER-48MFI0jFR2R
RRRRR-A-RRq*R
RRR2R;
RMRC8FROlMbFC;M0
R
RRo#HMRNDNk_NG:RRR8#0_oDFHPO_CFO0sH5I8q0E-84RF0IMF2Rj;R
RRo#HMRNDLk_NG:RRR8#0_oDFHPO_CFO0sH5I8A0E-84RF0IMF2Rj;R
RRo#HMRNDNRLRR:RRR8#0_oDFHPO_CFO0sI5NHE80*HLI8-0E4FR8IFM0R;j2
RRR#MHoNsDRCD#k0RR:#_08DHFoOC_POs0F5HNI8+0EL8IH04E-RI8FMR0Fj
2;
R--0RECV#Hs0sRNO0EHCkO0sVCRF0sRElCRkHD0bRD$-MRNRsNsNL$RN8#CRDlk0DHbH
Cs
oLCH
MRR-RR-IR1NqbRR8NMRHARVCRMO#C#N3s$RR
RRqHVDoNsC:sARRHV5HNI8R0E>IRLHE802CRoMNCs0RC
RRRRRsVFDbFF.V:RFHsRRRHMjFR0RHLI8-0E4CRoMNCs0RC
RRRRRRRRNs00H0LkC3R\s	NM\VRFRosC#:qRRLDNCHDR#;Rj
SSSNs00H0LkC3R\sFClPMC_FN_IsRM\FsVRCqo#RD:RNDLCRRH#4R;
RRRRRRRRNs00H0LkC3R\s	NM\VRFRosC#:ARRLDNCHDR#;Rj
SSSNs00H0LkC3R\sFClPMC_FN_IsRM\FsVRCAo#RD:RNDLCRRH#4R;
RRRRRoLCHRM
RRRRRRRRs#CoqR:RbCHbL
kVRRRRRRRRRsbF0NRlbR5
RRRRRRRRRQRRRR=>A25H,R
RRRRRRRRRRRRm=N>R_GNk5
H2RRRRRRRRR
2;RRRRRRRRRosC#RA:RbbHCVLk
RRRRRRRRFRbsl0RN
b5RRRRRRRRRRRRQ>R=RHq52R,
RRRRRRRRRmRRRR=>Lk_NG25H
RRRRRRRR;R2
RRRRCRRMo8RCsMCNR0CVDFsF.Fb;R

RRRRRsVFDbFF4V:RFHsRRRHML8IH00ERFIRNHE80-o4RCsMCN
0CRRRRRRRRR0N0skHL0\CR3MsN	F\RVCRsoR#A:NRDLRCDHj#R;S
SS0N0skHL0\CR3lsCF_PCMIF_N\sMRRFVs#CoARR:DCNLD#RHR
4;RRRRRCRLo
HMRRRRRRRRRosC#RA:RbbHCVLk
RRRRRRRRFRbsl0RN
b5RRRRRRRRRRRRQ>R=RHq52R,
RRRRRRRRRmRRRR=>Lk_NG25H
RRRRRRRR;R2
RRRRCRRMo8RCsMCNR0CVDFsF4Fb;R
RR8CMRMoCC0sNCVRHqsDNoACs;R

R-R-RCz#R&qRRIARHF0Ek#0RIbNbH3Mo
RRRH#VqlDNDC:sARRHV5HNI8R0E<L=RI0H8Eo2RCsMCN
0CRRRRRFRVsFDFbRN:VRFsHMRHR0jRFIRNHE80-o4RCsMCN
0CRRRRRRRRR0N0skHL0\CR3MsN	F\RVCRsoR#B:NRDLRCDHj#R;S
SS0N0skHL0\CR3lsCF_PCMIF_N\sMRRFVs#CoBRR:DCNLD#RHR
4;RRRRRRRRR0N0skHL0\CR3MsN	F\RVCRsoR#1:NRDLRCDHj#R;S
SS0N0skHL0\CR3lsCF_PCMIF_N\sMRRFVs#Co1RR:DCNLD#RHR
4;RRRRRCRLo
HMRRRRRRRRRosC#RB:RbbHCVLk
RRRRRRRRFRbsl0RN
b5RRRRRRRRRRRRQ>R=RHq52R,
RRRRRRRRRmRRRR=>Nk_NG25H
RRRRRRRR;R2
RRRRRRRRCRso:#1RHRbbkCLVR
RRRRRRbRRFRs0l5Nb
RRRRRRRRRRRR=QR>5RAH
2,RRRRRRRRRRRRm>R=RNL_kHG52R
RRRRRR2RR;R
RRRRRCRM8oCCMsCN0RsVFDbFFN
;
RRRRRFRVsFDFbRL:VRFsHMRHRHNI8R0E0LFRI0H8ER-4oCCMsCN0
RRRRRRRR0RN0LsHkR0C\N3sMR	\FsVRC7o#RD:RNDLCRRH#jS;
S0SN0LsHkR0C\C3slCFP__MFIMNs\VRFRosC#:7RRLDNCHDR#;R4
RRRRLRRCMoH
RRRRRRRRCRso:#7RHRbbkCLVR
RRRRRRbRRFRs0l5Nb
RRRRRRRRRRRR=QR>5RAH
2,RRRRRRRRRRRRm>R=RNL_kHG52R
RRRRRR2RR;R
RRRRRCRM8oCCMsCN0RsVFDbFFLR;
RMRC8CRoMNCs0HCRVlq#NCDDs
A;
RRRw#Hs0C10bw:RH0s#u8sFk#O0
RRRRoRRCsMCHlORN5bR
RRRRRRRRHRI8q0ERR=>I0H8E
q,RRRRRRRRR8IH0REA=I>RHE80AR
RRRRR2R
RRRRRb0FsRblNRR5
RRRRRRRRq>R=RNN_k
G,RRRRRRRRR=AR>_RLN,kG
RRRRRRRRARqRR=>NRL
RRRRR
2;
RRRqC88sCasC:.RR8N8CssaCRC
RRRRRMoCCOsHRblNRR5
RRRRRRRRI0H8E=qR>HRI8q0E,R
RRRRRRIRRHE80A>R=R8IH0
EARRRRR
R2RRRRRFRbsl0RN5bR
RRRRRRRRARqRR=>N
L,RRRRRRRRRFbs80kORR=>skC#DR0
RRRRR
2;
RRRRmu)7=R<R#sCk5D0I0H8ER-48MFI0jFR2C;
MD8RFOoH;-

-*R**************************************************************R*R---
--R
-DRLF_O	l0kDRONsECH0Os0kCV#RFmsRsRON6-
-R-
-R****************************************************************-RR-N

sHOE00COkRsCLODF	k_lDF0RVzRvpHaR#S

-b-RkFsb#RC:skC0sRM#0RECMRCII0H8ENRL#RC8FCMRG#OC#HRL0L#RCoHMRCbs#0CM
RRRVOkM0MHFR#bN#8WH05ER
RRRRORRF0M#NRM0lIF8HE80RH:RMo0CC
s;RRRRRFROMN#0MF0RDH8W8R0E:MRH0CCosS2
S0sCkRsMHCM0oRCsHS#
LHCoM-RR-NRb#H#W8
0ERRRRRVRHR8lFI0H8ERR>.ER0CRMR-l-RFR#00CN	RH0E#sRLNEMO
SSSskC0sFMRDH8W8;0E
CSSDV#HR8lFI0H8ERR=.ER0CSM
SCSs0MksR8FDW0H8E;-.
CSSDV#HR8lFI0H8ERR=4ER0CSM
SCSs0MksR8FDW0H8E;-4
CSSDV#HR8lFI0H8ERR=jER0CSM
SCSs0MksR8FDW0H8ES;
S#CDCSRRSSSSRR--0#EHRRH##CkbskVDF
k#SsSSCs0kMDRF88WH0
E;SMSC8VRH;C
SMb8RNW##HE80;S

-b-RkFsb#RC:skC0sRM#4VRHRCMC8FR0RR8FbCHbDHHMMSo
VOkM0MHFRNNMDC$#_bHMkI0_HE805HNI8L,RIRH8:MRH0CCoss2RCs0kMMRH0CCos#RH
CSLo
HMSVSHRN55IRH8>(R42MRN8LR5IRH8>(R4202RE
CMSsSSCs0kM;R4
RRRRCRRMH8RVS;
S0sCkRsMjS;
CRM8NDMN$_#CHkMb0H_I8;0E
R
RRR--V8HMRC0ERN#lDsDCR8IH05ERI0H8EsRFRHNI820E
RRRVOkM0MHFRVHM58IH0RE,N8IH0:ERR0HMCsoC2CRs0MksR0HMCsoCR
H#RLRRCMoH
RRRRHRRVIR5HE80RN<RI0H8E02RE
CMRRRRRRRRR0sCkRsMI0H8ER;
RRRRR#CDCR
RRRRRRsRRCs0kMIRNHE80;R
RRRRRCRM8H
V;RCRRMH8RM
V;
RRRO#FM00NMRvWzRRRR:MRH0CCos=R:R;4(
SSSSRSS
RRRO#FM00NMRHNI8RCR:MRH0CCos=R:RVHM58IH0RE,N8IH0;E2
FSOMN#0ML0RICH8RRR:HCM0oRCs:H=RMIV5HE80,IRLHE802S;
SSSSSRR
RFROMN#0MN0RlRF8RRR:HCM0oRCs:N=RICH8-5555HNI8WC+z4v-2z/Wv42-2z*Wv
2;RORRF0M#NRM0L8lFR:RRR0HMCsoCRR:=L8IHC5-55I5LH+8CW-zv4W2/z-v24W2*z;v2
SSSSRSS
RRRO#FM00NMRHNI8RRS:MRH0CCos=R:R#bN#8WH0NE5l,F8RHNI8;C2
RRRO#FM00NMRHLI8RRS:MRH0CCos=R:R#bN#8WH0LE5l,F8RHLI8;C2
R
RRMOF#M0N0CRMCb8_HDbCHRMC:MRH0CCos=R:RNNMDC$#_bHMkI0_HE805HNI8,0ERHLI820E;S
SSRSSR
SRSo#HMRNDCR4RRSRRR#:R0D8_FOoH_OPC05Fs4FR8IFM0R;j2
HS#oDMNRRC.RRRRSRR:#_08DHFoOC_POs0F584RF0IMF2Rj;S
SSRSSR
SRR#RRHNoMD0RqsRHlR:RRR8#0_oDFHPO_CFO0sI5NH-8C4FR8IFM0R;j2
RRR#MHoNADR0lsHRRRR:0R#8F_Do_HOP0COFLs5ICH8-84RF0IMF2Rj;R

RHR#oDMNRsqbHRlCRRR:#_08DHFoOC_POs0F5HNI8R-48MFI0jFR2R;
RHR#oDMNRsAbHRlCRRR:#_08DHFoOC_POs0F5HLI8R-48MFI0jFR2R;
RHR#oDMNRF1EsR0uRRR:#_08DHFoOC_POs0F5HNI8I+LH48-RI8FMR0Fj
2;SSSSS
SRR#RRHNoMDCR)#0kD4:RRR8#0_oDFHPO_CFO0sI5NH+8CL8IHCR-48MFI0jFR2R;
RHR#oDMNR#)CkGD0RRR:#_08DHFoOC_POs0F5HNI8LC+ICH8-84RF0IMF2Rj;R
RRo#HMRND)kC#DR0NR#:R0D8_FOoH_OPC05FsN8IHCI+LH-8C4FR8IFM0R;j2
RRR#MHoN)DRCD#k0RLR:0R#8F_Do_HOP0COFNs5ICH8+HLI84C-RI8FMR0Fj
2;R#RRHNoMDCR)#0kDC:RRR8#0_oDFHPO_CFO0sI5NH+8CL8IHCR-48MFI0jFR2=R:R05FE#CsRR=>'2j';R

RHR#oDMNRFus8N4_kRG,u8sF4C_s#RRR:0R#8F_Do_HOP0COFNs5ICH8+HLI84C-RI8FMR0Fj
2;R#RRHNoMDsRuFR84R:RRR8#0_oDFHPO_CFO0sI5NH+8CL8IHCR-48MFI0jFR2R;
RHR#oDMNRFus8R.RRRR:#_08DHFoOC_POs0F58IH04E-RI8FMR0Fj
2;
FSOlMbFCRM0ep.Am
BiSCSoMHCsO
R5SNSSI0H8ERR:HCM0oRCs:N=RI;H8
SSSL8IH0:ERR0HMCsoCRR:=L8IH;S
SSCMC8H_bbHCDM:CRR0HMCsoCRR:=M8CC_bbHCMDHC
2;SFSbs50R
SSSqRRRRH:RM#RR0D8_FOoH_OPC05FsN8IH-84RF0IMF2Rj;S
SSRARRRR:HRMR#_08DHFoOC_POs0F5HLI8R-48MFI0jFR2S;
S)Sum:7RR0FkR8#0_oDFHPO_CFO0sI5NHL8+I-H84FR8IFM0R2j2;C
SMO8RFFlbM0CM;L

CMoHR-R-RFLDOl	_k
D0
-S-RsbkbCF#:NR0	OCRNRsCF0VRE4CRR8NMRL.-HO0RN##C
-S-Rb0$CRRR:FROlMLHNF0HM
NDSR--HkMb0:#RRRq,A-
S-kRF00bk#u:R)
m7SR--0lsHRC0ERbHMkR0#0LFRCFRMR8IHC0sRERNM0RECFbk0kS0
HoV_CRM:H5VRM8CC_bbHCMDHCRR=4o2RCsMCN
0CSsS0H0lHqV:RFHsRRRHMjFR0RHNI84C-RMoCC0sNCS
SS0N0skHL0\CR3MsN	F\RVCRsoR#q:NRDLRCDHj#R;S
SS0N0skHL0\CR38bFCRl\FsVRCqo#RD:RNDLCRRH#HS;
S0SN0LsHkR0C\F3b8LClkR#\FsVRCqo#RD:RNDLCRRH#";q"
SSSNs00H0LkC3R\lkF8DRC\FsVRCqo#RD:RNDLCRRH#"pvza
";SNSS0H0sLCk0Rs\3CPlFCF_M_sINMF\RVCRsoR#q:NRDLRCDH4#R;S
SLHCoMS
SSosC#Rq:RbbHCVLk
SSSSsbF0NRlbS5
SSSSQ>R=RHq52S,
SSSSm>R=Rsq0HHl52S
SS;S2
CSSMo8RCsMCNR0C0lsHH;0q
R
RSsS0H0lHAV:RFHsRRRHMjFR0RHLI84C-RMoCC0sNCS
SS0N0skHL0\CR3MsN	F\RVCRsoR#A:NRDLRCDHj#R;S
SS0N0skHL0\CR38bFCRl\FsVRCAo#RD:RNDLCRRH#HS;
S0SN0LsHkR0C\F3b8LClkR#\FsVRCAo#RD:RNDLCRRH#";A"
SSSNs00H0LkC3R\lkF8DRC\FsVRCAo#RD:RNDLCRRH#"pvza
";SNSS0H0sLCk0Rs\3CPlFCF_M_sINMF\RVCRsoR#A:NRDLRCDH4#R;S
SLHCoMS
SSosC#RA:RbbHCVLk
SSSSsbF0NRlbS5
SSSSQ>R=RHA52S,
SSSSm>R=RsA0HHl52S
SS;S2
CSSMo8RCsMCNR0C0lsHH;0A
MSC8CRoMNCs0HCRVC_oM
;
S_HVojCM:VRHRC5MCb8_HDbCHRMC=2RjRMoCC0sNCS
SqH0sl=R<RNq5ICH8-84RF0IMF2Rj;S
SAH0sl=R<RLA5ICH8-84RF0IMF2Rj;C
SMo8RCsMCNR0CHoV_C;Mj
-
S-CRslCFPRC0ER0CGsLNRHR0#N00REpCR1CARMR8
RsRbkHMC0b:RsCFO#5#RqH0slA,R0lsH2L
SCMoHR-R-RFbsO#C#RkbsM0CH
HSSVlRNF=8RR04RE
CMSCSS4=R<R''jRq&R0lsH5;j2
SSSqHbsl<CR=0Rqs5HlN8IHCR-48MFI04FR2S;
S#CDHNVRlRF8=RR.0MEC
RRRRRRRR4RCRR<=qH0slR548MFI0jFR2S;
SbSqsCHlRR<=qH0slI5NH-8C4FR8IFM0R;.2
RRRRCRRD
#CSCSS4=R<R''jR'&Rj
';SqSSblsHC=R<Rsq0H
l;SMSC8VRH;S

SRHVL8lFR4=RRC0EMS
SSRC.<'=Rj&'RRsA0Hjl52S;
SbSAsCHlRR<=AH0slI5LH-8C4FR8IFM0R;42
CSSDV#HRFLl8RR=.ER0CRM
RRRRRRRRC<.R=0RAs5Hl4FR8IFM0R;j2
SSSAHbsl<CR=0RAs5HlL8IHCR-48MFI0.FR2R;
RRRRR#CDCS
SSRC.<'=Rj&'RR''j;S
SSsAbHRlC<A=R0lsH;S
SCRM8H
V;S8CMRFbsO#C#RkbsM0CH;S

-v-RkHD0bRD$L0$RECCRGN0sR0LH#VRHRRICECNPRCFMRRFs0RIFCsG0NHRL0F#RV
RqS_HVNR4:H5VRN8lFR4=R2CRoMNCs0SC
S_HVNj4L:VRHRl5LF<8R=RRjFLsRlRF8>2R.RMoCC0sNCS
SS#)CkND0RR<=Bemh_71a_tpmQeB_ mBa),5jRHNI8LC+ICH82ERIC5MRCj452RR='2j'RS
SSSSSRDRC# CRXAa5blsHCN,RICH8+HLI8;C2
RRRRCRRMo8RCsMCNR0CHNV_4;Lj
HSSV4_NLR4:H5VRL8lFR4=R2CRoMNCs0SC
SCS)#0kDN=R<RhBmea_17m_pt_QBea Bmj)5,IRNH+8CL8IHCI2RERCM55C4j=2RR''j2SR
SSSSSCRRDR#C 5XaAHbsl&CRR''j,IRNH+8CL8IHC
2;RRRRRMRC8CRoMNCs0HCRV4_NL
4;SVSH_LN4.H:RVLR5lRF8=2R.RMoCC0sNCS
SS#)CkND0RR<=Bemh_71a_tpmQeB_ mBa),5jRHNI8LC+ICH82ERIC5MRCj452RR='2j'RS
SSSSSRDRC# CRXAa5blsHCRR&'Rj'&jR''N,RICH8+HLI8;C2
RRRRCRRMo8RCsMCNR0CHNV_4;L.
MSC8CRoMNCs0HCRV4_N;H
SV._N:VRHRl5NF=8RRR.2oCCMsCN0
RRRR#RRHNoMDFRM1VEH0#,RE0HVCR8,NC888RR:#_08DHFoOC_POs0F5HNI8LC+ICH8-84RF0IMF2Rj;L
SCMoH
HSSV._NLRj:H5VRL8lFRR<=jsRFRFLl8RR>.o2RCsMCN
0CRSRRS1MFE0HVRR<= 5XaAHbslRC,N8IHCI+LH28C;R
RRRRRCRM8oCCMsCN0R_HVNj.L;S
SHNV_.:L4RRHV5FLl8RR=4o2RCsMCN
0CRSRRS1MFE0HVRR<= 5XaAHbsl&CRR''j,IRNH+8CL8IHC
2;RRRRRMRC8CRoMNCs0HCRV._NL
4;SVSH_LN..H:RVLR5lRF8=2R.RMoCC0sNCR
RRMSSFH1EV<0R=XR ab5AsCHlR'&Rj&'RR''j,IRNH+8CL8IHC
2;RRRRRMRC8CRoMNCs0HCRV._NL
.;RSRS#VEH0RC8<M=RFH#EVN05ICH8+HLI8.C-RI8FMR0Fj&2RR''j;S
SNC888RRR<M=RFH1EV+0RRH#EV80C;R
RRCS)#0kDN=R<RhBmea_17m_pt_QBea Bmj)5,HNI8LC+ICH82ERIC5MRC=4RRj"j"S2
SSSSRDRC#MCRFH1EVI0RERCM5RC4=jR"4
"2SSSSSCRRDR#C#VEH0RC8IMECR45CR"=R42j"
SSSSRSRCCD#R8N8C
8;S8CMRMoCC0sNCVRH_;N.
-
S-kRvDb0HDL$R$ER0CGRC0RsNL#H0RRHVIECRNRPCFRMCF0sRICFRGN0sR0LH#VRFRSA
HLV_4H:RVLR5lRF8=2R4RMoCC0sNCS
SHLV_4:NjRRHV5FNl8=R<RFjRslRNF>8RRR.2oCCMsCN0
SSS)kC#DR0L<B=Rm_he1_a7pQmtB _eB)am5Rj,N8IHCI+LH28CRCIEMCR5.25jR'=RjR'2
SSSSRSSR#CDCXR ab5qsCHl,IRNH+8CL8IHC
2;RRRRRMRC8CRoMNCs0HCRV4_LN
j;SVSH_NL44H:RVNR5lRF8=2R4RMoCC0sNCS
SS#)CkLD0RR<=Bemh_71a_tpmQeB_ mBa),5jRHNI8LC+ICH82ERIC5MRCj.52RR='2j'RS
SSSSSRDRC# CRXqa5blsHCRR&',j'RHNI8LC+ICH82R;
RRRRR8CMRMoCC0sNCVRH_NL44S;
S_HVL.4N:VRHRl5NF=8RRR.2oCCMsCN0
SSS)kC#DR0L<B=Rm_he1_a7pQmtB _eB)am5Rj,N8IHCI+LH28CRCIEMCR5.25jR'=RjR'2
SSSSRSSR#CDCXR ab5qsCHlR'&Rj&'RR''j,IRNH+8CL8IHC
2;RRRRRMRC8CRoMNCs0HCRV4_LN
.;S8CMRMoCC0sNCVRH_;L4
VSH_:L.RRHV5FLl8RR=.o2RCsMCN
0CRRRRRHR#oDMNR1MFE0HV,ER#HCV08N,R888CR#:R0D8_FOoH_OPC05FsN8IHCI+LH-8C4FR8IFM0R;j2
CSLo
HMSVSH_NL.jH:RVNR5lRF8<j=RRRFsN8lFR.>R2CRoMNCs0RC
RSRSMEF1HRV0< =RXqa5blsHCN,RICH8+HLI8;C2
RRRRCRRMo8RCsMCNR0CHLV_.;Nj
HSSV._LNR4:H5VRN8lFR4=R2CRoMNCs0RC
RSRSMEF1HRV0< =RXqa5blsHCRR&',j'RHNI8LC+ICH82R;
RRRRR8CMRMoCC0sNCVRH_NL.4S;
S_HVL..N:VRHRl5NF=8RRR.2oCCMsCN0
RRRSFSM1VEH0=R<Ra X5sqbHRlC&jR''RR&',j'RHNI8LC+ICH82R;
RRRRR8CMRMoCC0sNCVRH_NL..S;
SH#EV80CRR<=MEF1H5V0N8IHCI+LH-8C.FR8IFM0RRj2&jR''R;
RRRRR8N8CR8RRR<=MEF1HRV0+ER#HCV08S;
S#)CkLD0RR<=Bemh_71a_tpmQeB_ mBa),5jRHNI8LC+ICH82ERIC5MRC=.RRj"j"S2
SSSSRDRC#MCRFH1EVI0RERCM5RC.=jR"4
"2SSSSSCRRDR#C#VEH0RC8IMECR.5CR"=R42j"
SSSSRSRCCD#R8N8C
8;S8CMRMoCC0sNCVRH_;L.
-
S-kRvDb0HD0$RECCRGN0sR0LH#FR0oEC0CHsRVCRIRPENCGRC0#sNRRHMqMRN8
RAS_HVCR#:H5VR5FNl8R=4FNsRl=F8.N2RM58RL8lF=F4RslRLF.8=2o2RCsMCN
0CSCS)#0kDC25dRR<=C4452MRN84RC5Rj2NRM8C4.52MRN8.RC5;j2
)SSCD#k0.C52=R<R45C5R42NRM850MFR5C4jR22NRM8C4.52F2RsS
SSSSSRCR54254R8NMR5C.4N2RM58RMRF0Cj.52;22
)SSCD#k04C52=R<R45C5R42NRM850MFR5C.4R22NRM8Cj.52F2RsS
SSSSSRCR54254R8NMRF5M04RC52j2R8NMR5C.jR22FSs
SSSSS5RR50MFR5C44R22NRM8Cj452MRN8.RC5242R
FsSSSSSRSR55C4jN2RMC8R.254R8NMRF5M0.RC52j22S;
S#)CkCD05Rj2<C=R425jR8NMR5C.j
2;SVSH_#sCCH:RVNR5ICH8+HLI8>CRRRc2oCCMsCN0
SSS)kC#D50CN8IHCRR+L8IHCRR-4FR8IFM0RRc2<B=Rm_he1_a7pQmtB _eB)am5Rj,N8IHCI+LHR8C-;c2
CSSMo8RCsMCNR0CHsV_C;#C
MSC8CRoMNCs0HCRV#_C;S

LDlk0H:RVIRNHR8C>RR.NRM8L8IHCRR>.CRoMNCs0SC
SDlk0RGG:.ReABpmiS
SSMoCCOsHRblNRS5
SSSSSHNI8R0E=N>RI,H8
SSSSLSSI0H8E>R=RHLI8S,
SSSSSCMC8H_bbHCDM=CR>CRMCb8_HDbCH2MC
SSSb0FsRblNRS5
SSSSqRRRRR=>qHbsl
C,SSSSSRARR>R=RsAbH,lC
SSSS)Sum=7R>ER1Fus02S;
CRM8oCCMsCN0RkLlD
0;
GSC08CMHR0:bOsFCR##5F1Es20u
CSLoRHMRR--bOsFCR##CCG0M08H
)SSCD#k0<4R=XR aE51Fus0,IRNH+8CL8IHC
2;S8CMRFbsO#C#R0CGCHM80
;
SlNLF:8jRRHV5FNl8R>.FNsRl=F8jN2RM58RL8lF>F.RslRLFj8=2CRoMNCs0SC
S#)CkGD0RR<=)kC#D;04
MSC8CRoMNCs0NCRL8lFj
;
RNRSL8lF4H:RVNR5l=F84MRN8LR5l>F8.sRFRFLl82=j2sRFRN55l>F8.sRFRFNl82=jR8NMRFLl82=4RMoCC0sNCS
S)kC#DR0G<)=RCD#k0N45ICH8+HLI8.C-RI8FMR0Fj&2RR''j;C
SMo8RCsMCNR0CNFLl8
4;
LSNl.F8:VRHRl5NF48=R8NMRFLl82=4RRFs5FNl8R=.NRM85FLl8R>.FLsRl=F8jR22F5sR5FNl8R>.FNsRl=F8jN2RML8Rl=F8.o2RCsMCN
0CSCS)#0kDG=R<R#)Ck4D05HNI8LC+ICH8-8dRF0IMF2RjR"&Rj;j"
MSC8CRoMNCs0NCRL8lF.
;
SlNLF:8dRRHV5FNl8R=.NRM8L8lF=R42F5sRN8lF=N4RML8Rl=F8.o2RCsMCN
0CSCS)#0kDG=R<R#)Ck4D05HNI8LC+ICH8-8cRF0IMF2RjR"&Rj"jj;C
SMo8RCsMCNR0CNFLl8
d;
SRRNFLl8Rc:H5VRN8lF=N.RML8Rl=F8.o2RCsMCN
0CSCS)#0kDG=R<R#)Ck4D05HNI8LC+ICH8-86RF0IMF2RjR"&Rjjjj"S;
CRM8oCCMsCN0RlNLF;8c
H
SVC_oMNCs0RC:H5VR5l5NF>8RRRj2NRM85FNl8RR<dR22F5sR5FLl8RR>jN2RM58RL8lFRd<R2R22oCCMsCN0
CSLo
HMSVSH_N#00:C4RRHV5l5NF>8RRRj2NRM85FNl8RR<dN2RM58RL8lFRj>R2MRN8LR5lRF8<2Rd2CRoMNCs0SC
SsSuF_84NRkG<R=R)kC#DR0N+CR)#0kDLRR+)kC#D;0C
CSSMo8RCsMCNR0CH#V_0CN04S;
S_HV#00NCR.:H5VR5FNl8RR>jN2RM58RN8lFRd<R2MRN85R5L8lFR.>R2sRFRl5LF=8RR2j22CRoMNCs0SC
SsSuF_84NRkG<R=R)kC#D;0N
CSSMo8RCsMCNR0CH#V_0CN0.S;
S_HV#00NCRd:H5VR5FLl8RR>jN2RM58RL8lFRd<R2MRN85R5N8lFR.>R2sRFRl5NF=8RR2j22CRoMNCs0SC
SsSuF_84NRkG<R=R)kC#D;0L
CSSMo8RCsMCNR0CH#V_0CN0d
;
SVSH_bbH4H:RVMR5C_C8bCHbDCHMR4=R2CRoMNCs0SC
SkSLV0Fkb:k0RsVFRHHRMRRj0NFRI0H8ERR+L8IH04E-RMoCC0sNCS
SS0SN0LsHkR0C\N3sMR	\FsVRC1o#RD:RNDLCRRH#4S;
SNSS0H0sLCk0RL\3CMoH_C0sCF\RVCRsoR#1:NRDLRCDH4#R;S
SS0SN0LsHkR0C\C3slCFP__MFIMNs\VRFRosC#:1RRLDNCHDR#;R4
SSSLHCoMS
SSCSso:#1RHRbbkCLVS
SSFSbsl0RN
b5SSSSSRSQ=u>Rs4F8_GNk5,H2
SSSSmSSRR=>u8sF4C_s#25H
SSSS2SS;S
SS8CMRMoCC0sNCkRLV0Fkb;k0
CSSMo8RCsMCNR0CHbV_H;b4
HSSVH_bbRj:H5VRM8CC_bbHCMDHCRR=jo2RCsMCN
0CSuSSs4F8_#sC5HNI8R0E+IRLHE80R4-RRI8FMR0Fj<2R=SR
SuSSs4F8_GNk5HNI8R0E+IRLHE80R4-RRI8FMR0FjR2;
CSSMo8RCsMCNR0CHbV_H;bj
S
Su8sF4=R<R#)CkGD0Ru+Rs4F8_#sC;C
SMo8RCsMCNR0CHoV_CsMCN;0C
H
SVC_oMNCs04C_:VRHRN55lRF8>2R.R8NMRl5LF>8RR2.2RMoCC0sNCS
Su8sF4=R<R#)CkGD0;C
SMo8RCsMCNR0CHoV_CsMCN_0C4
;
RC
SGM0C8Fbs8b:RsCFO#5#Ru8sF4S2
LHCoM-RR-sRbF#OC#GRC08CMb8sF
HSSVHRI8R0E>IRNHR8C+IRLHR8C0MEC
SSSu8sF.=R<Ra X5Fus8R4,I0H8E
2;SDSC#SC
SsSuFR8.<u=Rs4F858IH04E-RI8FMR0Fj
2;SMSC8VRH;C
SMb8RsCFO#C#RGM0C8Fbs8
;
S_HVbNHb4H:RVMR5C_C8bCHbDCHMR4=R2CRoMNCs0SC
SVLkFbk0kR0:VRFsHMRHR0jRFHRI8-0E4CRoMNCs0SC
S0SN0LsHkR0C\N3sMR	\FsVRC1o#RD:RNDLCRRH#.S;
S0SN0LsHkR0C\M3C8s_0CRC\FsVRC1o#RD:RNDLCRRH#.S;
S0SN0LsHkR0C\F3b8\ClRRFVs#Co1RR:DCNLD#RHR
H;SNSS0H0sLCk0Rb\3Fl8CL\k#RRFVs#Co1RR:DCNLD#RHR)"um;7"
SSSNs00H0LkC3R\sFClPMC_FN_IsRM\FsVRC1o#RD:RNDLCRRH#4S;
SoLCHSM
SCSso:#1RHRbbkCLVS
SSFSbsl0RN
b5SSSSSRSQ=u>Rs.F85,H2
SSSSmSSRR=>u7)m5
H2SSSS2S;
S8CMRMoCC0sNCkRLV0Fkb;k0
MSC8CRoMNCs0HCRVH_bb;N4
VSH_bbHNRj:H5VRM8CC_bbHCMDHCRR=jo2RCsMCN
0CS)Sum<7R=sRuF58.I0H8ER-48MFI0jFR2S;
CRM8oCCMsCN0R_HVbNHbj
;
CRM8LODF	k_lD
0;




