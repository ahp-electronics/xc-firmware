
@ER--vkF8D:CRROkbM30sPRE8
-
-RMwkOF0HMk:RbFROkCM0sFRl8CkDRMoCC0sNF
sR
R--
-
-RMtCCOsH#
R
-I-RHE80RM-RkClLsVRFRkOFMs0CR0LH#
R
-s-RC0#CbRN0-CRs#RC0b0N0CRsMVRFsCENOR0LHR-

-0R#8F_Do_HOP0COFIs5HE80RI8FMR0FjR2,C33oRj"jjRj"
-
-Ru MFRDN-FRbDHNs0F$RVhR RMbHR-

-RRjNHO0PDCRF
IR
R--4ORN0CHPRoEHE
R
-.-RRRMF 5hROODF	DRNI#N$RNCML8DC2
R
-B-RDFsuD-NRRDbFN0sH$VRFR1)  baRH
MR
R--jORN0CHPRIDFR-

-RR4NHO0PECRHRoE
-
-RM.RF R)1R a5RMFsCC#0HRbM
2R
R--pF8uD-NRRDbFN0sH$VRFRqpm7HRbM
R
-j-RR0NOHRPCDRFI
-
-RN4ROP0HCHREo
ER
R--.FRMRqpm7NR5D$IN#FROkHM0MRo2
-
-R	BD C8oRN-ROP0HC8RCoFCRVpRBi
R
-j-RRDVNDoHMRoC8C
R
-4-RR#sHHRMoCC8oR-

-bRz7MFI7RHs-FROkRM08CHsOF0HM
R
-j-RRkOFM80RFRIM
-
-RO4RF0kMRRkb
-
-R-

-FRusR0#
-
-Ra7qqRR-8NN0RbHMkR0#VRFs#O$MEMsFFRk#D8FNR-

-RRT-FROkCM0skRF00bk#
R
-p-RmRq7-MRCNCLDRM#$OFEsM#FkRNDF8ERICNMROP0HC
,R
R--CCD#RNCMLRDCOMFk0oHMRb5F0MHFNVDRk0MOH2FMR-

-hR RC-RMDNLCDROFRO	IMECR0NOHRPC50FbHNFMDkRVMHO0FRM2
-
-R1)  -aRR$N#MsOEFkMF#CRs#RC050FbHNFMDkRVMHO0FRM2
-
-RiBpRO-RD	FORbHMk
0R
R--BamzRO-RN$ssR0FkbRk0
-
-RhBQRO-RN$ssRbHMk
0R
R--zhu7RE-RNIs8H8sCRR0F'R4'
-
-R-

--R----------------------------------------------------------R--



DsHLNRs$HCCC;kR
#HCRC3CC#_08DHFoO4_4nNc3DRD;
Ck#RsIF	C3oMObN	CNo3DND;
R

M
C0$H0RBzuhRa)H
#R
MoCCOsH58IH0:ERR0HMCsoCRR:=.
;R
#sCCN0b0RR:OMFk0ICsFRs8:j=R;-R-R8#0_oDFHPO_CFO0sH5I8-0E4FR8IFM0RRj2
s--C0#CbRN0:MRH0CCos=R:RRj;-#-R0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2
R
 FMuD:NRR0HMCsoCRR:=4-;R-,Rj4R,.NHO0PDCRFRI,EEHo,FRMM
CR
sBDuNFDRH:RMo0CC:sR=;R4RR--j,,4.ORN0CHPRIDF,HREoRE,MCFMRp

8DuFNRR:HCM0oRCs:4=R;-R-R4j,,N.ROP0HCFRDIE,RH,oERMMFC
R
B D	8RoC:MRH0CCos=R:RR4;-j-R,s4RHM#HoV,RNHDDMCoR8RoC
b
z7MFI7RHs:MRH0CCos=R:R-4R-,Rj4FROkRM08MFI,bRkR2

;
R
b0Fs5a7qqRR:H#MR0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2
;R
:TRR0FkR8#0_oDFHPO_CFO0sH5I8-0E4FR8IFM0R;j2Rp

mRq7:MRHR8#0_oDFHRO;
h
 RH:RM0R#8F_Do;HOR)

 a1 :MRHR8#0_oDFHRO;
p
BiRR:H#MR0D8_FOoH;
R
BamzRF:Rk#0R0D8_FOoH;
R
BRQh:MRHR8#0_oDFHRO;
u
z7:hRRRHM#_08DHFoO
R
2
;R
8CMRBzuh;a)RN

sHOE00COkRsCpze_uaBh)R_)FzVRuaBh)#RH
F
OlMbFCRM0z_Bup
1ARbRRF5s0
RRRR7RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR:RRHMR1RRap7_mBtQ;R
RRRRR1R7RRRRRRRRRRRRRRRRRRRRRRRRRR:RRRMRHRRRR1_a7pQmtBR;
RRRRRqpm7RRRRRRRRRRRRRRRRRRRRRRRRRRR:HRRMRRRR71a_tpmQ
B;RRRRRYRBQ)AqRRRRRRRRRRRRRRRRRRRRRRRRRR:RHRMRRaR17m_pt;QB
RRRR1RRjRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR:R0FkR1RRap7_mBtQ;R
RRRRRBamzRRRRRRRRRRRRRRRRRRRRRRRRR:RRRkRF0RRR1_a7pQmtB
2;CRM8ObFlFMMC0
;
ObFlFMMC0BRBzB_zuR
RRsbF0R5
RRRRRR7RRRRRRRRRRRRRRRRRRRRRRRRRRRRR:HRRMRRRR71a_tpmQ
B;RRRRR7R1RRRRRRRRRRRRRRRRRRRRRRRRRRRRRR:RHRMRRaR17m_pt;QB
RRRRpRRmRq7RRRRRRRRRRRRRRRRRRRRRRRRRRR:RRHMR1RRap7_mBtQ;R
RRRRRBRQhRRRRRRRRRRRRRRRRRRRRRRRRR:RRRMRHRRRR1_a7pQmtBR;
RRRRRR1jRRRRRRRRRRRRRRRRRRRRRRRRRRRR:FRRkR0RR71a_tpmQ
B;RRRRRmRBzRaRRRRRRRRRRRRRRRRRRRRRRRRRRR:RFRk0RaR17m_pt2QB;M
C8FROlMbFC;M0
F
OlMbFCRM07BwwA
)]RbRRF5s0
RRRRBRR RRRRRRRRRRRRRRRRRRRRRRRRRRRRRR:RRHMR1RRap7_mBtQ;R
RRRRR7RRRRRRRRRRRRRRRRRRRRRRRRRRRR:RRRMRHRRRR1_a7pQmtBR;
RRRRRiBpRRRRRRRRRRRRRRRRRRRRRRRRRRRR:HRRMRRRR71a_tpmQ
B;RRRRRRR)RRRRRRRRRRRRRRRRRRRRRRRRRRRRRR:RHRMRRaR17m_pt;QB
RRRRTRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR:R0FkR1RRap7_mBtQ2C;
MO8RFFlbM0CM;


ObFlFMMC0wR7w1BA]R
RRsbF0R5
RRRRRRB RRRRRRRRRRRRRRRRRRRRRRRRRRRR:HRRMRRRR71a_tpmQ
B;RRRRRRR7RRRRRRRRRRRRRRRRRRRRRRRRRRRRRR:RHRMRRaR17m_pt;QB
RRRRBRRpRiRRRRRRRRRRRRRRRRRRRRRRRRRRRR:RRHMR1RRap7_mBtQ;R
RRRRR1RRRRRRRRRRRRRRRRRRRRRRRRRRRR:RRRMRHRRRR1_a7pQmtBR;
RRRRRRTRRRRRRRRRRRRRRRRRRRRRRRRRRRRR:FRRkR0RR71a_tpmQ;B2
8CMRlOFbCFMM
0;
RRRRRRRRo#HMRNDOsNs$RR:#_08DHFoOC_POs0F5HRI8-0E4FR8IFM0R2jR;R
RRRRRRHR#oDMNR#T_H:oRR8#0_oDFHPO_CFO0sI5RHE80-84RF0IMFRRj2R;
RRRRR#RRHNoMD_R1#RHo:0R#8F_Do_HOP0COFRs5I0H8ER-48MFI0jFRR
2;RRRRRRRR#MHoNDDRFOoH4RRRR#:R0k8_DHFoO=R:R''4;R
RRRRRRHR#oDMNRoDFHROjR:RRR8#0_FkDoRHO:'=Rj
';RRRRRRRR#MHoNODRD#	_HRoRR#:R0k8_DHFoO=R:R''j;-RR-DROFRO	F
VVRRRRRRRR#MHoNODRD#s_HRoRR#:R0k8_DHFoO=R:R''j;-RR-DROCRNs8NH#L8DC
RRRRRRRRo#HMRNDC#M_HRoRRRR:#_08koDFH:OR=4R''R;R-O-RD	FORNCML8DC
RRRRRRRRo#HMRNDO_HM#RHoR:RRR8#0_FkDoRHO:'=RjR';RR--OODF	MRCNCLD8R
RRRRRRHR#oDMNR_D8#RHoR:RRR8#0_FkDoRHO:'=RjR';RR--D8FNR#8HNCLD8R
RRRRRRHR#oDMNR	OD__CM#RHoR:RRR8#0_FkDoRHO:'=RjR';RR--D8FNR#8HNCLD8L

CMoH
R
RRRRRRNRVDMDHoD_O	H:RVBR5D8	 o=CRRRj2oCCMsCN0
RRRRRRRRORRD#	_H<oR=FRM0pRBiR;
RRRRRCRRMo8RCsMCN;0C
RRRRRRRR#sHH_MoO:D	RRHV5	BD C8oR4=R2CRoMNCs0RC
RRRRRRRRR	OD_o#HRR<=B;pi
RRRRRRRR8CMRMoCC0sNCR;
RRRRRR
RRRRRRORN0CHP_IDF_sOD:VRHRD5BsDuFNRR=jo2RCsMCN
0CRRRRRRRRRDROsH_#o=R<R0MFR1)  
a;RRRRRRRRCRM8oCCMsCN0;R
RRRRRRORN0CHP_oEHED_OsH:RVBR5DFsuD=NRRR42oCCMsCN0
RRRRRRRRORRD#s_H<oR= R)1; a
RRRRRRRR8CMRMoCC0sNCR;
RRRRRMRRFD_OsH:RVBR5DFsuD=NRRR.2oCCMsCN0
RRRRRRRRORRD#s_H<oR=FRDojHO;R
RRRRRRMRC8CRoMNCs0
C;
RRRRRRR
RRRRRRRR0NOH_PCD_FIDR8:H5VRpF8uD=NRRRj2oCCMsCN0
RRRRRRRRDRR8H_#o=R<R0MFRqpm7S;
SCRRMH_#o=R<R; h
RSSRMOH_o#HRR<=BRQhNRM8D#8_H
o;RRRRRRRRCRM8oCCMsCN0;R
RRRRRRORN0CHP_oEHE8_D:VRHR85puNFDR4=R2CRoMNCs0RC
RRRRRRRRR_D8#RHo<p=Rm;q7
RSSR_CM#RHo< =RhS;
SORRH#M_H<oR=QRBhMRN8FRM08RD_o#H;R
RRRRRRMRC8CRoMNCs0
C;RRRRRRRRMDF_8H:RVpR58DuFNRR=.o2RCsMCN
0CRRRRRRRRR8RD_o#HRR<=DHFoO
j;SRSRC#M_H<oR=hR ;SR
SORRH#M_H<oR=QRBhR;
RRRRRCRRMo8RCsMCN;0C
S
SNHO0PDC_FOI_DC	_MH:RV R5MDuFNRR=jo2RCsMCN
0CRRRRRRRRRDRO	M_C_o#HRR<=C#M_H
o;RRRRRRRRCRM8oCCMsCN0;R
RRRRRRORN0CHP_oEHED_O	M_C:VRHRM5 uNFDR4=R2CRoMNCs0RC
RRRRRRRRR	OD__CM#RHo<M=RFC0RMH_#oR;
RRRRRCRRMo8RCsMCN;0C
RRRRRRRR_MFO_D	CRM:H5VR FMuD=NRRR.2oCCMsCN0
RRRRRRRRORRDC	_MH_#o=R<RoDFH;Oj
RRRRRRRR8CMRMoCC0sNC
;
S4Sz:BRBzB_zumRu)vaRq1u5j=RR>_R1#5HojR2,
SSSSSSSBamzRR=>OsNs$25j,SR
SSSSSRS7=T>R_o#H5,j2RS
SSSSSSR17=7>Rq5aqjR2,
SSSSSSSp7mqRR=>D#8_HRo,
SSSSSSSBRQh=O>RH#M_H;o2
S
SHoV_CRM:H5VRsCC#00bN5Rj2=jR''o2RCsMCN
0CSRRRRRRRR:z.Rw7wB]A)R)umaqRvuRR5RRRT=R>RTH_#o25j,RR
RRRSRRRRRRRRRRRRRRRRRRRRRRRRRRRRR=7R>1RR_o#H5,j2RR
RRRSRRRRRRRRRRRRRRRRRRRRRRRRRRpRBi>R=RDRO	H_#o
,RRSRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR)R=R>RO_Ds#,HoRR
RRRSRRRRRRRRRRRRRRRRRRRRRRRRRR RBR>R=RDRO	M_C_o#HR
2;SMSC8CRoMNCs0HCRVC_oM
;
SVSH_MoC4H:RVsR5C0#Cb5N0j=2RR''42CRoMNCs0SC
RRRRRRRRz:.NRw7wB]A1R)umaqRvuRR5RRRT=R>RTH_#o25j,RR
RRRSRRRRRRRRRRRRRRRRRRRRRRRRRRRRR=7R>1RR_o#H5,j2RR
RRRSRRRRRRRRRRRRRRRRRRRRRRRRRRpRBi>R=RDRO	H_#o
,RRSRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR1R=R>RO_Ds#,HoRR
RRRSRRRRRRRRRRRRRRRRRRRRRRRRRR RBR>R=RDRO	M_C_o#HR
2;SMSC8CRoMNCs0HCRVC_oM
4;
RRRRRRRR:p4RsVFRHHRMRR40IFRHE80-o4RCsMCN
0CRRRRRRRRRRRRRRRRpz4_4B:RBzz_BuuRmR)av5qu1RjR=1>R_o#H5,H2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRzBma>R=RsONsH$52
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR7=T>R_o#H5,H2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR1RR7>R=Ra7qq25H,RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRmRpq=7R>8RD_o#H,RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRBRRQ=hR>NROs5s$H2-42S;
SVSH_MoCGH:RVsR5C0#Cb5N0H=2RR''j2CRoMNCs0RC
RRRRRRRRRRRRRpRR4._z:wR7w)BA]mRu)vaRq5uRT=RR>_RT#5HoHR2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR7RR=>1H_#o25H,RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRBRRp=iR>DRO	H_#o
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR)R=O>RD#s_HRo,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRB RR=>O_D	C#M_H2oR;S
SS8CMRMoCC0sNCVRH_MoCGS;
SVSH_MoC$H:RVsR5C0#Cb5N0H=2RR''42CRoMNCs0RC
RRRRRRRRRRRRRpRR4W_z:wR7w1BA]mRu)vaRq5uRT=RR>_RT#5HoHR2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR7RR=>1H_#o25H,RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRBRRp=iR>DRO	H_#o
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR1R=O>RD#s_HRo,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRB RR=>O_D	C#M_H2oR;S
SS8CMRMoCC0sNCVRH_MoC$R;
RRRRRCRRMo8RCsMCN;0C
R
RRRRRRRRT<T=R_o#H;R
RRRRRRmRBz<aR=NROs5s$I0H8E2-4;C

Mp8Reu_zB)ha_
);
