--
@ER--B$FbsEHo0OR52gR4g-cRRj.jd$R1MHbDO$H0ROQM
R--fN]C8:CsR#//$DMbH0OH$N/lb0DN.Uj4J4.b/blNb#Cs/0N0/LDH/MoC_OFsN/.Ns_NlsPI3E48yR-f
-


---
-HR1lCbDRv)qR0IHEHR#MCoDR7q7)1 1RsVFR0LFECRsNN8RMI8RsCH0
R--aoNsC:0RROpkCRM0-)RmB.qRq-
-

--
LDHs$NsRCHCCk;
#HCRC3CC#_08DHFoO4_4nNc3D
D;kR#CHCCC38#0_oDFH#O_HCoM8D3NDD;
HNLssF$Rs.ON;#
kCsRFO3N.FNsOObFl3DND;M
C0$H0Rv)q_R)WHR#
RoRRCsMCH5OR
RRRRRRRRlVNH:D$Rs#0HRMo:"=RMCFM"R;
RRRRRIRRHE80RH:RMo0CC:sR=;R4RR
RRRRRR8RN8HsI8R0E:MRH0CCos=R:RRc;RRRRR-RR-HRLoMRCFEkoRsVFRb8C0RE
RRRRR8RRCEb0RH:RMo0CC:sR=4RRnR;
RRRRR8RRF_k0sRCo:FRLFNDCM=R:RDVN#RC;RRRR-E-RNF#Rkk0b0CRsoR
RRRRRRHR8MC_soRR:LDFFCRNM:V=RNCD#;RRRR-RR-NRE#NR80HNRM0bkRosC
RRRRRRRR8N8sC_soRR:LDFFCRNM:V=RNCD#RRRRR-R-R8ENR8N8s#C#RosC
RRRRRRRR
2;RRRRb0FsRR5
RRRRR7RRmRza:kRF00R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj;R
RRRRRRQR7h:RRRRHM#_08DHFoOC_POs0F58IH04E-RI8FMR0Fj
2;RRRRRRRRq)77RH:RM0R#8F_Do_HOP0COFNs58I8sHE80-84RF0IMF2Rj;R
RRRRRR RWRRR:H#MR0D8_FOoH;RRRRRRR-I-RsCH0RNCMLRDCVRFss
NlRRRRRRRRBRpi:MRHR8#0_oDFHRO;RRRRR-R-RFODOV	RFssRNRl,Ns88,HR8MR
RRRRRRBRmp:iRRRHM#_08DHFoORRRRRRR-F-RbO0RD	FORsVFRk8F0R
RRRRRR;R2
8CMR0CMHR0$)_qv)
W;

---w-RH0s#RbHlDCClM00NHRFMl0k#RRLCODNDCN8RsjOE

--NEsOHO0C0CksRONsEFjRVqR)vW_)R
H#O#FM00NMRlMk_DOCD8#_CRCb:MRH0CCos=R:R855CEb0R4-R2n/42R;RRRRRRR--yVRFRIsF#VRFRw)B4cnXZCRODRD#M8CCCO8
F0M#NRM0M_klODCD#H_I8:CRR0HMCsoCRR:=5H5I8R0E-2R4/;c2RRRRRRRR-y-RRRFVOkFDlRM#F)VRBnw4XRcZODCD#CRMC88C
0--$RbCF_k0L_k#0C$bRRH#NNss$MR5kOl_C#DDRI8FMR0FjI,RHE80-84RF0IMF2RjRRFV#_08DHFoO-;
-o#HMRNDF_k0LRk#:kRF0k_L#$_0bRC;RRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFRk8F0HR5M0bkRR0F0-sH#00NC
#2#MHoNFDRkC0_MRR:#_08DHFoOC_POs0F5lMk_DOCD8#_CRCb8MFI0jFR2R;RRRRRR-R-RNCML#DCRsVFRH0s-N#00
C##MHoNIDRbCC_MRR:#_08DHFoOC_POs0F5lMk_DOCD8#_CRCb8MFI0jFR2R;RRRRRR-R-RHIs0CCRMDNLCV#RFCsRNROEsRFIF)VRqOvRC#DD
o#HMRNDHsM_C:oRR8#0_oDFHPO_CFO0sH5I8+0EdFR8IFM0R;j2RRRRRRRRR-R-RCk#8FR0RosCHC#0sQR7h#R
HNoMDkRF0C_soRR:#_08DHFoOC_POs0F58IH0dE+RI8FMR0FjR2;RRRRRRRR-k-R#RC80sFRC#oH0RCs7amz
o#HMRNDNs8_C:oRR8#0_oDFHPO_CFO0s85N8HsI8-0E4FR8IFM0R;j2RRRRR-R-RCk#8FR0RosCHC#0s7Rq7#)
HNoMDFRDI8_N8:sRR8#0_oDFHPO_CFO0sR5d8MFI0jFR2R;RRRRRRRRRRRRR-N-R8R8sL#H0RbHMk00RFqR)vCRODRD#5LcRHR0#skCJH8sC2L

CMoH
R
RR-R-RRQVNs88I0H8ERR<c#RN#MHoR''jRR0Fk#MkCL8RH
0#RRRRzR4R:VRHR85N8HsI8R0E=2R4RMoCC0sNCR
RRRRRRFRDI8_N8<sR=jR"jRj"&8RN_osC5;j2
RRRR8CMRMoCC0sNC4Rz;R
RR.RzRRR:H5VRNs88I0H8ERR=.o2RCsMCN
0CRRRRRRRRD_FINs88RR<=""jjRN&R8C_soR548MFI0jFR2R;
RCRRMo8RCsMCNR0Cz
.;RRRRzRdR:VRHR85N8HsI8R0E=2RdRMoCC0sNCR
RRRRRRFRDI8_N8<sR=jR''RR&Ns8_C.o5RI8FMR0Fj
2;RRRRCRM8oCCMsCN0R;zd
RRRRRzcRH:RVNR58I8sHE80Rd>R2CRoMNCs0RC
RRRRRDRRFNI_8R8s<N=R8C_soR5d8MFI0jFR2R;
RCRRMo8RCsMCNR0Cz
c;
RRRRR--Q5VR8_HMs2CoRosCHC#0sQR7h#RkHRMoB
piRRRRzR6R:VRHRH58MC_soo2RCsMCN
0CRRRRRRRRbOsFCR##5iBp,QR7hL2RCMoH
RRRRRRRRRRRRRHV5iBpR'=R4N'RMB8RpCi'P0CM2ER0CRM
RRRRRRRRRRRRRHRRMC_so=R<Rj5"j"jjR7&RQ;h2
RRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMRFbsO#C#;R
RRMRC8CRoMNCs0zCR6R;
RzRRn:RRRRHV50MFRM8H_osC2CRoMNCs0RC
RRRRRRRRRHRRMC_so=R<Rj5"j"jjR7&RQ;h2
RRRR8CMRMoCC0sNCnRz;R

R-RR-VRQRF58ks0_CRo2sHCo#s0CRz7ma#RkHRMomiBp
RRRRRz(RH:RV8R5F_k0s2CoRMoCC0sNCR
RRRRRRsRbF#OC#mR5B,piR0Fk_osC2CRLo
HMRRRRRRRRRRRRH5VRmiBpR'=R4N'RMm8RB'piCMPC002RE
CMRRRRRRRRRRRRRRRR7amzRR<=F_k0s5CoI0H8ER-48MFI0jFR2R;
RRRRRRRRRCRRMH8RVR;
RRRRRCRRMb8RsCFO#
#;RRRRRRRRCRM8oCCMsCN0R;z(
RRRRRzURH:RVMR5F80RF_k0s2CoRMoCC0sNCR
RRRRRRRRRRmR7z<aR=kRF0C_soH5I8-0E4FR8IFM0R;j2
RRRR8CMRMoCC0sNCURz;R

R-RR-VRQR85N8ss_CRo2sHCo#s0CR7q7)#RkHRMoB
piRRRRzRgR:VRHR85N8ss_CRo2oCCMsCN0
RRRRRRRRFbsO#C#Rp5Biq,R727)RoLCHRM
RRRRRRRRRHRRVBR5p=iRR''4R8NMRiBp'CCPMR020MEC
RRRRRRRRRRRRRRRR_N8sRCo<q=R757)Ns88I0H8ER-48MFI0jFR2R;
RRRRRRRRRCRRMH8RVR;
RRRRRCRRMb8RsCFO#
#;RRRRCRM8oCCMsCN0R;zg
RRRRjz4RH:RVMR5FN0R8_8ss2CoRMoCC0sNCR
RRRRRRRRRR8RN_osCRR<=q)77;R
RRMRC8CRoMNCs0zCR4
j;RRRRRRRR
RRRRR--tCCMsCN0RC0ERv)qRDOCDN#RM#8RCODC0FRDo
HORRRRzR44:FRVsRRHHMMRkOl_C#DD_C8CbFR8IFM0RojRCsMCN
0CRRRR-Q-RVNR58I8sHE80Rc>R2CRMC08RFsROCCN0RHIs0CCRMDNLCMRN8kRF00bkRNCMLRDC#CCDOD0RFOoH
RRRRRRRR.z4RH:RVNR58I8sHE80Rc>R2CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_M25HRR<='Rj'IMECR85N_osC58N8s8IH04E-RI8FMR0Fc=2RRRH2CCD#R''4;R
RRRRRRRRRRRRRRbRICM_C5RH2<'=R4I'RERCM5_N8s5CoNs88I0H8ER-48MFI0cFR2RR=HC2RDR#C';j'
RRRRRRRRRRRR8CMRMoCC0sNC4Rz.R;
R-RR-VRQR85N8HsI8R0E<c=R2FRMRHIs0CCRMDNLCsRFR0FkbRk0CLMND#CRCODC0FRDoRHOM8CCCR8
RzRR4:dRRRHV58N8s8IH0<ER=2RcRMoCC0sNCR
RRRRRRRRRRkRF0M_C5RH2<'=Rj
';RRRRRRRRRRRRRRRRI_bCCHM52=R<R''4;R
RRRRRRRRRRMRC8CRoMNCs0zCR4
d;RRRR-t-RMNCs00CRE)CRqOvRC#DDR0IHEsR0H0-#N#0C
RRRRRRRRcz4RV:RF[sRRRHMM_klODCD#H_I88CRF0IMFRRjoCCMsCN0
RRRRRRRRRRRRqz)v):RBnw4XRcZ
RRRRRRRRRRRRsbF0NRlbaR5)=QR>kRF0M_C5,H2Rj7QRR=>HsM_C5o5c2*[27,RQ=4R>MRH_osC5*5c[42+27,RQ=.R>MRH_osC5*5c[.2+2
,RRRRRRRRRRRRRRRRRRRRRRRRRRQR7d>R=R_HMs5Co5[c*22+d,7Rqj>R=RIDF_8N8s25j,7Rq4>R=RIDF_8N8s254,7Rq.>R=RIDF_8N8s25.,R
RRRRRRRRRRRRRRRRRRRRRRRRRqR7d=D>RFNI_858sdR2,Wh) RR=>WR ,WRu =I>RbCC_M25H,iRBRR=>B,piRj7mRR=>F_k0s5Co5c[*2
2,RRRRRRRRRRRRRRRRRRRRRRRRRmR74>R=R0Fk_osC5*5[c42+27,Rm=.R>kRF0C_so[55*+c2.R2,7Rmd=F>Rks0_C5o5[2*c+2d2;R
RRRRRRRRRRMRC8CRoMNCs0zCR4
c;RRRRRRRRCRM8oCCMsCN0R4z4;R
RRRRRRRRRRRRRRRRRRRRRRRRRR
RRCRM8NEsOHO0C0CksRONsE
j;
