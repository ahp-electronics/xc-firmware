--$Header: //synplicity/maplat2018q2p1/designware/dw04.vhd#1 $
@E---------------------------------------------------------------------------------------------------

---w-RHRDCRRRRR:RRRj8IcE3P8-
-R#7CHRoMRRRRRB:RFNM0HRM#4L6RNO#HR#7CHWoMNRsCObFlFMMC0
#R-B-RFNlbMR$RR:RRRM1$bODHHR0$Q3MO
R--7CN0RRRRRRRR:kRqo6R.,jR.j
UR-q-RkF0EsRRRR:RRRD1CPRNl)-R
-CResF#HMRRRRRR:d
34---
-------------------------------------------------------------------------------------------------D-
HNLssQ$R ,  7)Wq W,7j
c;kR#CQ   38#0_oDFH4O_43ncN;DD
Ck#Rq7W)7 3WObN	CNo#D3NDk;
#7CRW3jc7cWj_lOFbCFMM30#N;DD
M
C0$H0Rj7WcN_bsC_oM#RH
MoCCOsHRH5I8R0E:hRQa  t)=R:RRU;b_Ns0C$bRQ:Rhta  :)R=2R4;b

FRs0508NNRHM:MRHR8#0_oDFHPO_CFO0sH5I8-0E4FR8IFM0R;j2
RRRRbRRN0sH$RR:FRk0#_08DHFoOR
RR;R2
-
-R0N0skHL08CRCNODsHN0FVMRF#sRHDMoCFR#kCsOR#8CHIoMN
sCRRRRRRRRNs00H0LkC$R#Mk_LHHD0Mk_8R#:R0MsHoR;
RRRRRNRR0H0sLCk0RM#$_HLkDM0H_R8kF7VRW_jcb_NsoRCM:MRC0$H0RRH#"NIC	
";
M
C8WR7jbc_Nos_C
M;
s
NO0EHCkO0ssCR0FDRVWR7jbc_Nos_CHMR#-

-0RN0LsHkR0C8DCON0sNHRFMVRFs#oHMD#CRFOksCCR8#MHoICNsR0
N0LsHkR0C#_$MLDkH0_HM8:kRRs#0H;Mo
0N0skHL0#CR$LM_k0HDH8M_kVRFRDs0RN:RsHOE00COkRsCH"#RI	CN"R;

R--wRFs#oHMD#CRFOksCWR7,sRNO0EHCkO0s#CREDFk8CRLRl8klN$
0H0sLCk0RM#$_NLDOL	_F:GRRFLFDMCN;0
N0LsHkR0C#_$MLODN	F_LGVRFRDs0RN:RsHOE00COkRsCH0#Rs;kC
L

CMoH
C

Ms8R0
D;
----------------------------------------------------------------------------------------D-
HNLssQ$R ,  7)Wq W,7j
c;kR#CQ   38#0_oDFH4O_43ncN;DD
Ck#Rq7W)7 3WObN	CNo#D3NDk;
#7CRW3jc7cWj_lOFbCFMM30#N;DD
M
C0$H0R_7WCROOHo#
CsMCH5ORI0H8ERR:Q hatR ):n=RcO;REH	L0:#RRaQh )t RR:=U#;R$_M8#RCD:hRQa  t)=R:R;j2
F
bs50RoRCM:MRHR8#0_oDFHRO;
RRRRORRFCssOM0_RH:RM0R#8F_Do;HO
RRRR8RRNH0NMRR:H#MR0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2R;
RRRRR	OEH:MRRRHM#_08DHFoOC_POs0F5	OEL#H0-84RF0IMF2Rj;R
RRRRRC_ss8CC0O:0RR0FkR8#0_oDFH
O;RRRRRsRCsk_lDD0bRF:Rk#0R0D8_FOoH;RR
RRRRR08NN0FkRF:Rk#0R0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2R;
RRRRR	OEFRk0:kRF00R#8F_Do_HOP0COFOs5EH	L04#-RI8FMR0Fj;22
-

-0RN0LsHkR0C8DCON0sNHRFMVRFs#oHMD#CRFOksCCR8#MHoICNs
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kRR:#H0sM
o;RRRRRRRRNs00H0LkC$R#Mk_LHHD0Mk_8RRFV7CW_O:ORR0CMHR0$H"#RI	CN"
;

8CMR_7WC;OO
N

sHOE00COkRsCsR0DF7VRWO_CO#RH
-
-R0N0skHL08CRCNODsHN0FVMRF#sRHDMoCFR#kCsOR#8CHIoMNRsC
0N0skHL0#CR$LM_k0HDH8M_kRR:#H0sM
o;Ns00H0LkC$R#Mk_LHHD0Mk_8RRFVsR0D:sRNO0EHCkO0sHCR#IR"C"N	;

R-w-RF#sRHDMoCFR#kCsOR,7WRONsECH0Os0kCER#F8kDRRLC8lkl$0
N0LsHkR0C#_$MLODN	F_LGRR:LDFFC;NM
0N0skHL0#CR$LM_D	NO_GLFRRFVsR0D:sRNO0EHCkO0sHCR#sR0k
C;
C
Lo
HM
M
C80RsD
;
---------------------------------------------------------------------------------------------------------
--
LDHs$NsR Q  W,7q,) 7cWj;#
kC RQ # 30D8_FOoH_n44cD3NDk;
#7CRW q)3b7WNNO	o3C#N;DD
Ck#Rj7WcW37jOc_FFlbM0CM#D3ND
;
CHM007$RWN_0b#RH
MoCCOsHRH5I8R0E:hRQa  t)=R:RRU;H:8RRaQh )t RR:=jP;
CHs#F:MRRaQh )t RR:=jb;RNRs0:hRQa  t)=R:R
j;l_NMMRkl:hRQa  t)=R:RRj;#O$M_8lFCRR:Q hatR ):j=RR
2;
sbF00R5O:	RRRHM#_08DHFoO0;Rs_#0MRR:H#MR0D8_FOoH;l
0#RR:H#MR0D8_FOoH;8R0HRR:H#MR0D8_FOoH;F
#RH:RM0R#8F_Do;HORbL$N_###:CDRRHM#_08DHFoO#;
CHM0M_CDPRND:MRHR8#0_oDFHPO_CFO0sH5I8-0E.FR8IFM0R;j2
FODO8	_sRR:FRk0#_08DHFoO#;RE0HV_R8s:kRF00R#8F_Do;HO
8kbN_0C8:sRR0FkR8#0_oDFHRO;0R8F:kRF00R#8F_Do;HO
F08_RCM:kRF00R#8F_Do;HO
b0N_N#00:CRR0FkR8#0_oDFHPO_CFO0s654RI8FMR0Fj
2;CCG0#:0RR0FkR8#0_oDFH
O;#bNl_NDF8RR:FRk0#_08DHFoOH;
Ms#0kHO0FRM#:kRF00R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj;$
#MOO_Nkb0sCC_MRR:FRk0#_08DHFoO#;
$_MOkNb808C_sRR:FRk0#_08DHFoO0;
CR#0:MRHR8#0_oDFH2OR;-

-0RN0LsHkR0C8DCON0sNHRFMVRFs#oHMD#CRFOksCCR8#MHoICNs
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kRR:#H0sM
o;RRRRRRRRNs00H0LkC$R#Mk_LHHD0Mk_8RRFV70W_N:bRR0CMHR0$H"#RI	CN"
;

8CMR_7W0;Nb
N

sHOE00COkRsCsR0DF7VRWN_0b#RH
-
-R0N0skHL08CRCNODsHN0FVMRF#sRHDMoCFR#kCsOR#8CHIoMNRsC
0N0skHL0#CR$LM_k0HDH8M_kRR:#H0sM
o;Ns00H0LkC$R#Mk_LHHD0Mk_8RRFVsR0D:sRNO0EHCkO0sHCR#IR"C"N	;

R-w-RF#sRHDMoCFR#kCsOR,7WRONsECH0Os0kCER#F8kDRRLC8lkl$0
N0LsHkR0C#_$MLODN	F_LGRR:LDFFC;NM
0N0skHL0#CR$LM_D	NO_GLFRRFVsR0D:sRNO0EHCkO0sHCR#sR0k
C;
C
Lo
HM
M
C80RsD
;

H
DLssN$ RQ 7 ,W q),j7Wck;
#QCR 3  #_08DHFoO4_4nNc3D
D;kR#C7)Wq W37b	NON#oC3DND;#
kCWR7j7c3W_jcObFlFMMC0N#3D
D;
0CMHR0$7LW_OR_4Hb#
FRs05bON0Cks_	ODRH:RM0R#8F_Do;HOR8kbN_0CORD	:MRHR8#0_oDFH
O;O0Nbk_sCC:MRRRHM#_08DHFoOk;Rb08NCM_CRH:RM0R#8F_Do;HO
H#EV80_sRR:H#MR0D8_FOoH;FRl8:CRRRHM#_08DHFoO#;
HRR:H#MR0D8_FOoH;NR80HN_MRR:H#MR0D8_FOoH;N
80FN_k:0RR0FkR8#0_oDFHRO;#:FRR0FkR8#0_oDFH2OR;-

-0RN0LsHkR0C8DCON0sNHRFMVRFs#oHMD#CRFOksCCR8#MHoICNs
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kRR:#H0sM
o;RRRRRRRRNs00H0LkC$R#Mk_LHHD0Mk_8RRFV7LW_OR_4:MRC0$H0RRH#"NIC	
";
8CMR_7WL4O_;


NEsOHO0C0CksRDs0RRFV7LW_OR_4H
#
-N-R0H0sLCk0RO8CDNNs0MHFRsVFRM#HoRDC#sFkO8CRCo#HMsINCNR
0H0sLCk0RM#$_HLkDM0H_R8k:0R#soHM;0
N0LsHkR0C#_$MLDkH0_HM8FkRV0RsDRR:NEsOHO0C0CksRRH#"NIC	
";R-
-RswFRM#HoRDC#sFkO7CRWN,RsHOE00COkRsC#kEFDL8RCkR8l
l$Ns00H0LkC$R#MD_LN_O	LRFG:FRLFNDCMN;
0H0sLCk0RM#$_NLDOL	_FFGRV0RsDRR:NEsOHO0C0CksRRH#0Csk;


LHCoMC

Ms8R0
D;
H
DLssN$ RQ 7 ,W q),j7Wck;
#QCR 3  #_08DHFoO4_4nNc3D
D;kR#C7)Wq W37b	NON#oC3DND;#
kCWR7j7c3W_jcObFlFMMC0N#3D
D;
0CMHR0$7LW_OR_.Hb#
FRs05bON0Cks_	ODRH:RM0R#8F_Do;HO
8kbN_0CORD	:MRHR8#0_oDFH
O;O0Nbk_sCC:MRRRHM#_08DHFoOk;
b08NCM_CRH:RM0R#8F_Do;HO
H#EV80_sRR:H#MR0D8_FOoH;F
l8:CRRRHM#_08DHFoO#;
HRR:H#MR0D8_FOoH;N
80HN_MRR:H#MR0D8_FOoH;N
80FN_k:0RR0FkR8#0_oDFH
O;#:FRR0FkR8#0_oDFH2OR;-

-0RN0LsHkR0C8DCON0sNHRFMVRFs#oHMD#CRFOksCCR8#MHoICNs
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kRR:#H0sM
o;RRRRRRRRNs00H0LkC$R#Mk_LHHD0Mk_8RRFV7LW_OR_.:MRC0$H0RRH#"NIC	
";
8CMR_7WL.O_;N

sHOE00COkRsCsR0DF7VRWO_L_H.R#-

-0RN0LsHkR0C8DCON0sNHRFMVRFs#oHMD#CRFOksCCR8#MHoICNsR0
N0LsHkR0C#_$MLDkH0_HM8:kRRs#0H;Mo
0N0skHL0#CR$LM_k0HDH8M_kVRFRDs0RN:RsHOE00COkRsCH"#RI	CN"R;

R--wRFs#oHMD#CRFOksCWR7,sRNO0EHCkO0s#CREDFk8CRLRl8klN$
0H0sLCk0RM#$_NLDOL	_F:GRRFLFDMCN;0
N0LsHkR0C#_$MLODN	F_LGVRFRDs0RN:RsHOE00COkRsCH0#Rs;kC
L

CMoH
8CMRDs0;


DsHLNRs$Q   ,q7W)7 ,W;jc
Ck#R Q  03#8F_Do_HO4c4n3DND;#
kCWR7q3) 7NWbOo	NCN#3D
D;kR#C7cWj3j7WcF_OlMbFC#M03DND;C

M00H$WR7__LOd#RH
sbF0OR5Nkb0sOC_D:	RRRHM#_08DHFoOO;RNkb0sCC_MRR:H#MR0D8_FOoH;E
#H_V08:sRRRHM#_08DHFoOl;RFR8C:MRHR8#0_oDFH
O;#:HRRRHM#_08DHFoO8;RN_0NH:MRRRHM#_08DHFoO8;
N_0NFRk0:kRF00R#8F_Do;HORR#F:kRF00R#8F_DoRHO2
;
-N-R0H0sLCk0RO8CDNNs0MHFRsVFRM#HoRDC#sFkO8CRCo#HMsINCR
RRRRRR0RN0LsHkR0C#_$MLDkH0_HM8:kRRs#0H;Mo
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kVRFR_7WLdO_RC:RM00H$#RHRC"IN;	"
C

M78RWO_L_
d;
ONsECH0Os0kC0RsDVRFR_7WLdO_R
H#
R--Ns00H0LkCCR8OsDNNF0HMFRVsHR#MCoDRk#FsROC8HC#oNMIs
CRNs00H0LkC$R#Mk_LHHD0Mk_8R#:R0MsHoN;
0H0sLCk0RM#$_HLkDM0H_R8kFsVR0:DRRONsECH0Os0kC#RHRC"IN;	"
-R
-FRwsHR#MCoDRk#FsROC7RW,NEsOHO0C0CksRF#EkRD8L8CRk$ll
0N0skHL0#CR$LM_D	NO_GLFRL:RFCFDN
M;Ns00H0LkC$R#MD_LN_O	LRFGFsVR0:DRRONsECH0Os0kC#RHRk0sC
;
LHCoMC

Ms8R0
D;
H
DLssN$ RQ 7 ,W q),j7Wck;
#QCR 3  #_08DHFoO4_4nNc3D
D;kR#C7)Wq W37b	NON#oC3DND;#
kCWR7j7c3W_jcObFlFMMC0N#3D
D;
0CMHR0$7LW_OR_cHb#
FRs05bON0Cks_	ODRH:RM0R#8F_Do;HO
bON0Cks_RCM:MRHR8#0_oDFH
O;#VEH0s_8RH:RM0R#8F_Do;HO
R#H:MRHR8#0_oDFH
O;8NN0_RHM:MRHR8#0_oDFH
O;#:FRR0FkR8#0_oDFH
O;8NN0_0FkRF:Rk#0R0D8_FOoHR
2;
R--Ns00H0LkCCR8OsDNNF0HMFRVsHR#MCoDRk#FsROC8HC#oNMIsRC
RRRRRNRR0H0sLCk0RM#$_HLkDM0H_R8k:0R#soHM;R
RRRRRR0RN0LsHkR0C#_$MLDkH0_HM8FkRVWR7__LOcRR:CHM00H$R#IR"C"N	;C

M78RWO_L_
c;
ONsECH0Os0kC0RsDVRFR_7WLcO_R
H#
R--Ns00H0LkCCR8OsDNNF0HMFRVsHR#MCoDRk#FsROC8HC#oNMIs
CRNs00H0LkC$R#Mk_LHHD0Mk_8R#:R0MsHoN;
0H0sLCk0RM#$_HLkDM0H_R8kFsVR0:DRRONsECH0Os0kC#RHRC"IN;	"
-R
-FRwsHR#MCoDRk#FsROC7RW,NEsOHO0C0CksRF#EkRD8L8CRk$ll
0N0skHL0#CR$LM_D	NO_GLFRL:RFCFDN
M;Ns00H0LkC$R#MD_LN_O	LRFGFsVR0:DRRONsECH0Os0kC#RHRk0sC
;
LHCoMM
C80RsD
;

LDHs$NsR Q  W,7q,) 7cWj;#
kC RQ # 30D8_FOoH_n44cD3NDk;
#7CRW q)3b7WNNO	o3C#N;DD
Ck#Rj7WcW37jOc_FFlbM0CM#D3ND
;
CHM007$RWO_L_H6R#F
bs50RO0Nbk_sCORD	:MRHR8#0_oDFHRO;kNb80OC_D:	RRRHM#_08DHFoOO;
Nkb0sCC_MRR:H#MR0D8_FOoH;bRk8CN0_RCM:MRHR8#0_oDFH
O;#VEH0s_8RH:RM0R#8F_Do;HOR8lFCRR:H#MR0D8_FOoH;M
H00C#RH:RM0R#8F_Do;HORR#H:MRHR8#0_oDFH
O;8NN0_RHM:MRHR8#0_oDFHRO;8NN0_0FkRF:Rk#0R0D8_FOoH;F
#RF:Rk#0R0D8_FOoHR
2;
R--Ns00H0LkCCR8OsDNNF0HMFRVsHR#MCoDRk#FsROC8HC#oNMIsRC
RRRRRNRR0H0sLCk0RM#$_HLkDM0H_R8k:0R#soHM;R
RRRRRR0RN0LsHkR0C#_$MLDkH0_HM8FkRVWR7__LO6RR:CHM00H$R#IR"C"N	;


CRM87LW_O;_6
s
NO0EHCkO0ssCR0FDRVWR7__LO6#RH
-
-R0N0skHL08CRCNODsHN0FVMRF#sRHDMoCFR#kCsOR#8CHIoMNRsC
0N0skHL0#CR$LM_k0HDH8M_kRR:#H0sM
o;Ns00H0LkC$R#Mk_LHHD0Mk_8RRFVsR0D:sRNO0EHCkO0sHCR#IR"C"N	;

R-w-RF#sRHDMoCFR#kCsOR,7WRONsECH0Os0kCER#F8kDRRLC8lkl$0
N0LsHkR0C#_$MLODN	F_LGRR:LDFFC;NM
0N0skHL0#CR$LM_D	NO_GLFRRFVsR0D:sRNO0EHCkO0sHCR#sR0k
C;
C
Lo
HM
8CMRDs0;D

HNLssQ$R ,  7)Wq W,7j
c;kR#CQ   38#0_oDFH4O_43ncN;DD
Ck#Rq7W)7 3WObN	CNo#D3NDk;
#7CRW3jc7cWj_lOFbCFMM30#N;DD
M
C0$H0R_7WL(O_R
H#b0FsRN5Obs0kCD_O	RR:H#MR0D8_FOoH;bRk8CN0_	ODRH:RM0R#8F_Do;HO
bON0Cks_RCM:MRHR8#0_oDFHRO;kNb80CC_MRR:H#MR0D8_FOoH;E
#H_V08:sRRRHM#_08DHFoOl;RF48CRH:RM0R#8F_Do;HO
8lFC:.RRRHM#_08DHFoO#;RHRR:H#MR0D8_FOoH;H
bMM_HbRk0:MRHR8#0_oDFHRO;O0FMs_FDFRk0:MRHR8#0_oDFH
O;Fbk0k80_NR0N:MRHR8#0_oDFHRO;HHO_M0bkRF:Rk#0R0D8_FOoH;N
80FN_k:0RR0FkR8#0_oDFHRO;#:FRR0FkR8#0_oDFH2OR;-

-0RN0LsHkR0C8DCON0sNHRFMVRFs#oHMD#CRFOksCCR8#MHoICNs
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kRR:#H0sM
o;RRRRRRRRNs00H0LkC$R#Mk_LHHD0Mk_8RRFV7LW_OR_(:MRC0$H0RRH#"NIC	
";
M
C8WR7__LO(
;
NEsOHO0C0CksRDs0RRFV7LW_OR_(H
#
-N-R0H0sLCk0RO8CDNNs0MHFRsVFRM#HoRDC#sFkO8CRCo#HMsINCNR
0H0sLCk0RM#$_HLkDM0H_R8k:0R#soHM;0
N0LsHkR0C#_$MLDkH0_HM8FkRV0RsDRR:NEsOHO0C0CksRRH#"NIC	
";R-
-RswFRM#HoRDC#sFkO7CRWN,RsHOE00COkRsC#kEFDL8RCkR8l
l$Ns00H0LkC$R#MD_LN_O	LRFG:FRLFNDCMN;
0H0sLCk0RM#$_NLDOL	_FFGRV0RsDRR:NEsOHO0C0CksRRH#0Csk;


LHCoMM
C80RsD
;

-

------------------------------------------------------------------------------------------------
H
DLssN$ RQ 7 ,W q),j7Wck;
#QCR 3  #_08DHFoO4_4nNc3D
D;kR#C7)Wq W37b	NON#oC3DND;#
kCWR7j7c3W_jcObFlFMMC0N#3D;D

0CMHR0$7UW_LL4j_O8CR
H#
MoCCOsHRL5R$#0CRH:RMo0CC:sR=;R.
RRRRRRRR	RR.6U__DFM$RR:HCM0oRCs:j=R;R
SR_CMlCF8RH:RMo0CC:sR=;Rj
RSRH0MH_8lFCRR:HCM0oRCs:j=R
RRRRRRRR
2;
sbF0RRRRO5RD:	RRRHM#_08DHFoOR;
RRRRRRRRR0s#_:MRRRHM#_08DHFoOR;
RRRRRRRRRHHM08_s_:MRRRHM#_08DHFoOR;
RRRRRRRRRHHM08_s_DPNRH:RM0R#8F_Do;HO
RRRRRRRR8RRN_0NH:MRRRHM#_08DHFoOC_POs0F50L$C4#*jR-48MFI0jFR2R;
RRRRRRRRRsCsF:sRR0FkR8#0_oDFH
O;RRRRRRRRR8RsRF:Rk#0R0D8_FOoH;R
RRRRRRRRR	E_ON:sRR0FkR8#0_oDFHPO_CFO0s$5L0-C#4FR8IFM0R;j2
RRRRRRRR8RRN_0NFRk0:kRF00R#8F_Do_HOP0COFLs5$#0C*4U-RI8FMR0Fj
2;SsRR8s_CsRR:FRk0#_08DHFoOS;
RFRO8CC_s:sRR0FkR8#0_oDFH
O;SCRRMDNLCRR:H#MR0D8_FOoH
RRRRRRRR
2;
R--Ns00H0LkCCR8OsDNNF0HMFRVsHR#MCoDRk#FsROC8HC#oNMIsRC
RRRRRNRR0H0sLCk0RM#$_HLkDM0H_R8k:0R#soHM;R
RRRRRR0RN0LsHkR0C#_$MLDkH0_HM8FkRVWR7_4ULj8L_C:ORR0CMHR0$H"#RI	CN"
;
CRM87UW_LL4j_O8C;N

sHOE00COkRsCsR0DF7VRWL_U4_jL8RCOH
#
-N-R0H0sLCk0RO8CDNNs0MHFRsVFRM#HoRDC#sFkO8CRCo#HMsINCNR
0H0sLCk0RM#$_HLkDM0H_R8k:0R#soHM;0
N0LsHkR0C#_$MLDkH0_HM8FkRV0RsDRR:NEsOHO0C0CksRRH#"NIC	
";R-
-RswFRM#HoRDC#sFkO7CRWN,RsHOE00COkRsC#kEFDL8RCkR8l
l$Ns00H0LkC$R#MD_LN_O	LRFG:FRLFNDCMN;
0H0sLCk0RM#$_NLDOL	_FFGRV0RsDRR:NEsOHO0C0CksRRH#0Csk;L

CMoH
M
C80RsD
;
-=-==============================================================================
==
H
DLssN$ RQ 7 ,W q),j7Wck;
#QCR 3  #_08DHFoO4_4nNc3D
D;kR#C7)Wq W37b	NON#oC3DND;#
kCWR7j7c3W_jcObFlFMMC0N#3D
D;
0CMHR0$7UW_LL4j_OCMR
H#
MoCCOsHRL5R$#0CRH:RMo0CC:sR=nR4;R
RRRRRRRRR	_.U6M_FD:$RR0HMCsoCRR:=jS;
RMRC_8lFCRR:HCM0oRCs:4=R;R
SRHHM0F_l8:CRR0HMCsoCRR:=4;R2
F
bsR0RRO5RD:	RRRHM#_08DHFoOR;
RRRRRRRRs_#0MRR:H#MR0D8_FOoH;R
RRRRRRHRRM_H0sM8_RH:RM0R#8F_Do;HO
RRRRRRRRMRHHs0_8N_PDRR:H#MR0D8_FOoH;R
RRRRRR	RR_NOEsRR:H#MR0D8_FOoH_OPC05FsLC$0#R-48MFI0jFR2R;
RRRRRRRR8NN0_RHM:MRHR8#0_oDFHPO_CFO0s$5L0*C#UR-48MFI0jFR2R;
RRRRRRRRs:8RR0FkR8#0_oDFH
O;RRRRRRRRR08NNk_F0RR:FRk0#_08DHFoOC_POs0F50L$C4#*jR-48MFI0jFR2S;
RNCMLRDC:MRHR8#0_oDFHRO
RRRRR2RR;-
-R0N0skHL08CRCNODsHN0FVMRF#sRHDMoCFR#kCsOR#8CHIoMN
sCRRRRRRRRNs00H0LkC$R#Mk_LHHD0Mk_8R#:R0MsHoR;
RRRRRNRR0H0sLCk0RM#$_HLkDM0H_R8kF7VRWL_U4_jLCRMO:MRC0$H0RRH#"NIC	
";
8CMR_7WUjL4LM_CO
;
NEsOHO0C0CksRDs0RRFV7UW_LL4j_OCMR
H#
R--Ns00H0LkCCR8OsDNNF0HMFRVsHR#MCoDRk#FsROC8HC#oNMIs
CRNs00H0LkC$R#Mk_LHHD0Mk_8R#:R0MsHoN;
0H0sLCk0RM#$_HLkDM0H_R8kFsVR0:DRRONsECH0Os0kC#RHRC"IN;	"
-R
-FRwsHR#MCoDRk#FsROC7RW,NEsOHO0C0CksRF#EkRD8L8CRk$ll
0N0skHL0#CR$LM_D	NO_GLFRL:RFCFDN
M;Ns00H0LkC$R#MD_LN_O	LRFGFsVR0:DRRONsECH0Os0kC#RHRk0sC
;
LHCoM


CRM8s;0D



DsHLNRs$Q   ,q7W)7 ,W;jc
Ck#R Q  03#8F_Do_HO4c4n3DND;#
kCWR7q3) 7NWbOo	NCN#3D
D;kR#C7cWj3j7WcF_OlMbFC#M03DND;C

M00H$WR7_OOs_HbR#o

CsMCH5OR8NN0_8IH0:ERRaQh )t RR:=4Rg;b$FD_x#HCRR:Q hatR ):6=R;s
OOV_OoRR:Q hatR ):(=R;HRL0s_F8RCs:hRQa  t)=R:R
j;b$FD_COFV:jRRaQh )t RR:=6b;RF_D$OVFC4RR:Q hatR ):j=R;F
bDO$_F.CVRQ:Rhta  :)R=;RjRDbF$F_OCRVd:hRQa  t)=R:R2j
;b

FRs0508NNM_HRH:RM0R#8F_Do_HOP0COF8s5N_0NI0H8ER-48MFI0jFR2O;
sHO_MRR:H#MR0D8_FOoH_OPC05Fsb$FD_x#HCR-48MFI0jFR2O;
sFO_	RR:FRk0#_08DHFoOO;
sFO_k:0RR0FkR8#0_oDFHPO_CFO0sF5bD#$_H-xC4FR8IFM0RRj22
;
-N-R0H0sLCk0RO8CDNNs0MHFRsVFRM#HoRDC#sFkO8CRCo#HMsINCR
RRRRRR0RN0LsHkR0C#_$MLDkH0_HM8:kRRs#0H;Mo
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kVRFR_7WO_sObRR:CHM00H$R#IR"C"N	;C

M78RWs_OO;_b
s
NO0EHCkO0ssCR0FDRVWR7_OOs_HbR#-

-0RN0LsHkR0C8DCON0sNHRFMVRFs#oHMD#CRFOksCCR8#MHoICNsR0
N0LsHkR0C#_$MLDkH0_HM8:kRRs#0H;Mo
0N0skHL0#CR$LM_k0HDH8M_kVRFRDs0RN:RsHOE00COkRsCH"#RI	CN"R;

R--wRFs#oHMD#CRFOksCWR7,sRNO0EHCkO0s#CREDFk8CRLRl8klN$
0H0sLCk0RM#$_NLDOL	_F:GRRFLFDMCN;0
N0LsHkR0C#_$MLODN	F_LGVRFRDs0RN:RsHOE00COkRsCH0#Rs;kC
oLCH
M
CRM8s;0D



DsHLNRs$Q   ,q7W)7 ,W;jc
Ck#R Q  03#8F_Do_HO4c4n3DND;#
kCWR7q3) 7NWbOo	NCN#3D
D;kR#C7cWj3j7WcF_OlMbFC#M03DND;C

M00H$WR7jOc_s.OdR
H#
MoCCOsHR85
N_0NI0H8EF_bIRCs:hRQa  t)=R:R
6;lCF8_D#CCRO0:hRQa  t)=R:R2d
;b

FRs05_
8H:MRRRHM#_08DHFoOC_POs0F5*.*8NN0_8IH0bE_FsIC-84RF0IMF2Rj;D
O	RR:H#MR0D8_FOoH;C
s#_C0hRR:H#MR0D8_FOoH;M
CNCLDRH:RM0R#8F_Do;HO
0L$CH_0l:CRRRHM#_08DHFoO#;
00NsRH:RM0R#8F_Do;HO
N8sH:MRRRHM#_08DHFoO8;
_0FkRF:Rk#0R0D8_FOoH_OPC05Fs.8**N_0NI0H8EF_bI-Cs4FR8IFM0R;j2
ONOkDlkNM0HoRR:FRk0#_08DHFoO8;
sMNHHRMo:kRF00R#8F_Do;HO
OOs_RF	:kRF00R#8F_Do;HO
OOs_osCRF:Rk#0R0D8_FOoH_OPC05Fsd84RF0IMF2Rj

2;-N-R0H0sLCk0RO8CDNNs0MHFRsVFRM#HoRDC#sFkO8CRCo#HMsINCR
RRRRRR0RN0LsHkR0C#_$MLDkH0_HM8:kRRs#0H;Mo
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kVRFRj7Wcs_OORd.:MRC0$H0RRH#"NIC	
";
8CMRj7Wcs_OO;d.
s
NO0EHCkO0ssCR0FDRVWR7jOc_s.OdR
H#
R--Ns00H0LkCCR8OsDNNF0HMFRVsHR#MCoDRk#FsROC8HC#oNMIs
CRNs00H0LkC$R#Mk_LHHD0Mk_8R#:R0MsHoN;
0H0sLCk0RM#$_HLkDM0H_R8kFsVR0:DRRONsECH0Os0kC#RHRC"IN;	"
-R
-FRwsHR#MCoDRk#FsROC7RW,NEsOHO0C0CksRF#EkRD8L8CRk$ll
0N0skHL0#CR$LM_D	NO_GLFRL:RFCFDN
M;Ns00H0LkC$R#MD_LN_O	LRFGFsVR0:DRRONsECH0Os0kC#RHRk0sCL;
CMoH
M
C80RsD
;

=--=========================================0CMHR0$NRM8NEsOHO0C0CksRsVFRj8IcE_#Ns8_C=oR========================
H
DLssN$ RQ 
 ;kR#CQ   38#0_oDFH4O_43ncN;DD
Ck#RCHCC03#8F_Do_HOkHM#o8MC3DND;C

M00H$WR7j#c_E_N8sRCoHo#
CsMCH
O5SHSI8S0ESRR:uQm1a QeRR:=cS;
S8LD_N#E8C_soRR:hzqa)RqpRR:=jS
S2S;
b0Fs5SR
S08NNRHMSRS:H#MR0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2S;
S##$_	ODRRS:H#MR0D8_FOoH;S
S#8EN_	ODRRS:H#MR0D8_FOoH;S
SsCC#0SRS:MRHR8#0_oDFH
O;SQS1RSSS:MRHR8#0_oDFH
O;S S1RSSS:MRHR8#0_oDFH
O;S$S##k_F0:RSR0FkR8#0_oDFHPO_CFO0sH5I8-0E4FR8IFM0R;j2
#SSE_N8FRk0SF:Rk#0R0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2S;
SR1mS:SSR0FkR8#0_oDFHSO
SS2;
-
-R0N0skHL08CRCNODsHN0FVMRF#sRHDMoCFR#kCsOR#8CHIoMN
sCRRRRRRRRNs00H0LkC$R#Mk_LHHD0Mk_8R#:R0MsHoR;
RRRRRNRR0H0sLCk0RM#$_HLkDM0H_R8kF7VRW_jc#8EN_osCRC:RM00H$#RHRC"IN;	"
M
C8WR7j#c_E_N8sRCo;N

sHOE00COkRsCsR0DF7VRW_jc#8EN_osCR#RHR-

-0RN0LsHkR0C8DCON0sNHRFMVRFs#oHMD#CRFOksCCR8#MHoICNsR0
N0LsHkR0C#_$MLDkH0_HM8:kRRs#0H;Mo
0N0skHL0#CR$LM_k0HDH8M_kVRFRDs0RN:RsHOE00COkRsCH"#RI	CN"R;

R--wRFs#oHMD#CRFOksCWR7,sRNO0EHCkO0s#CREDFk8CRLRl8klN$
0H0sLCk0RM#$_NLDOL	_F:GRRFLFDMCN;0
N0LsHkR0C#_$MLODN	F_LGVRFRDs0RN:RsHOE00COkRsCH0#Rs;kC
C
Lo
HM
8CMRDs0;


-=-=========================================CHM00N$RMN8RsHOE00COkRsCVRFs8cIj_M#$O=R======================
==DsHLNRs$HCCC,$R#MHbDV
$;kR#CHCCC38#0_oDFH4O_43ncN;DD
Ck#RM#$bVDH$03N0LsHk#0C3DND;C

M00H$WR7j#c_$RMOHo#
CsMCH5OR
MSSkNl_#O$MRRS:uQm1a QeRc:=RS;
S8sCkRM8SRS:uQm1a QeR4:=
2SS;b

F5s0
#SN$SMO:RHMR8#0_oDFHPO_CFO0sk5Ml#_N$-MO4FR8IFM0R;j2
SRRs_CVOSD	:RHMR8#0_oDFH
O;S#sCC:0SHRMR#_08DHFoOS;
CFsssFS:k#0R0D8_FOoH;#
S$SMO:0FkR8#0_oDFHPO_CFO0sk5Ml#_N$-MO4FR8IFM0R
j2S;R2
-
-R0N0skHL08CRCNODsHN0FVMRF#sRHDMoCFR#kCsOR#8CHIoMN
sCRRRRRRRRNs00H0LkC$R#Mk_LHHD0Mk_8R#:R0MsHoR;
RRRRRNRR0H0sLCk0RM#$_HLkDM0H_R8kF7VRW_jc#O$MRC:RM00H$#RHRC"IN;	"
M
C8WR7j#c_$;MO
s
NO0EHCkO0ssCR0FDRVWR7j#c_$RMOH
#
-N-R0H0sLCk0RO8CDNNs0MHFRsVFRM#HoRDC#sFkO8CRCo#HMsINCNR
0H0sLCk0RM#$_HLkDM0H_R8k:0R#soHM;0
N0LsHkR0C#_$MLDkH0_HM8FkRV0RsDRR:NEsOHO0C0CksRRH#"NIC	
";R-
-RswFRM#HoRDC#sFkO7CRWN,RsHOE00COkRsC#kEFDL8RCkR8l
l$Ns00H0LkC$R#MD_LN_O	LRFG:FRLFNDCMN;
0H0sLCk0RM#$_NLDOL	_FFGRV0RsDRR:NEsOHO0C0CksRRH#0Csk;


LHCoMC

Ms8R0
D;








