--
@ER--B$FbsEHo0OR52gR4g-cRRj.jd$R1MHbDO$H0ROQM
R--fN]C8:CsR#//$DMbH0OH$N/lb0DN.Uj4J4.b/blNb#Cs/0DN0CHO/LDH/MoC_PDNNl4/k3D0PyE84
Rf-
-

LDHs$NsR Q  k;
#QCR 3  #_08DHFoO4_4nNc3D
D;
C

M00H$zRvpHaR#
R
oCCMs5HORR
RRRRRRHRI8R0E:MRH0CCos=R:R;4dRR
RRRRRRIRNHE80RH:RMo0CC:sR=;R6RR
RRRRRRIRLHE80RH:RMo0CC:sR=RRU
RRRRRRRRRRRRRRRR2RR;
R
b0Fs5
R
RRRRRRRRqH:RM0R#8F_Do_HOP0COFNs5I0H8E4R-RI8FMR0FjR2;
RRRRRRRRRA:H#MR0D8_FOoH_OPC05FsL8IH0-ER4FR8IFM0R;j2RR
RRRRRR)Rum:7RR0FkR8#0_oDFHPO_CFO0sH5I8R0E-84RF0IMF2RjR2

;
R
CRM8vazp;
R

ONsECH0Os0kCuRpvz_vpFaRVzRvpHaR#


ObFlFMMC0uRpvz_vpRa
RCRoMHCsO5RR
RRRRRRRRRRRRRRRD_bl0C$bR#:R0MsHo=R:Rb"Dlk_lD;0"
RRRRRRRRRRRRRRRD_blI0H8E:NRR#bFHP0HCR;
RRRRRRRRRRRRRbRDlH_I8L0ERb:RF0#HH;PCRRRRRRRRR
RRRRRRRRRRRRRRRDRRbIl_HE80bRR:bHF#0CHP;RR
RRRRRRRRRRRRRbRDlH_EMR0RR#:R0MsHo=R:Ru"1 " 72R;
RFRbs
05RRRRRNR80RNNRRRRRRRRRRRRRRR:RRHMR1RRap7_mBtQ_Be a5m)D_blI0H8E4N-RI8FMR0Fj
2;RRRRRNR80RNLRRRRRRRRRRRRRRR:RRHMR1RRap7_mBtQ_Be a5m)D_blI0H8E4L-RI8FMR0Fj
2;RRRRRCRs#0kDRRRRRRRRRRRRRRR:R0FkR1RRap7_mBtQ_Be a5m)D_blI0H8E4b-RI8FMR0Fj;22
8CMRlOFbCFMM
0;
oLCH
M
RRRRR:z4p_uvvazpRMoCCOsHRblN5lDb_8IH0RENRR=>N8IH0
E,RRRRRRRRRRRRRRRRRRRRRRRRRlDb_8IH0RELRRRRRR=>L8IH0
E,RRRRRRRRRRRRRRRRRRRRRRRRRlDb_8IH0REbRRRRRR=>I0H8ER,
RRRRRRRRRRRRRRRRRRRRRRRRD_blE0HMRRRRRRRR=">R1 u 7
"2RRRRRRRRRRRRRRRRRsbF0NRlbN580RNNRRRRRRRRRR=>qR,
RRRRRRRRRRRRRRRRRRRRRRRRR08NNRLRRRRRRRRR=A>R,R
RRRRRRRRRRRRRRRRRRRRRRRRRskC#DR0RRRRRR=RR>)Rum;72
C

Mp8Ruvv_z;pa




