--*****************************************************
@Ea--HC0D:RRRR_#LH_OCObFlFMMC0##_$PM3E
8R-k-q0sEF:RRR[FoDM-o
-MwkOF0HMH:RMN#0MN0H0NCRD0DREOCRC#DDRRFV0REC#HL_O#C_$PM3RLDHs$NsR-
-BbFlN:M$RHR1DFHOMkADCCRaOFEMDHFoCR#,Q3MO
Q--h:QaRRRRRLwCR,4URj.jU-
-*****************************************************D*
HNLssH$RCRCC;#
kCCRHC#C30D8_FOoH_n44cD3ND
;
b	NONRoCBumvmhh aH1R#0
N0LsHkR0C#_$MLODN	F_LGRR:LDFFC;NM
0N0skHL0#CR$DM_HOL_CRDD:FRLFNDCMN;
0H0sLCk0R_GOlRNb:0R#soHM;0
N0LsHkR0C#_$MLODN	F_LGVRFRlOFbCFMMR0#:NRbOo	NC#RHRk0sCN;
0H0sLCk0RM#$_LDH_DOCDVRFRlOFbCFMMR0#:NRbOo	NC#RHRk0sC
;
ObFlFMMC0AR1_)Bq)
YRRRRRRRRRRFRbsR05
RRRRRRRRRRRRRRRRRBm:kRF00R#8F_DoRHORR;
RRRRRRRRRRRRRQRRjRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRRQR4:RRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRRBQ:MRHR0R#8F_DoRHO
RRRRRRRRRRRRRRR2C;
MO8RFFlbM0CM;O

FFlbM0CMR_1AB)q)Yh_Q_Xvz
RRRRRRRRoRRCsMCH5ORRQB_hRQa:HRL0C_POs0F5RR4RI8FMR0Fj22RR
R;RRRRRRRRRFRbsR05
RRRRRRRRRRRRRRRRsONsH$_M_H0FRk0:FRRk#0R0D8_FOoHRR;
RRRRRRRRRRRRRORRN$ss_HHM0M_HRRR:RRHMR8#0_oDFH
ORRRRRRRRRRRRRR2RR;M
C8FROlMbFC;M0
F
OlMbFCRM01pA_z
acRRRRRRRRRCRoMHCsORR5p_zaQahQRL:RHP0_CFO0s45R68RRF0IMF2RjR;2R
RRRRRRRRbRRF5s0RR
RRRRRRRRRRRRRRRRmRF:Rk#0R0D8_FOoHRR;
RRRRRRRRRRRRRQRRjRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRRQ:4RRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRRQ.:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRdRQRH:RM#RR0D8_FOoHRR
RRRRRRRRRRRRRR
2;CRM8ObFlFMMC0N;
0H0sLCk0R_GOlRNbF1VRAz_pa:cRRlOFbCFMMH0R#DR"k;0"
F
OlMbFCRM017A_wRw
RRRRRRRRRsbF0
5RRRRRRRRRRRRRRRRRTRR:FRk0#_08DHFoO
R;RRRRRRRRRRRRRRRRBRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRR7RR:HRMR#_08DHFoORR
RRRRRRRRRRRRR;R2
8CMRlOFbCFMM
0;
lOFbCFMM10RAw_7w
1)RRRRRRRRRFRbsR05
RRRRRRRRRRRRRRRR:TRR0FkR8#0_oDFH;OR
RRRRRRRRRRRRRRRR:BRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRR:7RRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRR:)RRRHMR8#0_oDFH
ORRRRRRRRRRRRRR2RR;M
C8FROlMbFC;M0
F
OlMbFCRM017A_w1w1
RRRRRRRRbRRF5s0RR
RRRRRRRRRRRRRRRRT:kRF00R#8F_DoRHO;R
RRRRRRRRRRRRRRRRB:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRRR7:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRRR1:MRHR0R#8F_DoRHO
RRRRRRRRRRRRRRR2C;
MO8RFFlbM0CM;O

FFlbM0CMR_1A7)ww
RRRRRRRRbRRF5s0RR
RRRRRRRRRRRRRRRRT:kRF00R#8F_DoRHO;R
RRRRRRRRRRRRRRRRB:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRRR7:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRRR):MRHR0R#8F_DoRHO
RRRRRRRRRRRRRRR2C;
MO8RFFlbM0CM;O

FFlbM0CMR_1A71ww
RRRRRRRRbRRF5s0RR
RRRRRRRRRRRRRRRRT:kRF00R#8F_DoRHO;R
RRRRRRRRRRRRRRRRB:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRRR7:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRRR1:MRHR0R#8F_DoRHO
RRRRRRRRRRRRRRR2C;
MO8RFFlbM0CM;O

FFlbM0CMR_1A7 ww
RRRRRRRRbRRF5s0RR
RRRRRRRRRRRRRRRRT:kRF00R#8F_DoRHO;R
RRRRRRRRRRRRRRRRB:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRRR :MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRRR7:MRHR0R#8F_DoRHO
RRRRRRRRRRRRRRR2C;
MO8RFFlbM0CM;O

FFlbM0CMR_1A7 ww1R)
RRRRRRRRRsbF0
5RRRRRRRRRRRRRRRRRTRR:FRk0#_08DHFoO
R;RRRRRRRRRRRRRRRRBRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRR RR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRR7RR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRR)RR:HRMR#_08DHFoORR
RRRRRRRRRRRRR;R2
8CMRlOFbCFMM
0;
lOFbCFMM10RAw_7w1 1
RRRRRRRRbRRF5s0RR
RRRRRRRRRRRRRRRRT:kRF00R#8F_DoRHO;R
RRRRRRRRRRRRRRRRB:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRRR :MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRRR7:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRRR1:MRHR0R#8F_DoRHO
RRRRRRRRRRRRRRR2C;
MO8RFFlbM0CM;O

FFlbM0CMR_1A7 ww)R
RRRRRRRRRb0Fs5RR
RRRRRRRRRRRRRTRRRF:Rk#0R0D8_FOoHRR;
RRRRRRRRRRRRRBRRRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRR RRRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRR7RRRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRR)RRRH:RM#RR0D8_FOoHRR
RRRRRRRRRRRRRR
2;CRM8ObFlFMMC0
;
ObFlFMMC0AR1_w7w R1
RRRRRRRRRsbF0
5RRRRRRRRRRRRRRRRRTRR:FRk0#_08DHFoO
R;RRRRRRRRRRRRRRRRBRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRR RR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRR7RR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRR1RR:HRMR#_08DHFoORR
RRRRRRRRRRRRR;R2
8CMRlOFbCFMM
0;
lOFbCFMM10RAw_7wRh
RRRRRRRRRsbF0
5RRRRRRRRRRRRRRRRRTRR:FRk0#_08DHFoO
R;RRRRRRRRRRRRRRRRBRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRR7RR:HRMR#_08DHFoORR
RRRRRRRRRRRRR;R2
8CMRlOFbCFMM
0;
lOFbCFMM10RAw_7w)h1
RRRRRRRRbRRF5s0RR
RRRRRRRRRRRRRRRRT:kRF00R#8F_DoRHO;R
RRRRRRRRRRRRRRRRB:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRRR7:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRRR):MRHR0R#8F_DoRHO
RRRRRRRRRRRRRRR2C;
MO8RFFlbM0CM;O

FFlbM0CMR_1A7hww1R1
RRRRRRRRRsbF0
5RRRRRRRRRRRRRRRRRTRR:FRk0#_08DHFoO
R;RRRRRRRRRRRRRRRRBRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRR7RR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRR1RR:HRMR#_08DHFoORR
RRRRRRRRRRRRR;R2
8CMRlOFbCFMM
0;
lOFbCFMM10RAw_7w
h)RRRRRRRRRFRbsR05
RRRRRRRRRRRRRRRR:TRR0FkR8#0_oDFH;OR
RRRRRRRRRRRRRRRR:BRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRR:7RRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRR:)RRRHMR8#0_oDFH
ORRRRRRRRRRRRRR2RR;M
C8FROlMbFC;M0
F
OlMbFCRM017A_w1wh
RRRRRRRRbRRF5s0RR
RRRRRRRRRRRRRRRRT:kRF00R#8F_DoRHO;R
RRRRRRRRRRRRRRRRB:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRRR7:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRRR1:MRHR0R#8F_DoRHO
RRRRRRRRRRRRRRR2C;
MO8RFFlbM0CM;O

FFlbM0CMR_1A7hww R
RRRRRRRRRb0Fs5RR
RRRRRRRRRRRRRTRRRF:Rk#0R0D8_FOoHRR;
RRRRRRRRRRRRRBRRRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRR RRRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRR7RRRH:RM#RR0D8_FOoHRR
RRRRRRRRRRRRRR
2;CRM8ObFlFMMC0
;
ObFlFMMC0AR1_w7wh) 1
RRRRRRRRbRRF5s0RR
RRRRRRRRRRRRRRRRT:kRF00R#8F_DoRHO;R
RRRRRRRRRRRRRRRRB:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRRR :MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRRR7:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRRR):MRHR0R#8F_DoRHO
RRRRRRRRRRRRRRR2C;
MO8RFFlbM0CM;O

FFlbM0CMR_1A7hww 
11RRRRRRRRRFRbsR05
RRRRRRRRRRRRRRRR:TRR0FkR8#0_oDFH;OR
RRRRRRRRRRRRRRRR:BRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRR: RRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRR:7RRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRR:1RRRHMR8#0_oDFH
ORRRRRRRRRRRRRR2RR;M
C8FROlMbFC;M0
F
OlMbFCRM017A_w wh)R
RRRRRRRRRb0Fs5RR
RRRRRRRRRRRRRTRRRF:Rk#0R0D8_FOoHRR;
RRRRRRRRRRRRRBRRRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRR RRRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRR7RRRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRR)RRRH:RM#RR0D8_FOoHRR
RRRRRRRRRRRRRR
2;CRM8ObFlFMMC0
;
ObFlFMMC0AR1_w7wh
 1RRRRRRRRRFRbsR05
RRRRRRRRRRRRRRRR:TRR0FkR8#0_oDFH;OR
RRRRRRRRRRRRRRRR:BRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRR: RRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRR:7RRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRR:1RRRHMR8#0_oDFH
ORRRRRRRRRRRRRR2RR;M
C8FROlMbFC;M0
F
OlMbFCRM01)A_qivchR)
RRRRRRRRRMoCCOsHRQ5Rh_QajRR:L_H0P0COFRs5.R66RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRRRRRQQhaR_4:HRL0C_POs0F56R.68RRF0IMF2RjR
;RRRRRRRRRRRRRRRRRRRRRQahQ_:.RR0LH_OPC05FsR6.6RFR8IFM0RRj2;RR
RRRRRRRRRRRRRRRRRQRRh_QadRR:L_H0P0COFRs5.R66RI8FMR0Fj;2RRR
RRRRRRRRRRRRRRRRRRhRQQca_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2RR;
RRRRRRRRRRRRRRRRRRRRQQhaR_6:HRL0C_POs0F56R.68RRF0IMF2RjRR;
RRRRRRRRRRRRRRRRRQRRh_QanRR:L_H0P0COFRs5.R66RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRRRRRQQhaR_(:HRL0C_POs0F56R.68RRF0IMF2RjRR;
RRRRRRRRRRRRRRRRRQRRh_QaURR:L_H0P0COFRs5.R66RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRRRRRQQhaR_g:HRL0C_POs0F56R.68RRF0IMF2RjRR;
RRRRRRRRRRRRRRRRRQRRh_QaqRR:L_H0P0COFRs5.R66RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRRRRRQQhaR_A:HRL0C_POs0F56R.68RRF0IMF2RjRR;
RRRRRRRRRRRRRRRRRQRRh_QaBRR:L_H0P0COFRs5.R66RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRRRRRQQhaR_7:HRL0C_POs0F56R.68RRF0IMF2RjRR;
RRRRRRRRRRRRRRRRRQRRh_Qa RR:L_H0P0COFRs5.R66RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRRRRRQQhaR_w:HRL0C_POs0F56R.68RRF0IMF2RjRR
RRRRRRRRRRRRRRRRR2
R;RRRRRRRRRFRbsR05
RRRRRRRRRRRRRRRRq)7a:qRR0FkR8#0_oDFHPO_CFO0s45R68RRF0IMF2RjRR;
RRRRRRRRRRRRR)RRBhpiRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRR)RRB piRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRR)RR RRRRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRR)RRq)77RH:RM#RR0D8_FOoH_OPC05FsRR(R8MFI0jFR2
R;RRRRRRRRRRRRRRRRWiBpRRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRRWiBp RR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRRWR RRRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRRW7q7)RR:HRMR#_08DHFoOC_POs0F5RR(RI8FMR0Fj;2R
RRRRRRRRRRRRRRRR1vqi:RRRRHMR8#0_oDFHPO_CFO0s45R68RRF0IMF2RjRR;
RRRRRRRRRRRRRWRR7qqaRH:RM#RR0D8_FOoH_OPC05FsRR46RI8FMR0FjR2
RRRRRRRRRRRRR;R2
8CMRlOFbCFMM
0;
lOFbCFMM10RAq_)vhciWR
RRRRRRRRRoCCMsRHO5hRQQja_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2
R;RRRRRRRRRRRRRRRRRRRRQahQ_:4RR0LH_OPC05FsR6.6RFR8IFM0RRj2;RR
RRRRRRRRRRRRRRRRRQRRh_Qa.RR:L_H0P0COFRs5.R66RI8FMR0Fj;2RRR
RRRRRRRRRRRRRRRRRRhRQQda_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2RR;
RRRRRRRRRRRRRRRRRRRRQQhaR_c:HRL0C_POs0F56R.68RRF0IMF2RjR
;RRRRRRRRRRRRRRRRRRRRRQahQ_:6RR0LH_OPC05FsR6.6RFR8IFM0RRj2;R
RRRRRRRRRRRRRRRRRRhRQQna_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2
R;RRRRRRRRRRRRRRRRRRRRQahQ_:(RR0LH_OPC05FsR6.6RFR8IFM0RRj2;R
RRRRRRRRRRRRRRRRRRhRQQUa_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2
R;RRRRRRRRRRRRRRRRRRRRQahQ_:gRR0LH_OPC05FsR6.6RFR8IFM0RRj2;R
RRRRRRRRRRRRRRRRRRhRQQqa_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2
R;RRRRRRRRRRRRRRRRRRRRQahQ_:ARR0LH_OPC05FsR6.6RFR8IFM0RRj2;R
RRRRRRRRRRRRRRRRRRhRQQBa_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2
R;RRRRRRRRRRRRRRRRRRRRQahQ_:7RR0LH_OPC05FsR6.6RFR8IFM0RRj2;R
RRRRRRRRRRRRRRRRRRhRQQ a_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2
R;RRRRRRRRRRRRRRRRRRRRQahQ_:wRR0LH_OPC05FsR6.6RFR8IFM0RRj2
RRRRRRRRRRRRRRRR2RRRR;
RRRRRRRRRsbF0
5RRRRRRRRRRRRRRRRR)a7qqRR:FRk0#_08DHFoOC_POs0F56R4RFR8IFM0RRj2;R
RRRRRRRRRRRRRRBR)pRiR:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRBR)pRi :MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRR R)RRRR:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRqR)7R7):MRHR0R#8F_Do_HOP0COFRs5(8RRF0IMF2RjRR;
RRRRRRRRRRRRRWRRBhpiRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRRWRRB piRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRRWRR RRRRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRRWRRq)77RH:RM#RR0D8_FOoH_OPC05FsRR(R8MFI0jFR2
R;RRRRRRRRRRRRRRRRviq1RRR:HRMR#_08DHFoOC_POs0F56R4RFR8IFM0RRj2;R
RRRRRRRRRRRRRR7RWqRaq:MRHR0R#8F_Do_HOP0COFRs54R6R8MFI0jFR2R
RRRRRRRRRRRRRR
2;CRM8ObFlFMMC0
;
ObFlFMMC0AR1_v)qc)ihhRW
RRRRRRRRRMoCCOsHRQ5Rh_QajRR:L_H0P0COFRs5.R66RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRRRRRQQhaR_4:HRL0C_POs0F56R.68RRF0IMF2RjR
;RRRRRRRRRRRRRRRRRRRRRQahQ_:.RR0LH_OPC05FsR6.6RFR8IFM0RRj2;RR
RRRRRRRRRRRRRRRRRQRRh_QadRR:L_H0P0COFRs5.R66RI8FMR0Fj;2RRR
RRRRRRRRRRRRRRRRRRhRQQca_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2RR;
RRRRRRRRRRRRRRRRRRRRQQhaR_6:HRL0C_POs0F56R.68RRF0IMF2RjRR;
RRRRRRRRRRRRRRRRRQRRh_QanRR:L_H0P0COFRs5.R66RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRRRRRQQhaR_(:HRL0C_POs0F56R.68RRF0IMF2RjRR;
RRRRRRRRRRRRRRRRRQRRh_QaURR:L_H0P0COFRs5.R66RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRRRRRQQhaR_g:HRL0C_POs0F56R.68RRF0IMF2RjRR;
RRRRRRRRRRRRRRRRRQRRh_QaqRR:L_H0P0COFRs5.R66RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRRRRRQQhaR_A:HRL0C_POs0F56R.68RRF0IMF2RjRR;
RRRRRRRRRRRRRRRRRQRRh_QaBRR:L_H0P0COFRs5.R66RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRRRRRQQhaR_7:HRL0C_POs0F56R.68RRF0IMF2RjRR;
RRRRRRRRRRRRRRRRRQRRh_Qa RR:L_H0P0COFRs5.R66RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRRRRRQQhaR_w:HRL0C_POs0F56R.68RRF0IMF2RjRR
RRRRRRRRRRRRRRRRR2
R;RRRRRRRRRFRbsR05
RRRRRRRRRRRRRRRRq)7a:qRR0FkR8#0_oDFHPO_CFO0s45R68RRF0IMF2RjRR;
RRRRRRRRRRRRR)RRBhpiRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRR)RRB piRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRR)RR RRRRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRR)RRq)77RH:RM#RR0D8_FOoH_OPC05FsRR(R8MFI0jFR2
R;RRRRRRRRRRRRRRRRWiBphRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRRWiBp RR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRRWR RRRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRRW7q7)RR:HRMR#_08DHFoOC_POs0F5RR(RI8FMR0Fj;2R
RRRRRRRRRRRRRRRR1vqi:RRRRHMR8#0_oDFHPO_CFO0s45R68RRF0IMF2RjRR;
RRRRRRRRRRRRRWRR7qqaRH:RM#RR0D8_FOoH_OPC05FsRR46RI8FMR0FjR2
RRRRRRRRRRRRR;R2
8CMRlOFbCFMM
0;
lOFbCFMM10RAq_)v
ciRRRRRRRRRCRoMHCsORR5QahQ_:jRR0LH_OPC05FsR6.6RFR8IFM0RRj2;R
RRRRRRRRRRRRRRRRRRhRQQ4a_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2RR;
RRRRRRRRRRRRRRRRRRRRQQhaR_.:HRL0C_POs0F56R.68RRF0IMF2RjR
;RRRRRRRRRRRRRRRRRRRRRQahQ_:dRR0LH_OPC05FsR6.6RFR8IFM0RRj2;RR
RRRRRRRRRRRRRRRRRQRRh_QacRR:L_H0P0COFRs5.R66RI8FMR0Fj;2RRR
RRRRRRRRRRRRRRRRRRhRQQ6a_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2
R;RRRRRRRRRRRRRRRRRRRRQahQ_:nRR0LH_OPC05FsR6.6RFR8IFM0RRj2;R
RRRRRRRRRRRRRRRRRRhRQQ(a_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2
R;RRRRRRRRRRRRRRRRRRRRQahQ_:URR0LH_OPC05FsR6.6RFR8IFM0RRj2;R
RRRRRRRRRRRRRRRRRRhRQQga_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2
R;RRRRRRRRRRRRRRRRRRRRQahQ_:qRR0LH_OPC05FsR6.6RFR8IFM0RRj2;R
RRRRRRRRRRRRRRRRRRhRQQAa_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2
R;RRRRRRRRRRRRRRRRRRRRQahQ_:BRR0LH_OPC05FsR6.6RFR8IFM0RRj2;R
RRRRRRRRRRRRRRRRRRhRQQ7a_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2
R;RRRRRRRRRRRRRRRRRRRRQahQ_: RR0LH_OPC05FsR6.6RFR8IFM0RRj2;R
RRRRRRRRRRRRRRRRRRhRQQwa_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2RR
RRRRRRRRRRRRRRRRR;2R
RRRRRRRRbRRF5s0RR
RRRRRRRRRRRRRR7R)qRaq:kRF00R#8F_Do_HOP0COFRs54R6R8MFI0jFR2
R;RRRRRRRRRRRRRRRR)iBpRRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRR)iBp RR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRR)R RRRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRR)7q7)RR:HRMR#_08DHFoOC_POs0F5RR(RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRpWBi:RRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRpWBi: RRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRRW R:RRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRR7Wq7:)RRRHMR8#0_oDFHPO_CFO0s(5RRFR8IFM0RRj2;R
RRRRRRRRRRRRRRqRv1RiR:MRHR0R#8F_Do_HOP0COFRs54R6R8MFI0jFR2
R;RRRRRRRRRRRRRRRRWa7qqRR:HRMR#_08DHFoOC_POs0F56R4RFR8IFM0R
j2RRRRRRRRRRRRR2RR;M
C8FROlMbFC;M0
F
OlMbFCRM01QA_mR
RRRRRRRRRoCCMsRHO5QRuhY_auR RRRR:L_H0P0COFRs568RRF0IMF2Rj;R
RRRRRRRRRRRRRRRRRRzRupupzR:RRR0LH;RR
RRRRRRRRRRRRRRRRRhRR at_)tQt :)RR0LH;RR
RRRRRRRRRRRRRRRRRQRRma_1qqh7):7RRs#0HRMo
RRRRRRRRRRRRRRRR2RRRR;
RRRRRRRRRsbF0
5RRRRRRRRRRRRRRRRRuiqBq_t uRQhRRRRR:RRRFHMk#0R0D8_FOoHRR;
RRRRRRRRRRRRRpRRq]aB_uQhzea_q pzRRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRRBBpmih_ q ApRRRRR:RRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRuQhzBa_pRiRRRRRRRRR:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRzRmaauz_iBpRRRRRRRRRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRRmRRzzauah_ q ApRRRRRRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRR7z_maR_4RRRRRRRRR:RRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRm7_zja_RRRRRRRRRRRR:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRR_R7Q4h_RRRRRRRRRRRRRF:Rk#0R0D8_FOoHRR;
RRRRRRRRRRRRR7RR__QhjRRRRRRRRRRRRRR:FRk0#_08DHFoORRRRRRRRRRRRRRRRRR
RRRRRRRRRRRRR;R2
8CMRlOFbCFMM
0;
lOFbCFMM10RAA_t_
QmRRRRRRRRRCRoMHCsORR5u_Qha YuRRRR:HRL0C_POs0F5RR6RI8FMR0Fj
2;RRRRRRRRRRRRRRRRRRRRupzpzRuRRL:RHR0;
RRRRRRRRRRRRRRRRRRRRth _Qa)t)t RL:RHR0;
RRRRRRRRRRRRRRRRRRRR_Qm1haq77q)R#:R0MsHoRR
RRRRRRRRRRRRRRRRR;2R
RRRRRRRRbRRF5s0RR
RRRRRRRRRRRRRRqRuBtiq Q_uhRRRRRRRR:RRRFHMk#0R0D8_FOoHRR;
RRRRRRRRRRRRRpRRq]aB_uQhzea_q pzRRRR:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRpRBm_Bi AhqpR RRRRRR:RRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRuQhzBa_pRiRRRRRRRRRRRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRRmuzazBa_pRiRRRRRRRRRRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRRmRRzzauah_ q ApRRRRRRRR:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRR_R7m_za4RRRRRRRRRRRR:RRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRm7_zja_RRRRRRRRRRRRRRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRR7h_Q_R4RRRRRRRRRRRRRRF:Rk#0R0D8_FOoHRR;
RRRRRRRRRRRRR7RR__QhjRRRRRRRRRRRRRRR:kRF00R#8F_DoRHO;R
RRRRRRRRRRRRRRpRtmpAq_wAzw_ )muzaz:aRR0FkR8#0_oDFHRORRRRRRRRRRRRRRRR
RRRRRRRRRRRRR;R2
8CMRlOFbCFMM
0;
lOFbCFMM10RAm_Q_
71RRRRRRRRRCRoMHCsORR5u_Qha YuRRRR:HRL0C_POs0F5RR6RI8FMR0Fj
2;RRRRRRRRRRRRRRRRRRRRh_ tat)QtR ):HRL0
;RRRRRRRRRRRRRRRRRRRRRQ1m_a7qhqR)7:0R#soHMRR
RRRRRRRRRRRRRRRRR2
R;RRRRRRRRRFRbsR05
RRRRRRRRRRRRRRRRBuqi qt_huQRRRRRRRR:MRHFRk0#_08DHFoO
R;RRRRRRRRRRRRRRRRuiqBq_t u_QhARRRR:RRRFHMk#0R0D8_FOoHRR;
RRRRRRRRRRRRRpRRq]aB_uQhzea_q pzRRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRRBBpmih_ q ApRRRRR:RRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRuQhzBa_pRiRRRRRRRRR:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRzRmaauz_iBpRRRRRRRRRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRRmRRzzauah_ q ApRRRRRRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRR7z_maR_4RRRRRRRRR:RRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRm7_zja_RRRRRRRRRRRR:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRR_R7Q4h_RRRRRRRRRRRRRF:Rk#0R0D8_FOoHRR;
RRRRRRRRRRRRR7RR__QhjRRRRRRRRRRRRRR:FRk0#_08DHFoORRRRRRRRRRRRRRRRRR
RRRRRRRRRRRRR;R2
8CMRlOFbCFMM
0;
lOFbCFMM10RAA_t
RRRRRRRRbRRF5s0RR
RRRRRRRRRRRRRRpRtmpAq_wAzw_ )muzazRaRRRRRR:RRR0FkR8#0_oDFH;OR
RRRRRRRRRRRRRRRR z1)Q_1tphq__amtApmqAp_z ww)RR:HRMR#_08DHFoORR
RRRRRRRRRRRRR;R2
8CMRlOFbCFMM
0;
lOFbCFMM#0RLD_bDF_Os
CRRCRoMHCsO
R5S Sw q7ABui_qRa]S:SSRs#0HRMoRR:="v1Qu"p ;S
S7q pY7_qKaz1va h_7vm SRS:0R#soHMR=R:R$"8MHNlOR";
wSSQ7X _p7 qqY_71Kzahv aSRS:MRH0CCos=R:RRj;
uSSpzpma]_uqS1 SRS:#H0sMRoR:"=RMCFM"S;
Se7Q)SSSSL:RHP0_CFO0sR5d8MFI0jFR2=R:Rj"jj;j"
7SSQSewS:SSR0LH_OPC05Fs6FR8IFM0RRj2:"=Rjjjjj;j"
7SSQSeTS:SSR0LH_OPC05Fs.FR8IFM0RRj2:"=Rj"jj;S
SwaQp ))_q htS:SSR0LH_OPC05Fs.FR8IFM0RRj2:"=Rj"jj;SR
Sq hA_p QtB qRa S:SSR0LHRR:=';j'
aSS _1av m7RSSS:HRL0=R:R''j;S
S  Xa)phq_e7QQ_7 waqBmS)RSH:RMo0CC:sR=RR4
RRRRRRR2R;
RsbF0RR5
RRRRRRRRw)  h) Bp Bi:SSRRHM#_08DHFoOR;
RRRRRuRRpzpma)Bm :SSR0FkR8#0_oDFH
O;RRRRRRRRumppzpatmpAqSRS:FRk0#_08DHFoOR;
RRRRR RRX aw q7ABSiS:MRHR8#0_oDFH
O;Sh7YqBvQ7q pY:SSRRHM#_08DHFoOC_POs0FRR5d8MFI0jFR2
R;RRRRRRRRAqYu1S1SSH:RM0R#8F_Do;HO
RRRRRRRR1)  SaSSH:RM0R#8F_Do;HO
RRRRRRRRBpmiSSS:kRF00R#8F_Do;HO
RRRRRRRRapqBh]Quezaq pzSRS:H#MR0D8_FOoH;1
S7SmSSF:Rk#0R0D8_FOoH;1
S7SQSSH:RM0R#8F_Do;HO
BS1pSiSSH:RM0R#8F_Do
HORRRRR2RR;M
C8FROlMbFC;M0
F
OlMbFCRM0#bL_DbD_NR8
RMoCCOsHRS5
S w 7BAqiq_uaS]RSRS:#H0sMRoR:"=R1uQvp; "
7SS Ypq_Kq7zv1a _hav m7R:SSRs#0HRMoRR:="h7YqBvQ"
;RSQSwX_ 77q pY7_qKaz1va hR:SSR0HMCsoCRR:=j
;RSpSupamz_qu]1S SS#:R0MsHo:RR=MR"F"MC;S
S7)QeSSSS:HRL0C_POs0F58dRF0IMF2RjRR:="jjjj
";SQS7eSwSSRS:L_H0P0COF6s5RI8FMR0Fj:2R=jR"jjjjj
";SQS7eSTSSRS:L_H0P0COF.s5RI8FMR0Fj:2R=jR"j;j"
wSSQ pa)q_)hSt SRS:L_H0P0COF.s5RI8FMR0Fj:2R=jR"j;j"RSR
Sq hA_p QtB qRa S:SSR0LHRR:=';j'
aSS _1av m7RSSS:HRL0=R:R''j;S
S  Xa)phq_e7QQ_7 waqBmS)RSH:RMo0CC:sR=RR4
RRRRRRR2R;
RsbF0RR5
RRRRRRRRBuqi qtuSQhSH:RM0FkR8#0_oDFH
O;RRRRRRRRumppzmaB)S S:kRF00R#8F_Do;HO
RRRRRRRRpupmtzapqmAp:SSR0FkR8#0_oDFH
O;RRRRRRRR wXa A 7qSBiSH:RM0R#8F_Do;HO
SRR7qYhv7QB YpqSRS:H#MR0D8_FOoH_OPC0RFs58dRF0IMF2RjRR;
RRRRRARRY1uq1SSS:MRHR8#0_oDFH
O;RRRRRRRR)  1aSSS:MRHR8#0_oDFH
O;RRRRRRRRpimBS:SSR0FkR8#0_oDFH
O;RRRRRRRRpBqa]uQhzqaepSz SH:RM0R#8F_Do;HO
1RS7SmSSF:Rk#0R0D8_FOoH;1
S7SQSSH:RM0R#8F_Do;HO
BS1pSiSSH:RM0R#8F_Do
HOS
2;CRM8ObFlFMMC0
;
ObFlFMMC0LR#_DbD_b._N
8RRCRoMHCsO
R5S Sw q7ABui_qRa]S:SSRs#0HRMoRR:="v1Qu"p ;S
S7q pY7_qKaz1va h_7vm SRS:0R#soHMR=R:R$"8MHNlOR";
wSSQ7X _p7 qqY_71Kzahv aSRS:MRH0CCos=R:RRj;
uSSpzpma]_uqS1 SRS:#H0sMRoR:"=RMCFM"S;
Se7Q)SSSSL:RHP0_CFO0sR5d8MFI0jFR2=R:Rj"jj;j"
7SSQSewS:SSR0LH_OPC05Fs6FR8IFM0RRj2:"=Rjjjjj;j"
7SSQSeTS:SSR0LH_OPC05Fs.FR8IFM0RRj2:"=Rj"jj;S
SwaQp ))_q htS:SSR0LH_OPC05Fs.FR8IFM0RRj2:"=Rj"jj;S
S AhqpQ _Bq tau _mq)aSRS:LRH0:'=Rj
';ShS q Ap_ QBt qa_)umaSAS:HRL0=R:R''j;S
Saa 1_7vm SRSSL:RH:0R=jR''S;
Sa X q)hpQ_7e Q7_BwqaRm)SRS:HCM0oRCs:4=RRR
RRRRRR;R2
bRRFRs05RR
RRRRRuRRqqBitQ uh:SSRFHMk#0R0D8_FOoH;R
RRRRRRpRupamzB m)q:SSR0FkR8#0_oDFH
O;RRRRRRRRumppzpatmpAqq:SSR0FkR8#0_oDFH
O;RRRRRRRRumppzmaB)S ASF:Rk#0R0D8_FOoH;R
RRRRRRpRupamztApmqSpASF:Rk#0R0D8_FOoH;R
RRRRRRXR a w 7BAqi:SSRRHM#_08DHFoOS;
7qYhv7QB YpqSRS:H#MR0D8_FOoH_OPC0RFs58dRF0IMF2RjRR;
RRRRRARRY1uq1SSS:MRHR8#0_oDFH
O;RRRRRRRR)  1aSSS:MRHR8#0_oDFH
O;RRRRRRRRpimBS:SSR0FkR8#0_oDFH
O;RRRRRRRRpBqa]uQhzqaepSz SH:RM0R#8F_Do;HO
SRR1S7mSRS:FRk0#_08DHFoOS;
1S7QSRS:H#MR0D8_FOoH;1
SBSpiSRS:H#MR0D8_FOoH
RRRRRRR2R;
RM
C8FROlMbFC;M0
0
N0LsHkR0C#_$MLODN	F_LGVRFRDNDRO:RFFlbM0CMRRH#0Csk;0
N0LsHkR0C#_$MD_HLODCDRRFVNRDD:FROlMbFCRM0H0#Rs;kC
8CMRvBmu mhh;a1




