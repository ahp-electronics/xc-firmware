--*****************************************************
@Ea--HC0D:RRRR_#LH_OCObFlFMMC0D#_OE3P8-R
-#7CH:oMR#RRLO_HCF_OlMbFC#M0_3DOPRE8
q--kF0EsR:RRD[oF
Mo-k-wMHO0FRM:BbFlFMMC0F#RVER0CERb$O#HNpDRFOoHRDBCD-
-BbFlN:M$RHR1DFHOMkADCCRaOFEMDHFoCR#,Q3MO
Q--h:QaRRRRRLwCR,4URj.jU-
-*****************************************************D*
HNLssH$RCRCC;#
kCCRHC#C30D8_FOoH_n44cD3ND
;
b	NONRoC#HL_OjCc_lOFbCFMM_0#DHOR#O

FFlbM0CMR7th
RRRRRRRRbRRF5s0RR
RRRRRRRRRRRRRRRRY:kRF0#RR0D8_FOoHRR
RRRRRRRRRRRRRR;R2
8CMRlOFbCFMM
0;
lOFbCFMMe0RBRB
RRRRRRRRRsbF0
5RRRRRRRRRRRRRRRRRYRR:FRk0R8#0_oDFH
ORRRRRRRRRRRRRRRRR2C;
MO8RFFlbM0CM;


ObFlFMMC0FRDo_HOODCD
RRRRRRRRbRRF5s0
RRRRRRRRRRRRsONsF$_k:0RR0FkR8#0_oDFH
O;RRRRRRRRRRRRDFO_kR0RRRR:FRk0#_08DHFoOR;
RRRRR
RRRRRRRRRRRRRROsNs$M_HRR:RH#MR0D8_FOoH;R
RRRRRRRRRRDRO	RRRR:RRRMRHR8#0_oDFH
O;RRRRRRRRRRRROLD	RRRRRR:RH#MR0D8_FOoH;R
RRRRRRRRRRMRHjRRRR:RRRMRHR8#0_oDFH
O;RRRRRRRRRRRRHRM4RRRRRR:RH#MR0D8_FOoH;R
RRRRRRRRRRMRH.RRRR:RRRMRHR8#0_oDFH
O;RRRRRRRRRRRRHRMdRRRRRR:RH#MR0D8_FOoH;R
RRRRRRRRRRsRbFRoRR:RRRMRHR8#0_oDFH
O;RRRRRRRRRRRRb#ks0RRRRR:RH#MR0D8_FOoH;R
RRRRRRRRRR_R#sRRRR:RRRMRHR8#0_oDFH
O;RRRRRRRRRRRRO0LHRRRRRR:RH#MR0D8_FOoH_OPC05Fs.8jRF0IMF2Rj
RRRRRRRRRRRR
2;CRM8ObFlFMMC0
;
ObFlFMMC0FRpoBHOC
DDRRRRRRRRRCRoMHCsORR5
RRRRRRRRSRRSSSS1_ Tv m7RRR:L_H0P0COFds5RI8FMR0Fj:2R=jR"j"jj;R
RRRRRRRRRRSRSS_SBmRhRRRRR:HRL0=R:R''j;RR
RRRRRRRRRSRRSpSSzQa_hRQaRL:RHP0_CFO0s654RI8FMR0Fj:2R="RXjjjj"R
RRRRRRRRRRRRRRRRR2
R;RRRRRRRRRFRbsR05
RRRRRRRRRRRRRRRRsONsF$_k:0RR0FkR0R#8F_DoRHO;R
RRRRRRRRRRRRRRORD_0FkRRRR:kRF0#RR0D8_FOoHR
;
RRRRRRRRRRRRRRRROsNs$M_HRRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRRORD	RRRRRRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRROLD	RRRRRRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRRHRMjRRRRRRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRRHRM4RRRRRRR:HRMR#_08DHFoORR;
RRRRRRRRRRRRRRRR.HMRRRRR:RRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRdHMRRRRR:RRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRs#_RRRRR:RRRRHMR8#0_oDFH
ORRRRRRRRRRRRRRRRR2C;
MO8RFFlbM0CM;O

FFlbM0CMReQh
RRRRRRRRbRRF5s0RR
RRRRRRRRRRRRRRRRQRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRRmRRRF:RkR0R#_08DHFoORR
RRRRRRRRRRRRR2RR;M
C8FROlMbFC;M0
F
OlMbFCRM0H_MPE
P0RRRRRRRRRFRbsR05
RRRRRRRRRRRRRRRRRQR:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRRRm:kRF0#RR0D8_FOoHRR
RRRRRRRRRRRRRR;R2
8CMRlOFbCFMM
0;
lOFbCFMMO0RF8sCV
VsRRRRRRRRRFRbs
05RRRRRRRRRRRRJRRRRRRR:kRF00R#8F_Do;HO
RRRRRRRRR
RRRRRRRRRRRR8RRRRRRR:H#MR0D8_FOoH;R
RRRRRRRRRRkRbsR#0RRR:H#MR0D8_FOoH;R
RRRRRRRRRR_R1)RRRRRR:H#MR0D8_FOoH;R
RRRRRRRRRRDRO	RRRRRR:H#MR0D8_FOoH;R
RRRRRRRRRRDRO	RLRRRR:H#MR0D8_FOoH;R
RRRRRRRRRRLROHR0RRRR:H#MR0D8_FOoH_OPC05Fs4FR8IFM0R
j2RRRRRRRRRRRR2C;
MO8RFFlbM0CM;O

FFlbM0CMRkOD0Rc
RRRRRRRRRsbF0R5
RRRRRRRRRDRRkR0c:kRF00R#8F_Do;HO
RRRRRRRRR
RRRRRRRRRRMRHj:RRRRHM#_08DHFoOR;
RRRRRRRRRHRRMR4R:MRHR8#0_oDFH
O;RRRRRRRRRRRRHRM.RH:RM0R#8F_Do;HO
RRRRRRRRRRRRdHMRRR:H#MR0D8_FOoH;R
RRRRRRRRRRMRHj:LRRRHM#_08DHFoOR;
RRRRRRRRRHRRMR4L:MRHR8#0_oDFH
O;RRRRRRRRRRRRHLM.RH:RM0R#8F_Do;HO
RRRRRRRRRRRRdHMLRR:H#MR0D8_FOoH;R
RRRRRRRRRRLROH:0RRRHM#_08DHFoOC_POs0F5R468MFI0jFR2R
RRRRRRRRRR;R2
8CMRlOFbCFMM
0;
lOFbCFMMO0RN$ss_oDFHRO
RRRRRRRRRsbF0R5
RRRRRRRRRORRFRk0:kRF00R#8F_Do;HO
RRRRRRRRR
RRRRRRRRRRNROs_s$HRMR:MRHR8#0_oDFH
O;RRRRRRRRRRRRNRRRRRRRRRR:H#MR0D8_FOoH;R
RRRRRRRRRR_RNLRNsRRRR:MRHR8#0_oDFH
O;RRRRRRRRRRRRLRRRRRRRRRR:H#MR0D8_FOoH;R
RRRRRRRRRR_RLLRNsRRRR:MRHR8#0_oDFH
O;RRRRRRRRRRRRPCo_MRRRRRR:H#MR0D8_FOoH
RRRRRRRRRRRR
2;CRM8ObFlFMMC0
;
ObFlFMMC0_RFl
kGRRRRRRRRRFRbs
05RRRRRRRRRRRRmRRRRF:Rk#0R0D8_FOoH;R
RRRRRRRR
RRRRRRRRRHRRMRjR:MRHR8#0_oDFH
O;RRRRRRRRRRRRHRM4RH:RM0R#8F_Do;HO
RRRRRRRRRRRRHOL0RR:H#MR0D8_FOoH;R
RRRRRRRRRRsRbF:oRRRHM#_08DHFoOR
RRRRRRRRRR;R2
8CMRlOFbCFMM
0;
lOFbCFMMq0Rh
7.RRRRRRRRRFRbsR05
RRRRRRRRRRRRRRRRRqR:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRRRARH:RM#RR0D8_FOoHR
;
RRRRRRRRRRRRRRRRm:RRR0FkR0R#8F_DoRHO
RRRRRRRRRRRRRRRR
2;CRM8ObFlFMMC0
;
ObFlFMMC0DRB	Gvk
RRRRRRRRbRRF5s0RR
RRRRRRRRRRRRRRRRQRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRRmRRRRR:FRk0R8#0_oDFH
ORRRRRRRRRRRRRRRRR2C;
MO8RFFlbM0CM;O

FFlbM0CMRv1)kRG
RRRRRRRRRsbF0
5RRRRRRRRRRRRRRRRRQ:RRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRRmR:kRF0#RR0D8_FOoHRR
RRRRRRRRRRRRRR;R2
8CMRlOFbCFMM
0;
lOFbCFMMt0RDpL.FDONv
kGRRRRRRRRRFRbsR05
RRRRRRRRRRRRRRRRRQR:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRRRmRF:RkR0R#_08DHFoORR
RRRRRRRRRRRRR2RR;M
C8FROlMbFC;M0
F
OlMbFCRM0Bk vGR
RRRRRRRRRb0Fs5RR
RRRRRRRRRRRRRQRRRRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRRm:RRR0FkR0R#8F_DoRHO
RRRRRRRRRRRRRRRR
2;CRM8ObFlFMMC0
;
ObFlFMMC0bR1N.M4v
kGRRRRRRRRRFRbsR05
RRRRRRRRRRRRRRRRRQR:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRRRmRF:RkR0R#_08DHFoORR
RRRRRRRRRRRRR2RR;M
C8FROlMbFC;M0
F
OlMbFCRM01.b40
FcRRRRRRRRRFRbsR05
RRRRRRRRRRRRRRRRRQR:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRRRmRF:RkR0R#_08DHFoORR
RRRRRRRRRRRRR2RR;M
C8FROlMbFC;M0
F
OlMbFCRM0mP8scR
RRRRRRRRRb0Fs5RR
RRRRRRRRRRRRRQRRRRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRRm:RRR0FkR0R#8F_DoRHO
RRRRRRRRRRRRRRRR
2;CRM8ObFlFMMC0
;
ObFlFMMC08Rms.P4
RRRRRRRRbRRF5s0RR
RRRRRRRRRRRRRRRRQRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRRmRRRRR:FRk0R8#0_oDFH
ORRRRRRRRRRRRRRRRR2C;
MO8RFFlbM0CM;O

FFlbM0CMROpFNkDvGR
RRRRRRRRRb0Fs5RR
RRRRRRRRRRRRRQRRRRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRRm:RRR0FkR0R#8F_DoRHO
RRRRRRRRRRRRRRRR
2;CRM8ObFlFMMC0
;
ObFlFMMC0bR1NvMckRG
RRRRRRRRRsbF0
5RRRRRRRRRRRRRRRRRQ:RRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRRmR:kRF0#RR0D8_FOoHRR
RRRRRRRRRRRRRR;R2
8CMRlOFbCFMM
0;
lOFbCFMMQ0RMGvk
RRRRRRRRbRRF5s0RR
RRRRRRRRRRRRRRRRQRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRRmRRRRR:FRk0R8#0_oDFH
ORRRRRRRRRRRRRRRRR2C;
MO8RFFlbM0CM;O

FFlbM0CMRQQFMGvk
RRRRRRRRbRRF5s0RR
RRRRRRRRRRRRRRRRQRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRRmRRRRR:FRk0R8#0_oDFH
ORRRRRRRRRRRRRRRRR2C;
MO8RFFlbM0CM;O

FFlbM0CMRFoH.sB0DVAk
RRRRRRRRbRRF5s0RR
RRRRRRRRRRRRRRRRQRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRRmRRRRR:FRk0R8#0_oDFH
ORRRRRRRRRRRRRRRRR2C;
MO8RFFlbM0CM;O

FFlbM0CMRFtDLvNDk
GRRRRRRRRRRFRbsR05
RRRRRRRRRRRRRRRRRQR:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRRRmRF:RkR0R#_08DHFoORR
RRRRRRRRRRRRR2RR;M
C8FROlMbFC;M0
F
OlMbFCRM0QbF1NvMck
GRRRRRRRRRRFRbsR05
RRRRRRRRRRRRRRRRRQR:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRRRmRF:RkR0R#_08DHFoORR
RRRRRRRRRRRRR2RR;M
C8FROlMbFC;M0
F
OlMbFCRM01MbNcGvk_
PRRRRRRRRRRFRbsR05
RRRRRRRRRRRRRRRRRQR:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRRRmRF:RkR0R#_08DHFoORR
RRRRRRRRRRRRR2RR;M
C8FROlMbFC;M0
F
OlMbFCRM01MbNcGvk__#jPRR
RRRRRRRRRsbF0
5RRRRRRRRRRRRRRRRRQ:RRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRRmR:kRF0#RR0D8_FOoHRR
RRRRRRRRRRRRRR;R2
8CMRlOFbCFMM
0;
lOFbCFMM10RbcNMv_kG#P4_RR
RRRRRRRRRb0Fs5RR
RRRRRRRRRRRRRQRRRRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRRm:RRR0FkR0R#8F_DoRHO
RRRRRRRRRRRRRRRR
2;CRM8ObFlFMMC0
;
ObFlFMMC0bR1NvMck#G_.R_P
RRRRRRRRbRRF5s0RR
RRRRRRRRRRRRRRRRQRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRRmRRRRR:FRk0R8#0_oDFH
ORRRRRRRRRRRRRRRRR2C;
MO8RFFlbM0CM;O

FFlbM0CMRN1bMkcvGd_#_
PRRRRRRRRRRFRbsR05
RRRRRRRRRRRRRRRRRQR:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRRRmRF:RkR0R#_08DHFoORR
RRRRRRRRRRRRR2RR;M
C8FROlMbFC;M0
F
OlMbFCRM01MbNcGvk_
ERRRRRRRRRRFRbsR05
RRRRRRRRRRRRRRRRRQR:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRRRmRF:RkR0R#_08DHFoORR
RRRRRRRRRRRRR2RR;M
C8FROlMbFC;M0
F
OlMbFCRM01MbNcGvk__#jERR
RRRRRRRRRsbF0
5RRRRRRRRRRRRRRRRRQ:RRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRRmR:kRF0#RR0D8_FOoHRR
RRRRRRRRRRRRRR;R2
8CMRlOFbCFMM
0;
lOFbCFMM10RbcNMv_kG#E4_RR
RRRRRRRRRb0Fs5RR
RRRRRRRRRRRRRQRRRRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRRm:RRR0FkR0R#8F_DoRHO
RRRRRRRRRRRRRRRR
2;CRM8ObFlFMMC0
;
ObFlFMMC0bR1NvMck#G_.R_E
RRRRRRRRbRRF5s0RR
RRRRRRRRRRRRRRRRQRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRRmRRRRR:FRk0R8#0_oDFH
ORRRRRRRRRRRRRRRRR2C;
MO8RFFlbM0CM;O

FFlbM0CMRN1bMkcvGd_#_
ERRRRRRRRRRFRbsR05
RRRRRRRRRRRRRRRRRQR:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRRRmRF:RkR0R#_08DHFoORR
RRRRRRRRRRRRR2RR;M
C8FROlMbFC;M0
F
OlMbFCRM01MbN4k.vGR_E
RRRRRRRRbRRF5s0RR
RRRRRRRRRRRRRRRRQRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRRmRRRRR:FRk0R8#0_oDFH
ORRRRRRRRRRRRRRRRR2C;
MO8RFFlbM0CM;O

FFlbM0CMRN1bMv4.k#G_jR_E
RRRRRRRRbRRF5s0RR
RRRRRRRRRRRRRRRRQRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRRmRRRRR:FRk0R8#0_oDFH
ORRRRRRRRRRRRRRRRR2C;
MO8RFFlbM0CM;O

FFlbM0CMRN1bMv4.k#G_4R_E
RRRRRRRRbRRF5s0RR
RRRRRRRRRRRRRRRRQRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRRmRRRRR:FRk0R8#0_oDFH
ORRRRRRRRRRRRRRRRR2C;
MO8RFFlbM0CM;O

FFlbM0CMRN1bMv4.k#G_.R_E
RRRRRRRRbRRF5s0RR
RRRRRRRRRRRRRRRRQRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRRmRRRRR:FRk0R8#0_oDFH
ORRRRRRRRRRRRRRRRR2C;
MO8RFFlbM0CM;O

FFlbM0CMRN1bMv4.k#G_dR_E
RRRRRRRRbRRF5s0RR
RRRRRRRRRRRRRRRRQRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRRmRRRRR:FRk0R8#0_oDFH
ORRRRRRRRRRRRRRRRR2C;
MO8RFFlbM0CM;O

FFlbM0CMRN1bMv4.k#G_cR_E
RRRRRRRRbRRF5s0RR
RRRRRRRRRRRRRRRRQRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRRmRRRRR:FRk0R8#0_oDFH
ORRRRRRRRRRRRRRRRR2C;
MO8RFFlbM0CM;O

FFlbM0CMRN1bMv4.k#G_6R_E
RRRRRRRRbRRF5s0RR
RRRRRRRRRRRRRRRRQRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRRmRRRRR:FRk0R8#0_oDFH
ORRRRRRRRRRRRRRRRR2C;
MO8RFFlbM0CM;O

FFlbM0CMRN1bMv4.k#G_nR_E
RRRRRRRRbRRF5s0RR
RRRRRRRRRRRRRRRRQRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRRmRRRRR:FRk0R8#0_oDFH
ORRRRRRRRRRRRRRRRR2C;
MO8RFFlbM0CM;O

FFlbM0CMRN1bMv4.k#G_(R_E
RRRRRRRRbRRF5s0RR
RRRRRRRRRRRRRRRRQRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRRmRRRRR:FRk0R8#0_oDFH
ORRRRRRRRRRRRRRRRR2C;
MO8RFFlbM0CM;O

FFlbM0CMRN1bMv4.k#G_UR_E
RRRRRRRRbRRF5s0RR
RRRRRRRRRRRRRRRRQRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRRmRRRRR:FRk0R8#0_oDFH
ORRRRRRRRRRRRRRRRR2C;
MO8RFFlbM0CM;O

FFlbM0CMRN1bMv4.k#G_gR_E
RRRRRRRRbRRF5s0RR
RRRRRRRRRRRRRRRRQRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRRmRRRRR:FRk0R8#0_oDFH
ORRRRRRRRRRRRRRRRR2C;
MO8RFFlbM0CM;O

FFlbM0CMRN1bMv4.k#G_4Ej_RR
RRRRRRRRRb0Fs5RR
RRRRRRRRRRRRRQRRRRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRRm:RRR0FkR0R#8F_DoRHO
RRRRRRRRRRRRRRRR
2;CRM8ObFlFMMC0
;
ObFlFMMC0bR1N.M4v_kG#_44ERR
RRRRRRRRRsbF0
5RRRRRRRRRRRRRRRRRQ:RRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRRmR:kRF0#RR0D8_FOoHRR
RRRRRRRRRRRRRR;R2
8CMRlOFbCFMM
0;
lOFbCFMM10Rb4NM.Gvk_
PRRRRRRRRRRFRbsR05
RRRRRRRRRRRRRRRRRQR:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRRRmRF:RkR0R#_08DHFoORR
RRRRRRRRRRRRR2RR;M
C8FROlMbFC;M0
F
OlMbFCRM01MbN4k.vGj_#_
PRRRRRRRRRRFRbsR05
RRRRRRRRRRRRRRRRRQR:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRRRmRF:RkR0R#_08DHFoORR
RRRRRRRRRRRRR2RR;M
C8FROlMbFC;M0
F
OlMbFCRM01MbN4k.vG4_#_
PRRRRRRRRRRFRbsR05
RRRRRRRRRRRRRRRRRQR:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRRRmRF:RkR0R#_08DHFoORR
RRRRRRRRRRRRR2RR;M
C8FROlMbFC;M0
F
OlMbFCRM01MbN4k.vG._#_
PRRRRRRRRRRFRbsR05
RRRRRRRRRRRRRRRRRQR:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRRRmRF:RkR0R#_08DHFoORR
RRRRRRRRRRRRR2RR;M
C8FROlMbFC;M0
F
OlMbFCRM01MbN4k.vGd_#_
PRRRRRRRRRRFRbsR05
RRRRRRRRRRRRRRRRRQR:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRRRmRF:RkR0R#_08DHFoORR
RRRRRRRRRRRRR2RR;M
C8FROlMbFC;M0
F
OlMbFCRM01MbN4k.vGc_#_
PRRRRRRRRRRFRbsR05
RRRRRRRRRRRRRRRRRQR:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRRRmRF:RkR0R#_08DHFoORR
RRRRRRRRRRRRR2RR;M
C8FROlMbFC;M0
F
OlMbFCRM01MbN4k.vG6_#_
PRRRRRRRRRRFRbsR05
RRRRRRRRRRRRRRRRRQR:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRRRmRF:RkR0R#_08DHFoORR
RRRRRRRRRRRRR2RR;M
C8FROlMbFC;M0
F
OlMbFCRM01MbN4k.vGn_#_
PRRRRRRRRRRFRbsR05
RRRRRRRRRRRRRRRRRQR:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRRRmRF:RkR0R#_08DHFoORR
RRRRRRRRRRRRR2RR;M
C8FROlMbFC;M0
F
OlMbFCRM01MbN4k.vG(_#_
PRRRRRRRRRRFRbsR05
RRRRRRRRRRRRRRRRRQR:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRRRmRF:RkR0R#_08DHFoORR
RRRRRRRRRRRRR2RR;M
C8FROlMbFC;M0
F
OlMbFCRM01MbN4k.vGU_#_
PRRRRRRRRRRFRbsR05
RRRRRRRRRRRRRRRRRQR:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRRRmRF:RkR0R#_08DHFoORR
RRRRRRRRRRRRR2RR;M
C8FROlMbFC;M0
F
OlMbFCRM01MbN4k.vGg_#_
PRRRRRRRRRRFRbsR05
RRRRRRRRRRRRRRRRRQR:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRRRmRF:RkR0R#_08DHFoORR
RRRRRRRRRRRRR2RR;M
C8FROlMbFC;M0
F
OlMbFCRM01MbN4k.vG4_#jR_P
RRRRRRRRbRRF5s0RR
RRRRRRRRRRRRRRRRQRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRRmRRRRR:FRk0R8#0_oDFH
ORRRRRRRRRRRRRRRRR2C;
MO8RFFlbM0CM;O

FFlbM0CMRN1bMv4.k#G_4P4_RR
RRRRRRRRRb0Fs5RR
RRRRRRRRRRRRRQRRRRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRRm:RRR0FkR0R#8F_DoRHO
RRRRRRRRRRRRRRRR
2;CRM8ObFlFMMC0
;
ObFlFMMC0$R#MOO_DC	_MDNLCRR
RRRRRRRRRsbF0
5RRRRRRRRRRRRRRRRR7:RRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRRhB:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRRRTRF:RkR0R#_08DHFoORR
RRRRRRRRRRRRR2RR;M
C8FROlMbFC;M0
F
OlMbFCRM01tA_.kaAV#RH
MoCCOsHR
5RSRSX:MRQ0CCos
R;SRSY:MRQ0CCosSR
R;R2
bRRF5s0
RRRR:mRR0FkR8#0_oDFH
O;RRRRQRR:H#MR0D8_FOoH
RRRR
2;CRM8ObFlFMMC0
;
CRM8;



