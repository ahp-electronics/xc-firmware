-- $Header: //synplicity/maplat2018q2p1/mappers/xilinx/lib/generic/gen_generic2/cmp_eq.vhd#1 $
@E


DsHLNRs$HCCC;kR
#HCRC3CC#_08DHFoO4_4nNc3D
D;
0CMHR0$CCJ_DCClMH0R#R
RRFRbsN05jL,RjN,R4L,R4D,R0RHM:MRHR8#0_oDFH
O;RRRRRRRRRRRRRFD0kR0:FRk0#_08DHFoO
2;CRM8CCJ_DCClM
0;
s
NO0EHCkO0sCCRJFMRVJRC_CCDl0CMR
H#So#HMRND0:4RR8#0_oDFH
O;SO
SFFlbM0CMRXvzBpY_
SRSb0FsRR5
RSRSSRpm:kRF00R#8F_Do;HO
RRRSBSSQRR:H#MR0D8_FOoH;R
RRSSS7:QRRRHM#_08DHFoOR;
RSRSS:1RRRHM#_08DHFoOS
RS
2;S8CMRlOFbCFMM
0;SN--0H0sLCk0RNLDOL	_FFGRVzRvXRBY:FROlMbFCRM0H0#Rs;kC
oLCHSM
0<4R=NR54MRGFLsR4N2RM58RNGjRMRFsL;j2
RRRRGlk_#HM0RR:vBzXY
_pRRRRRRRRb0FsRblN5=1R>4R0,RR
RRRRRpRRm>R=RFD0k
0,RRRRRRRRB=QR>0RDH
M,RRRRRRRR7=QR>jR''
2;CRM8C;JM
D

HNLssH$RC;CCR#
kCCRHC#C30D8_FOoH_n44cD3ND
;
CHM00C$RJD_CCMlC0M_FC0LHR
H#RRRRb0Fs5,NjR,LjRHD0MRR:H#MR0D8_FOoH;R
RRRRRRRRRRDRR00Fk:kRF00R#8F_Do2HO;M
C8JRC_CCDl0CM_CFML;H0
N

sHOE00COkRsCCRJMFCVRJD_CCMlC0M_FC0LHR
H#So#HMRND0:4RR8#0_oDFH
O;SO
SFFlbM0CMRXvzBpY_
SRSb0FsRR5
RSRSSRpm:kRF00R#8F_Do;HO
RRRSBSSQRR:H#MR0D8_FOoH;R
RRSSS7:QRRRHM#_08DHFoOR;
RSRSS:1RRRHM#_08DHFoOS
RS
2;S8CMRlOFbCFMM
0;SN--0H0sLCk0RNLDOL	_FFGRVzRvXRBY:FROlMbFCRM0H0#Rs;kC
oLCHSM
0<4R=NR5jMRGFLsRj
2;RRRRl_kGH0M#Rv:RzYXB_Rp
RRRRRbRRFRs0l5Nb1>R=R,04RR
RRRRRRmRpRR=>Dk0F0R,
RRRRRBRRQ>R=RHD0MR,
RRRRR7RRQ>R=R''j2C;
MC8RJ
M;
D

HNLssH$RC;CCR#
kCCRHC#C30D8_FOoH_n44cD3ND
;
CHM00B$Rv u_T#RH
RRRRMoCCOsH58IH0:ERR0HMCsoCR4:=2R;
RbRRF5s0qH:RM0R#8F_Do_HOP0COFIs5HE80RR-48MFI0jFR2R;
RRRRRRRRAH:RM0R#8F_Do_HOP0COFIs5HE80RR-48MFI0jFR2R;
RRRRRRRR :TRR0FkR8#0_oDFH;O2
8CMRuBv_; T
N

sHOE00COkRsCODCD_PDCCFDRVvRBuT_ R
H#
MVkOF0HMkRVMCO_sssF5_CJI0H8ERR:HCM0o2CsR0sCkRsM#H0sMHoR#C
Lo
HMRVRHRC55JH_I8R0E>U=R2MRN8CR5JH_I8R0E<n=RcR220MEC
RRRR0sCk5sM";"2
CRRD
#CRRRRskC0s"M5CFsss;"2
CRRMH8RVC;
MV8Rk_MOCFsssN;
0H0sLCk0RMoCC0sNFss_CsbF0RR:#H0sM
o;Ns00H0LkCCRoMNCs0_FssFCbsF0RVCRODDD_CDPCRN:RsHOE00COkRsCHV#Rk_MOCFsssH5I820E;S

O#FM00NMRCH0sHN0F:MRR0HMCsoCRR:=58IH0/E2.S;
O#FM00NMRlsCN8HMC:sRR0HMCsoCRR:=58IH0RE2lRF8.R;
R#RRHNoMDNR800N_l:bRR8#0_oDFHPO_CFO0sIR5HE80R4-RRI8FMR0Fj
2;
RRRRlOFbCFMMC0RJD_CCMlC0#RH
RRRRRRRRsbF0j5N,jRL,4RN,4RL,0RDHRM:H#MR0D8_FOoH;R
RRRRRRRRRRRRRRDRR00FkRF:Rk#0R0D8_FOoH2R;
RCRRMO8RFFlbM0CM;S

ObFlFMMC0JRC_CCDl0CM_CFMLRH0HR#
RRRRRbRRF5s0NRj,LRj,DM0H:MRHR8#0_oDFH
O;RRRRRRRRRRRRRRRRRFD0k:0RR0FkR8#0_oDFH;O2
RRRR8CMRlOFbCFMM
0;LHCoMz
SjRR:HRV5I0H8ERR>4o2RCsMCN
0CSoLCHRM
RzRRj:4RR_CJClDCC
M0RRRRRRRRRRRRRRRRb0FsRblN5S
SSjSNRR=>q25j,RR
RRRRRRRRRRRRRLRRj>R=RjA52S,
SNSS4>R=R4q52
,RRRRRRRRRRRRRRRRRL=4R>5RA4
2,RRRRRRRRRRRRRRRRDM0HRR=>',4'
RRRRRRRRRRRRRRRRFD0k=0R>NR800N_ljb52
2;S8CMRMoCC0sNC
;
RRRRRRRR
4SzRH:RVI5RHE80R4=R2CRoMNCs0SC
LHCoMS
S <TR=5RqjG2RMRFsA25j;C
SMo8RCsMCN;0C
R
RR.RzRV:RFLsRHH0_MG8CRRHM4FR0R05HC0sNHRFM-2R4RCRoMNCs0RC
RRRRRLRRCMoH
RRRRRRRRRRRR4z.RC:RJD_CCMlC0R
RRRRRRRRRRRRRRFRbsl0RN
b5SSSSN=jR>5Rq.H*L0M_H82CG,RR
RRRRRRRRRRRRRLRRj>R=R.A5*0LH_8HMC,G2
SSSSRN4=q>R5L.*HH0_MG8CR4+R2
,RRRRRRRRRRRRRRRRRL=4R>5RA.H*L0M_H8RCG+2R4,R
RRRRRRRRRRRRRR0RDH=MR>NR800N_lLb5HH0_MG8CR4-R2R,
RRRRRRRRRRRRRDRR00FkRR=>8NN0_b0l50LH_8HMC2G2;R
RRRRRRMRC8CRoMNCs0
C;
dSzRH:RVs5RCHlNMs8CR4=RR8NMR8IH0>ERRR42oCCMsCN0
CSLo
HMSdSz4RR:CCJ_DCClMF0_MHCL0S
SSsbF0NRlbS5
SNSSj>R=RIq5HE80R2-4,S
SSjSLRR=>AH5I8R0E-2R4,S
SS0SDH=MR>08NNl_0b05HC0sNHRFM-2R4,S
SS0SDFRk0= >RT
2;S8CMRMoCC0sNC
;
RRRRRRRR
cSzRH:RVC5slMNH8RCs=RRjNRM8I0H8E>RRRR42oCCMsCN0
CSLo
HMRRRRSR T<8=RN_0N05lbHs0CNF0HMRR-4R2;
C
SMo8RCsMCN;0C
M
C8ORRC_DDDCCPD
;

