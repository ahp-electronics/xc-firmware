module DCUA (
   // Channel and Dual Pins
   input  CH0_HDINP, CH1_HDINP, CH0_HDINN, CH1_HDINN, D_TXBIT_CLKP_FROM_ND, D_TXBIT_CLKN_FROM_ND, D_SYNC_ND, D_TXPLL_LOL_FROM_ND,
          CH0_RX_REFCLK, CH1_RX_REFCLK, CH0_FF_RXI_CLK, CH1_FF_RXI_CLK, CH0_FF_TXI_CLK, CH1_FF_TXI_CLK, CH0_FF_EBRD_CLK, CH1_FF_EBRD_CLK,
          CH0_FF_TX_D_0, CH1_FF_TX_D_0, CH0_FF_TX_D_1, CH1_FF_TX_D_1, CH0_FF_TX_D_2, CH1_FF_TX_D_2, CH0_FF_TX_D_3, CH1_FF_TX_D_3,
          CH0_FF_TX_D_4, CH1_FF_TX_D_4, CH0_FF_TX_D_5, CH1_FF_TX_D_5, CH0_FF_TX_D_6, CH1_FF_TX_D_6, CH0_FF_TX_D_7, CH1_FF_TX_D_7,
          CH0_FF_TX_D_8, CH1_FF_TX_D_8, CH0_FF_TX_D_9, CH1_FF_TX_D_9, CH0_FF_TX_D_10, CH1_FF_TX_D_10, CH0_FF_TX_D_11, CH1_FF_TX_D_11,
          CH0_FF_TX_D_12, CH1_FF_TX_D_12, CH0_FF_TX_D_13, CH1_FF_TX_D_13, CH0_FF_TX_D_14, CH1_FF_TX_D_14, CH0_FF_TX_D_15, CH1_FF_TX_D_15,
          CH0_FF_TX_D_16, CH1_FF_TX_D_16, CH0_FF_TX_D_17, CH1_FF_TX_D_17, CH0_FF_TX_D_18, CH1_FF_TX_D_18, CH0_FF_TX_D_19, CH1_FF_TX_D_19,
          CH0_FF_TX_D_20, CH1_FF_TX_D_20, CH0_FF_TX_D_21, CH1_FF_TX_D_21, CH0_FF_TX_D_22, CH1_FF_TX_D_22, CH0_FF_TX_D_23, CH1_FF_TX_D_23,
          CH0_FFC_EI_EN, CH1_FFC_EI_EN, CH0_FFC_PCIE_DET_EN, CH1_FFC_PCIE_DET_EN, CH0_FFC_PCIE_CT, CH1_FFC_PCIE_CT, CH0_FFC_SB_INV_RX, CH1_FFC_SB_INV_RX,
          CH0_FFC_ENABLE_CGALIGN, CH1_FFC_ENABLE_CGALIGN, CH0_FFC_SIGNAL_DETECT, CH1_FFC_SIGNAL_DETECT, CH0_FFC_FB_LOOPBACK, CH1_FFC_FB_LOOPBACK, CH0_FFC_SB_PFIFO_LP, CH1_FFC_SB_PFIFO_LP,
          CH0_FFC_PFIFO_CLR, CH1_FFC_PFIFO_CLR, CH0_FFC_RATE_MODE_RX, CH1_FFC_RATE_MODE_RX, CH0_FFC_RATE_MODE_TX, CH1_FFC_RATE_MODE_TX, CH0_FFC_DIV11_MODE_RX, CH1_FFC_DIV11_MODE_RX,
          CH0_FFC_DIV11_MODE_TX, CH1_FFC_DIV11_MODE_TX, CH0_FFC_RX_GEAR_MODE, CH1_FFC_RX_GEAR_MODE, CH0_FFC_TX_GEAR_MODE, CH1_FFC_TX_GEAR_MODE, CH0_FFC_LDR_CORE2TX_EN, CH1_FFC_LDR_CORE2TX_EN,
          CH0_FFC_LANE_TX_RST, CH1_FFC_LANE_TX_RST, CH0_FFC_LANE_RX_RST, CH1_FFC_LANE_RX_RST, CH0_FFC_RRST, CH1_FFC_RRST, CH0_FFC_TXPWDNB, CH1_FFC_TXPWDNB,
          CH0_FFC_RXPWDNB, CH1_FFC_RXPWDNB, CH0_LDR_CORE2TX, CH1_LDR_CORE2TX, D_SCIWDATA0, D_SCIWDATA1, D_SCIWDATA2, D_SCIWDATA3,
          D_SCIWDATA4, D_SCIWDATA5, D_SCIWDATA6, D_SCIWDATA7, D_SCIADDR0, D_SCIADDR1, D_SCIADDR2, D_SCIADDR3,
          D_SCIADDR4, D_SCIADDR5, D_SCIENAUX, D_SCISELAUX, CH0_SCIEN, CH1_SCIEN, CH0_SCISEL, CH1_SCISEL,
          D_SCIRD, D_SCIWSTN, D_CYAWSTN, D_FFC_SYNC_TOGGLE, D_FFC_DUAL_RST, D_FFC_MACRO_RST, D_FFC_MACROPDB, D_FFC_TRST,
          CH0_FFC_CDR_EN_BITSLIP, CH1_FFC_CDR_EN_BITSLIP, D_SCAN_ENABLE, D_SCAN_IN_0, D_SCAN_IN_1, D_SCAN_IN_2, D_SCAN_IN_3, D_SCAN_IN_4,
          D_SCAN_IN_5, D_SCAN_IN_6, D_SCAN_IN_7, D_SCAN_MODE, D_SCAN_RESET, D_CIN0, D_CIN1, D_CIN2,
          D_CIN3, D_CIN4, D_CIN5, D_CIN6, D_CIN7, D_CIN8, D_CIN9, D_CIN10,
          D_CIN11,
   output CH0_HDOUTP, CH1_HDOUTP, CH0_HDOUTN, CH1_HDOUTN, D_TXBIT_CLKP_TO_ND, D_TXBIT_CLKN_TO_ND, D_SYNC_PULSE2ND, D_TXPLL_LOL_TO_ND,
          CH0_FF_RX_F_CLK, CH1_FF_RX_F_CLK, CH0_FF_RX_H_CLK, CH1_FF_RX_H_CLK, CH0_FF_TX_F_CLK, CH1_FF_TX_F_CLK, CH0_FF_TX_H_CLK, CH1_FF_TX_H_CLK,
          CH0_FF_RX_PCLK, CH1_FF_RX_PCLK, CH0_FF_TX_PCLK, CH1_FF_TX_PCLK, CH0_FF_RX_D_0, CH1_FF_RX_D_0, CH0_FF_RX_D_1, CH1_FF_RX_D_1,
          CH0_FF_RX_D_2, CH1_FF_RX_D_2, CH0_FF_RX_D_3, CH1_FF_RX_D_3, CH0_FF_RX_D_4, CH1_FF_RX_D_4, CH0_FF_RX_D_5, CH1_FF_RX_D_5,
          CH0_FF_RX_D_6, CH1_FF_RX_D_6, CH0_FF_RX_D_7, CH1_FF_RX_D_7, CH0_FF_RX_D_8, CH1_FF_RX_D_8, CH0_FF_RX_D_9, CH1_FF_RX_D_9,
          CH0_FF_RX_D_10, CH1_FF_RX_D_10, CH0_FF_RX_D_11, CH1_FF_RX_D_11, CH0_FF_RX_D_12, CH1_FF_RX_D_12, CH0_FF_RX_D_13, CH1_FF_RX_D_13,
          CH0_FF_RX_D_14, CH1_FF_RX_D_14, CH0_FF_RX_D_15, CH1_FF_RX_D_15, CH0_FF_RX_D_16, CH1_FF_RX_D_16, CH0_FF_RX_D_17, CH1_FF_RX_D_17,
          CH0_FF_RX_D_18, CH1_FF_RX_D_18, CH0_FF_RX_D_19, CH1_FF_RX_D_19, CH0_FF_RX_D_20, CH1_FF_RX_D_20, CH0_FF_RX_D_21, CH1_FF_RX_D_21,
          CH0_FF_RX_D_22, CH1_FF_RX_D_22, CH0_FF_RX_D_23, CH1_FF_RX_D_23, CH0_FFS_PCIE_DONE, CH1_FFS_PCIE_DONE, CH0_FFS_PCIE_CON, CH1_FFS_PCIE_CON,
          CH0_FFS_RLOS, CH1_FFS_RLOS, CH0_FFS_LS_SYNC_STATUS, CH1_FFS_LS_SYNC_STATUS, CH0_FFS_CC_UNDERRUN, CH1_FFS_CC_UNDERRUN, CH0_FFS_CC_OVERRUN, CH1_FFS_CC_OVERRUN,
          CH0_FFS_RXFBFIFO_ERROR, CH1_FFS_RXFBFIFO_ERROR, CH0_FFS_TXFBFIFO_ERROR, CH1_FFS_TXFBFIFO_ERROR, CH0_FFS_RLOL, CH1_FFS_RLOL, CH0_FFS_SKP_ADDED, CH1_FFS_SKP_ADDED,
          CH0_FFS_SKP_DELETED, CH1_FFS_SKP_DELETED, CH0_LDR_RX2CORE, CH1_LDR_RX2CORE, D_SCIRDATA0, D_SCIRDATA1, D_SCIRDATA2, D_SCIRDATA3,
          D_SCIRDATA4, D_SCIRDATA5, D_SCIRDATA6, D_SCIRDATA7, D_SCIINT, D_SCAN_OUT_0, D_SCAN_OUT_1, D_SCAN_OUT_2,
          D_SCAN_OUT_3, D_SCAN_OUT_4, D_SCAN_OUT_5, D_SCAN_OUT_6, D_SCAN_OUT_7, D_COUT0, D_COUT1, D_COUT2,
          D_COUT3, D_COUT4, D_COUT5, D_COUT6, D_COUT7, D_COUT8, D_COUT9, D_COUT10,
          D_COUT11, D_COUT12, D_COUT13, D_COUT14, D_COUT15, D_COUT16, D_COUT17, D_COUT18,
          D_COUT19,
   // No of ports = 161 inputs + 129 outputs = 290

   // PLL Pins
   input  D_REFCLKI,
   output D_FFS_PLOL
   // No of ports = 1 inputs + 1 outputs = 2

   // Total no of ports = 292
  ); //synthesis syn_black_box

   // Ch_Dual_Attr
   parameter D_MACROPDB = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter D_IB_PWDNB = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter D_XGE_MODE = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter D_LOW_MARK = "DONTCARE"; //"DONTCARE" "0d0"-"0d15"
   parameter D_HIGH_MARK = "DONTCARE"; //"DONTCARE" "0d0"-"0d15"
   parameter D_BUS8BIT_SEL = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter D_CDR_LOL_SET = "DONTCARE"; //"DONTCARE" "0b00"-"0b11"
   parameter D_TXPLL_PWDNB = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter D_BITCLK_LOCAL_EN = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter D_BITCLK_ND_EN = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter D_BITCLK_FROM_ND_EN = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter D_SYNC_LOCAL_EN = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter D_SYNC_ND_EN = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH0_UC_MODE = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH1_UC_MODE = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH0_PCIE_MODE = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH1_PCIE_MODE = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH0_RIO_MODE = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH1_RIO_MODE = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH0_WA_MODE = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH1_WA_MODE = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH0_INVERT_RX = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH1_INVERT_RX = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH0_INVERT_TX = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH1_INVERT_TX = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH0_PRBS_SELECTION = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH1_PRBS_SELECTION = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH0_GE_AN_ENABLE = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH1_GE_AN_ENABLE = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH0_PRBS_LOCK = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH1_PRBS_LOCK = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH0_PRBS_ENABLE = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH1_PRBS_ENABLE = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH0_ENABLE_CG_ALIGN = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH1_ENABLE_CG_ALIGN = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH0_TX_GEAR_MODE = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH1_TX_GEAR_MODE = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH0_RX_GEAR_MODE = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH1_RX_GEAR_MODE = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH0_PCS_DET_TIME_SEL = "DONTCARE"; //"DONTCARE" "0b00"-"0b11"
   parameter CH1_PCS_DET_TIME_SEL = "DONTCARE"; //"DONTCARE" "0b00"-"0b11"
   parameter CH0_PCIE_EI_EN = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH1_PCIE_EI_EN = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH0_TX_GEAR_BYPASS = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH1_TX_GEAR_BYPASS = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH0_ENC_BYPASS = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH1_ENC_BYPASS = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH0_SB_BYPASS = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH1_SB_BYPASS = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH0_RX_SB_BYPASS = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH1_RX_SB_BYPASS = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH0_WA_BYPASS = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH1_WA_BYPASS = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH0_DEC_BYPASS = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH1_DEC_BYPASS = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH0_CTC_BYPASS = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH1_CTC_BYPASS = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH0_RX_GEAR_BYPASS = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH1_RX_GEAR_BYPASS = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH0_LSM_DISABLE = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH1_LSM_DISABLE = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH0_MATCH_2_ENABLE = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH1_MATCH_2_ENABLE = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH0_MATCH_4_ENABLE = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH1_MATCH_4_ENABLE = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH0_MIN_IPG_CNT = "DONTCARE"; //"DONTCARE" "0b00"-"0b11"
   parameter CH1_MIN_IPG_CNT = "DONTCARE"; //"DONTCARE" "0b00"-"0b11"
   parameter CH0_CC_MATCH_1 = "DONTCARE"; //"DONTCARE" "0x000"-"0x3ff"
   parameter CH1_CC_MATCH_1 = "DONTCARE"; //"DONTCARE" "0x000"-"0x3ff"
   parameter CH0_CC_MATCH_2 = "DONTCARE"; //"DONTCARE" "0x000"-"0x3ff"
   parameter CH1_CC_MATCH_2 = "DONTCARE"; //"DONTCARE" "0x000"-"0x3ff"
   parameter CH0_CC_MATCH_3 = "DONTCARE"; //"DONTCARE" "0x000"-"0x3ff"
   parameter CH1_CC_MATCH_3 = "DONTCARE"; //"DONTCARE" "0x000"-"0x3ff"
   parameter CH0_CC_MATCH_4 = "DONTCARE"; //"DONTCARE" "0x000"-"0x3ff"
   parameter CH1_CC_MATCH_4 = "DONTCARE"; //"DONTCARE" "0x000"-"0x3ff"
   parameter CH0_UDF_COMMA_MASK = "DONTCARE"; //"DONTCARE" "0x000"-"0x3ff"
   parameter CH1_UDF_COMMA_MASK = "DONTCARE"; //"DONTCARE" "0x000"-"0x3ff"
   parameter CH0_UDF_COMMA_A = "DONTCARE"; //"DONTCARE" "0x000"-"0x3ff"
   parameter CH1_UDF_COMMA_A = "DONTCARE"; //"DONTCARE" "0x000"-"0x3ff"
   parameter CH0_UDF_COMMA_B = "DONTCARE"; //"DONTCARE" "0x000"-"0x3ff"
   parameter CH1_UDF_COMMA_B = "DONTCARE"; //"DONTCARE" "0x000"-"0x3ff"
   parameter CH0_RX_DCO_CK_DIV = "DONTCARE"; //"DONTCARE" "0b000"-"0b111"
   parameter CH1_RX_DCO_CK_DIV = "DONTCARE"; //"DONTCARE" "0b000"-"0b111"
   parameter CH0_RCV_DCC_EN = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH1_RCV_DCC_EN = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH0_TPWDNB = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH1_TPWDNB = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH0_RATE_MODE_TX = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH1_RATE_MODE_TX = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH0_RTERM_TX = "DONTCARE"; //"DONTCARE" "0d0"-"0d31"
   parameter CH1_RTERM_TX = "DONTCARE"; //"DONTCARE" "0d0"-"0d31"
   parameter CH0_TX_CM_SEL = "DONTCARE"; //"DONTCARE" "0b00"-"0b11"
   parameter CH1_TX_CM_SEL = "DONTCARE"; //"DONTCARE" "0b00"-"0b11"
   parameter CH0_TDRV_PRE_EN = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH1_TDRV_PRE_EN = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH0_TDRV_SLICE0_SEL = "DONTCARE"; //"DONTCARE" "0b00"-"0b11"
   parameter CH1_TDRV_SLICE0_SEL = "DONTCARE"; //"DONTCARE" "0b00"-"0b11"
   parameter CH0_TDRV_SLICE1_SEL = "DONTCARE"; //"DONTCARE" "0b00"-"0b11"
   parameter CH1_TDRV_SLICE1_SEL = "DONTCARE"; //"DONTCARE" "0b00"-"0b11"
   parameter CH0_TDRV_SLICE2_SEL = "DONTCARE"; //"DONTCARE" "0b00"-"0b11"
   parameter CH1_TDRV_SLICE2_SEL = "DONTCARE"; //"DONTCARE" "0b00"-"0b11"
   parameter CH0_TDRV_SLICE3_SEL = "DONTCARE"; //"DONTCARE" "0b00"-"0b11"
   parameter CH1_TDRV_SLICE3_SEL = "DONTCARE"; //"DONTCARE" "0b00"-"0b11"
   parameter CH0_TDRV_SLICE4_SEL = "DONTCARE"; //"DONTCARE" "0b00"-"0b11"
   parameter CH1_TDRV_SLICE4_SEL = "DONTCARE"; //"DONTCARE" "0b00"-"0b11"
   parameter CH0_TDRV_SLICE5_SEL = "DONTCARE"; //"DONTCARE" "0b00"-"0b11"
   parameter CH1_TDRV_SLICE5_SEL = "DONTCARE"; //"DONTCARE" "0b00"-"0b11"
   parameter CH0_TDRV_SLICE0_CUR = "DONTCARE"; //"DONTCARE" "0b000"-"0b111"
   parameter CH1_TDRV_SLICE0_CUR = "DONTCARE"; //"DONTCARE" "0b000"-"0b111"
   parameter CH0_TDRV_SLICE1_CUR = "DONTCARE"; //"DONTCARE" "0b000"-"0b111"
   parameter CH1_TDRV_SLICE1_CUR = "DONTCARE"; //"DONTCARE" "0b000"-"0b111"
   parameter CH0_TDRV_SLICE2_CUR = "DONTCARE"; //"DONTCARE" "0b00"-"0b11"
   parameter CH1_TDRV_SLICE2_CUR = "DONTCARE"; //"DONTCARE" "0b00"-"0b11"
   parameter CH0_TDRV_SLICE3_CUR = "DONTCARE"; //"DONTCARE" "0b00"-"0b11"
   parameter CH1_TDRV_SLICE3_CUR = "DONTCARE"; //"DONTCARE" "0b00"-"0b11"
   parameter CH0_TDRV_SLICE4_CUR = "DONTCARE"; //"DONTCARE" "0b00"-"0b11"
   parameter CH1_TDRV_SLICE4_CUR = "DONTCARE"; //"DONTCARE" "0b00"-"0b11"
   parameter CH0_TDRV_SLICE5_CUR = "DONTCARE"; //"DONTCARE" "0b00"-"0b11"
   parameter CH1_TDRV_SLICE5_CUR = "DONTCARE"; //"DONTCARE" "0b00"-"0b11"
   parameter CH0_TDRV_DAT_SEL = "DONTCARE"; //"DONTCARE" "0b00"-"0b11"
   parameter CH1_TDRV_DAT_SEL = "DONTCARE"; //"DONTCARE" "0b00"-"0b11"
   parameter CH0_TX_DIV11_SEL = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH1_TX_DIV11_SEL = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH0_RPWDNB = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH1_RPWDNB = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH0_RATE_MODE_RX = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH1_RATE_MODE_RX = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH0_RX_DIV11_SEL = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH1_RX_DIV11_SEL = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH0_SEL_SD_RX_CLK = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH1_SEL_SD_RX_CLK = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH0_FF_RX_H_CLK_EN = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH1_FF_RX_H_CLK_EN = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH0_FF_RX_F_CLK_DIS = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH1_FF_RX_F_CLK_DIS = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH0_FF_TX_H_CLK_EN = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH1_FF_TX_H_CLK_EN = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH0_FF_TX_F_CLK_DIS = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH1_FF_TX_F_CLK_DIS = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH0_TDRV_POST_EN = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH1_TDRV_POST_EN = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH0_TX_POST_SIGN = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH1_TX_POST_SIGN = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH0_TX_PRE_SIGN = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH1_TX_PRE_SIGN = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH0_REQ_LVL_SET = "DONTCARE"; //"DONTCARE" "0b00"-"0b11"
   parameter CH1_REQ_LVL_SET = "DONTCARE"; //"DONTCARE" "0b00"-"0b11"
   parameter CH0_REQ_EN = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH1_REQ_EN = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH0_RTERM_RX = "DONTCARE"; //"DONTCARE" "0d0"-"0d31"
   parameter CH1_RTERM_RX = "DONTCARE"; //"DONTCARE" "0d0"-"0d31"
   parameter CH0_RXTERM_CM = "DONTCARE"; //"DONTCARE" "0b00"-"0b11"
   parameter CH1_RXTERM_CM = "DONTCARE"; //"DONTCARE" "0b00"-"0b11"
   parameter CH0_PDEN_SEL = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH1_PDEN_SEL = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH0_RXIN_CM = "DONTCARE"; //"DONTCARE" "0b00"-"0b11"
   parameter CH1_RXIN_CM = "DONTCARE"; //"DONTCARE" "0b00"-"0b11"
   parameter CH0_LEQ_OFFSET_SEL = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH1_LEQ_OFFSET_SEL = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH0_LEQ_OFFSET_TRIM = "DONTCARE"; //"DONTCARE" "0b000"-"0b111"
   parameter CH1_LEQ_OFFSET_TRIM = "DONTCARE"; //"DONTCARE" "0b000"-"0b111"
   parameter CH0_RLOS_SEL = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH1_RLOS_SEL = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH0_RX_LOS_LVL = "DONTCARE"; //"DONTCARE" "0b000"-"0b111"
   parameter CH1_RX_LOS_LVL = "DONTCARE"; //"DONTCARE" "0b000"-"0b111"
   parameter CH0_RX_LOS_CEQ = "DONTCARE"; //"DONTCARE" "0b00"-"0b11"
   parameter CH1_RX_LOS_CEQ = "DONTCARE"; //"DONTCARE" "0b00"-"0b11"
   parameter CH0_RX_LOS_HYST_EN = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH1_RX_LOS_HYST_EN = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH0_RX_LOS_EN = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH1_RX_LOS_EN = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH0_LDR_RX2CORE_SEL = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH1_LDR_RX2CORE_SEL = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH0_LDR_CORE2TX_SEL = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH1_LDR_CORE2TX_SEL = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter D_TX_MAX_RATE = "DONTCARE"; //"DONTCARE" "0.27"-"3.125"
   parameter CH0_CDR_MAX_RATE = "DONTCARE"; //"DONTCARE" "0.27"-"3.125"
   parameter CH1_CDR_MAX_RATE = "DONTCARE"; //"DONTCARE" "0.27"-"3.125"
   parameter CH0_TXAMPLITUDE = "DONTCARE"; //"DONTCARE" "0d0"-"0d1300"
   parameter CH1_TXAMPLITUDE = "DONTCARE"; //"DONTCARE" "0d0"-"0d1300"
   parameter CH0_TXDEPRE = "DONTCARE"; //"DONTCARE" "DISABLED" "0d0"-"0d11"
   parameter CH1_TXDEPRE = "DONTCARE"; //"DONTCARE" "DISABLED" "0d0"-"0d11"
   parameter CH0_TXDEPOST = "DONTCARE"; //"DONTCARE" "DISABLED" "0d0"-"0d11"
   parameter CH1_TXDEPOST = "DONTCARE"; //"DONTCARE" "DISABLED" "0d0"-"0d11"
   parameter CH0_PROTOCOL = "DONTCARE"; //"DONTCARE" "PCIE" "GBE" "SGMII" "XAUI" "SDI" "CPRI" "JESD204" "EDP" "G8B10B" "8BSER" "10BSER"
   parameter CH1_PROTOCOL = "DONTCARE"; //"DONTCARE" "PCIE" "GBE" "SGMII" "XAUI" "SDI" "CPRI" "JESD204" "EDP" "G8B10B" "8BSER" "10BSER"
   // No of parameters = 186

   // Analog_Attr
   parameter D_ISETLOS = "DONTCARE"; //"DONTCARE" "0d0"-"0d255"
   parameter D_SETIRPOLY_AUX = "DONTCARE"; //"DONTCARE" "0b00"-"0b11"
   parameter D_SETICONST_AUX = "DONTCARE"; //"DONTCARE" "0b00"-"0b11"
   parameter D_SETIRPOLY_CH = "DONTCARE"; //"DONTCARE" "0b00"-"0b11"
   parameter D_SETICONST_CH = "DONTCARE"; //"DONTCARE" "0b00"-"0b11"
   parameter D_REQ_ISET = "DONTCARE"; //"DONTCARE" "0b000"-"0b111"
   parameter D_PD_ISET = "DONTCARE"; //"DONTCARE" "0b00"-"0b11"
   parameter D_DCO_CALIB_TIME_SEL = "DONTCARE"; //"DONTCARE" "0b00"-"0b11"
   parameter CH0_CDR_CNT4SEL = "DONTCARE"; //"DONTCARE" "0b00"-"0b11"
   parameter CH1_CDR_CNT4SEL = "DONTCARE"; //"DONTCARE" "0b00"-"0b11"
   parameter CH0_CDR_CNT8SEL = "DONTCARE"; //"DONTCARE" "0b00"-"0b11"
   parameter CH1_CDR_CNT8SEL = "DONTCARE"; //"DONTCARE" "0b00"-"0b11"
   parameter CH0_DCOATDCFG = "DONTCARE"; //"DONTCARE" "0b00"-"0b11"
   parameter CH1_DCOATDCFG = "DONTCARE"; //"DONTCARE" "0b00"-"0b11"
   parameter CH0_DCOATDDLY = "DONTCARE"; //"DONTCARE" "0b00"-"0b11"
   parameter CH1_DCOATDDLY = "DONTCARE"; //"DONTCARE" "0b00"-"0b11"
   parameter CH0_DCOBYPSATD = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH1_DCOBYPSATD = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH0_DCOCALDIV = "DONTCARE"; //"DONTCARE" "0b000"-"0b111"
   parameter CH1_DCOCALDIV = "DONTCARE"; //"DONTCARE" "0b000"-"0b111"
   parameter CH0_DCOCTLGI = "DONTCARE"; //"DONTCARE" "0b000"-"0b111"
   parameter CH1_DCOCTLGI = "DONTCARE"; //"DONTCARE" "0b000"-"0b111"
   parameter CH0_DCODISBDAVOID = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH1_DCODISBDAVOID = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH0_DCOFLTDAC = "DONTCARE"; //"DONTCARE" "0b00"-"0b11"
   parameter CH1_DCOFLTDAC = "DONTCARE"; //"DONTCARE" "0b00"-"0b11"
   parameter CH0_DCOFTNRG = "DONTCARE"; //"DONTCARE" "0b000"-"0b111"
   parameter CH1_DCOFTNRG = "DONTCARE"; //"DONTCARE" "0b000"-"0b111"
   parameter CH0_DCOIOSTUNE = "DONTCARE"; //"DONTCARE" "0b000"-"0b111"
   parameter CH1_DCOIOSTUNE = "DONTCARE"; //"DONTCARE" "0b000"-"0b111"
   parameter CH0_DCOITUNE = "DONTCARE"; //"DONTCARE" "0b00"-"0b11"
   parameter CH1_DCOITUNE = "DONTCARE"; //"DONTCARE" "0b00"-"0b11"
   parameter CH0_DCOITUNE4LSB = "DONTCARE"; //"DONTCARE" "0b000"-"0b111"
   parameter CH1_DCOITUNE4LSB = "DONTCARE"; //"DONTCARE" "0b000"-"0b111"
   parameter CH0_DCOIUPDNX2 = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH1_DCOIUPDNX2 = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH0_DCONUOFLSB = "DONTCARE"; //"DONTCARE" "0b000"-"0b111"
   parameter CH1_DCONUOFLSB = "DONTCARE"; //"DONTCARE" "0b000"-"0b111"
   parameter CH0_DCOSCALEI = "DONTCARE"; //"DONTCARE" "0b00"-"0b11"
   parameter CH1_DCOSCALEI = "DONTCARE"; //"DONTCARE" "0b00"-"0b11"
   parameter CH0_DCOSTARTVAL = "DONTCARE"; //"DONTCARE" "0b000"-"0b111"
   parameter CH1_DCOSTARTVAL = "DONTCARE"; //"DONTCARE" "0b000"-"0b111"
   parameter CH0_DCOSTEP = "DONTCARE"; //"DONTCARE" "0b00"-"0b11"
   parameter CH1_DCOSTEP = "DONTCARE"; //"DONTCARE" "0b00"-"0b11"
   parameter CH0_BAND_THRESHOLD = "DONTCARE"; //"DONTCARE" "0d0"-"0d63"
   parameter CH1_BAND_THRESHOLD = "DONTCARE"; //"DONTCARE" "0d0"-"0d63"
   parameter CH0_AUTO_FACQ_EN = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH1_AUTO_FACQ_EN = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH0_AUTO_CALIB_EN = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH1_AUTO_CALIB_EN = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH0_CALIB_CK_MODE = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH1_CALIB_CK_MODE = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH0_REG_BAND_OFFSET = "DONTCARE"; //"DONTCARE" "0d0"-"0d15"
   parameter CH1_REG_BAND_OFFSET = "DONTCARE"; //"DONTCARE" "0d0"-"0d15"
   parameter CH0_REG_BAND_SEL = "DONTCARE"; //"DONTCARE" "0d0"-"0d63"
   parameter CH1_REG_BAND_SEL = "DONTCARE"; //"DONTCARE" "0d0"-"0d63"
   parameter CH0_REG_IDAC_SEL = "DONTCARE"; //"DONTCARE" "0d0"-"0d1023"
   parameter CH1_REG_IDAC_SEL = "DONTCARE"; //"DONTCARE" "0d0"-"0d1023"
   parameter CH0_REG_IDAC_EN = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter CH1_REG_IDAC_EN = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter D_CMUSETISCL4VCO = "DONTCARE"; //"DONTCARE" "0b000"-"0b111"
   parameter D_CMUSETI4VCO = "DONTCARE"; //"DONTCARE" "0b00"-"0b11"
   parameter D_CMUSETINITVCT = "DONTCARE"; //"DONTCARE" "0b00"-"0b11"
   parameter D_CMUSETZGM = "DONTCARE"; //"DONTCARE" "0b000"-"0b111"
   parameter D_CMUSETP2AGM = "DONTCARE"; //"DONTCARE" "0b000"-"0b111"
   parameter D_CMUSETP1GM = "DONTCARE"; //"DONTCARE" "0b000"-"0b111"
   parameter D_CMUSETI4CPZ = "DONTCARE"; //"DONTCARE" "0d0"-"0d15"
   parameter D_CMUSETI4CPP = "DONTCARE"; //"DONTCARE" "0d0"-"0d15"
   parameter D_CMUSETICP4Z = "DONTCARE"; //"DONTCARE" "0b000"-"0b111"
   parameter D_CMUSETICP4P = "DONTCARE"; //"DONTCARE" "0b00"-"0b11"
   parameter D_CMUSETBIASI = "DONTCARE"; //"DONTCARE" "0b00"-"0b11"
   parameter D_SETPLLRC = "DONTCARE"; //"DONTCARE" "0d0"-"0d63"
   parameter CH0_RX_RATE_SEL = "DONTCARE"; //"DONTCARE" "0d0"-"0d15"
   parameter CH1_RX_RATE_SEL = "DONTCARE"; //"DONTCARE" "0d0"-"0d15"
   // No of parameters = 74

   // PLL Attr
   parameter D_REFCK_MODE = "DONTCARE"; //"DONTCARE" "0b000"-"0b100"
   parameter D_TX_VCO_CK_DIV = "DONTCARE"; //"DONTCARE" "0b000"-"0b111"
   parameter D_PLL_LOL_SET = "DONTCARE"; //"DONTCARE" "0b00"-"0b11"
   parameter D_RG_EN = "DONTCARE"; //"DONTCARE" "0b0" "0b1"
   parameter D_RG_SET = "DONTCARE"; //"DONTCARE" "0b00"-"0b11"
   // No of parameters = 5

   // Total no of parameters = 265
endmodule

