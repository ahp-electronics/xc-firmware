module MUX2(O,I0,I1,S0);  // synthesis syn_black_box
input I0,I1,S0;
output O;
endmodule
module MUX4(O,I0,I1,I2,I3,S0,S1);  // synthesis syn_black_box
input I0,I1,I2,I3,S0,S1;
output O;
endmodule
module AND2 (O,I0,I1);   // synthesis syn_black_box
input I0,I1; 
output O; 
endmodule
module AND3 (O,I0,I1,I2);   // synthesis syn_black_box
input I0,I1,I2; 
output O; 
endmodule
module AND4 (O,I0,I1,I2,I3);   // synthesis syn_black_box
input I0,I1,I2,I3; 
output O; 
endmodule
module AND5 (O,I0,I1,I2,I3,I4);   // synthesis syn_black_box
input I0,I1,I2,I3,I4; 
output O; 
endmodule
module AND6 (O,I0,I1,I2,I3,I4,I5);   // synthesis syn_black_box
input I0,I1,I2,I3,I4,I5; 
output O; 
endmodule
module AND7 (O,I0,I1,I2,I3,I4,I5,I6);   // synthesis syn_black_box
input I0,I1,I2,I3,I4,I5,I6; 
output O; 
endmodule
module AND8 (O,I0,I1,I2,I3,I4,I5,I6,I7);   // synthesis syn_black_box
input I0,I1,I2,I3,I4,I5,I6,I7; 
output O; 
endmodule
module BI_DIR (O,I0,IO,OE);   // synthesis syn_black_box black_box_pad_pin="IO"
input I0,OE; 
inout IO; 
output O; 
endmodule
module BUFF (O,I0);   // synthesis syn_black_box
input I0; 
output O; 
endmodule
module BUFTH (O,I0,OE);  // synthesis syn_black_box black_box_pad_pin="O"
input I0,OE; 
output O; 
endmodule
module BUFTI (O,I0,OE);  // synthesis syn_black_box black_box_pad_pin="O"
input I0,OE; 
output O; 
endmodule
module BUFTL (O,I0,OE);  // synthesis syn_black_box black_box_pad_pin="O" 
input I0,OE; 
output O; 
endmodule
module CLKI(O,PAD);   // synthesis syn_black_box black_box_pad_pin="PAD"
input PAD; 
output O; 
endmodule
module DFF (Q,D,CLK);   // synthesis syn_black_box
input D,CLK; 
output Q; 
endmodule
module DFFC (Q,D,CLK,CE);   // synthesis syn_black_box
input D,CLK,CE; 
output Q; 
endmodule
module DFFCR (Q,D,CLK,CE,R);   // synthesis syn_black_box
input D,CLK,CE,R; 
output Q; 
endmodule
module DFFCRH (Q,D,CLK,CE,R);   // synthesis syn_black_box
input D,CLK,CE,R; 
output Q; 
endmodule
module DFFCRS (Q,D,CLK,CE,R,S);   // synthesis syn_black_box
input D,CLK,CE,R,S; 
output Q; 
endmodule
module DFFCRSH (Q,D,CLK,CE,R,S);   // synthesis syn_black_box
input D,CLK,CE,R,S; 
output Q; 
endmodule
module DFFCS (Q,D,CLK,CE,S);   // synthesis syn_black_box
input D,CLK,CE,S; 
output Q; 
endmodule
module DFFCSH (Q,D,CLK,CE,S);   // synthesis syn_black_box
input D,CLK,CE,S; 
output Q; 
endmodule
module DFFR (Q,D,CLK,R);   // synthesis syn_black_box
input D,CLK,R; 
output Q; 
endmodule
module DFFRH (Q,D,CLK,R);   // synthesis syn_black_box
input D,CLK,R; 
output Q; 
endmodule
module DFFRS (Q,D,CLK,R,S);   // synthesis syn_black_box
input D,CLK,R,S; 
output Q; 
endmodule
module DFFRSH (Q,D,CLK,R,S);   // synthesis syn_black_box
input D,CLK,R,S; 
output Q; 
endmodule
module DFFS (Q,D,CLK,S);   // synthesis syn_black_box
input D,CLK,S; 
output Q;
endmodule
module DFFSH (Q,D,CLK,S);   // synthesis syn_black_box
input D,CLK,S; 
output Q; 
endmodule
module DLAT (Q,D,LAT);   // synthesis syn_black_box
input D,LAT; 
output Q; 
endmodule
module DLATR (Q,D,LAT,R);   // synthesis syn_black_box
input D,LAT,R; 
output Q; 
endmodule 
module DLATRH (Q,D,LAT,R);   // synthesis syn_black_box
input D,LAT,R; 
output Q; 
endmodule 
module DLATRS (Q,D,LAT,R,S);   // synthesis syn_black_box
input D,LAT,R,S; 
output Q; 
endmodule 
module DLATRSH (Q,D,LAT,R,S);   // synthesis syn_black_box
input D,LAT,R,S; 
output Q; 
endmodule 
module DLATS (Q,D,LAT,S);   // synthesis syn_black_box
input D,LAT,S; 
output Q; 
endmodule 
module DLATSH (Q,D,LAT,S);   // synthesis syn_black_box
input D,LAT,S; 
output Q; 
endmodule 
module VCC (X);  // synthesis syn_black_box
output X; 
endmodule 
module GND (X);   // synthesis syn_black_box
output X; 
endmodule 
module GSRBUF (O,SRI);   // synthesis syn_black_box black_box_pad_pin="SRI"
input SRI; 
output O; 
endmodule 
module IBUF (O,I0);   // synthesis syn_black_box black_box_pad_pin="I0"
input I0; 
output O; 
endmodule 
module INV (O,I0);   // synthesis syn_black_box
input I0; 
output O; 
endmodule 
module INVTH (O,I0,OE);   // synthesis syn_black_box black_box_pad_pin="O"
input I0,OE; 
output O; 
endmodule 
module LVPECLIN (O,P_IN,N_IN);   // synthesis syn_black_box black_box_pad_pin="P_IN,N_IN"
input P_IN,N_IN; 
output O; 
endmodule 
module LVPECLOUT (P_OUT,N_OUT,I);   // synthesis syn_black_box black_box_pad_pin="P_OUT,N_OUT"
input I; 
output P_OUT,N_OUT; 
endmodule 
module LVPECLTRI (N_OUT,P_OUT,I,OE);    // synthesis syn_black_box black_box_pad_pin="P_OUT,N_OUT"
input I,OE; 
output N_OUT, P_OUT; 
endmodule 
module INVTL (O,I0,OE);    // synthesis syn_black_box black_box_pad_pin="O"
input I0,OE; 
output O; 
endmodule 
module NAN2 (O,I0,I1);   // synthesis syn_black_box
input I0,I1; 
output O; 
endmodule 
module NAN3 (O,I0,I1,I2);   // synthesis syn_black_box
input I0,I1,I2; 
output O; 
endmodule 
module NAN4 (O,I0,I1,I2,I3);   // synthesis syn_black_box
input I0,I1,I2,I3; 
output O; 
endmodule 
module NAN5 (O,I0,I1,I2,I3,I4);   // synthesis syn_black_box
input I0,I1,I2,I3,I4; 
output O; 
endmodule 
module NAN6 (O,I0,I1,I2,I3,I4,I5);   // synthesis syn_black_box
input I0,I1,I2,I3,I4,I5; 
output O; 
endmodule 
module NAN7 (O,I0,I1,I2,I3,I4,I5,I6);   // synthesis syn_black_box
input I0,I1,I2,I3,I4,I5,I6; 
output O; 
endmodule 
module NAN8 (O,I0,I1,I2,I3,I4,I5,I6,I7);   // synthesis syn_black_box
input I0,I1,I2,I3,I4,I5,I6,I7; 
output O; 
endmodule 
module NOR2 (O,I0,I1);   // synthesis syn_black_box
input I0,I1; 
output O; 
endmodule 
module NOR3 (O,I0,I1,I2);   // synthesis syn_black_box
input I0,I1,I2; 
output O; 
endmodule 
module NOR4 (O,I0,I1,I2,I3);   // synthesis syn_black_box
input I0,I1,I2,I3; 
output O; 
endmodule 
module NOR5 (O,I0,I1,I2,I3,I4);   // synthesis syn_black_box
input I0,I1,I2,I3,I4; 
output O; 
endmodule 
module NOR6 (O,I0,I1,I2,I3,I4,I5);   // synthesis syn_black_box
input I0,I1,I2,I3,I4,I5; 
output O; 
endmodule 
module NOR7 (O,I0,I1,I2,I3,I4,I5,I6);   // synthesis syn_black_box
input I0,I1,I2,I3,I4,I5,I6; 
output O; 
endmodule 
module NOR8 (O,I0,I1,I2,I3,I4,I5,I6,I7);   // synthesis syn_black_box
input I0,I1,I2,I3,I4,I5,I6,I7; 
output O; 
endmodule 
module OBUF (O,I0);    // synthesis syn_black_box black_box_pad_pin="O"
input I0; 
output O; 
endmodule 
module OR2 (O,I0,I1);   // synthesis syn_black_box
input I0,I1; 
output O; 
endmodule 
module OR3 (O,I0,I1,I2);   // synthesis syn_black_box
input I0,I1,I2; 
output O; 
endmodule 
module OR4 (O,I0,I1,I2,I3);   // synthesis syn_black_box
input I0,I1,I2,I3; 
output O; 
endmodule 
module OR5 (O,I0,I1,I2,I3,I4);   // synthesis syn_black_box
input I0,I1,I2,I3,I4; 
output O; 
endmodule 
module OR6 (O,I0,I1,I2,I3,I4,I5);   // synthesis syn_black_box
input I0,I1,I2,I3,I4,I5; 
output O; 
endmodule 
module OR7 (O,I0,I1,I2,I3,I4,I5,I6);   // synthesis syn_black_box
input I0,I1,I2,I3,I4,I5,I6; 
output O; 
endmodule 
module OR8 (O,I0,I1,I2,I3,I4,I5,I6,I7);   // synthesis syn_black_box
input I0,I1,I2,I3,I4,I5,I6,I7; 
output O; 
endmodule 
module TFF (Q,T,CLK);   // synthesis syn_black_box
input T,CLK; 
output Q; 
endmodule 
module TFFR (Q,T,CLK,R);   // synthesis syn_black_box
input T,CLK,R; 
output Q; 
endmodule 
module TFFRH (Q,T,CLK,R);   // synthesis syn_black_box
input T,CLK,R; 
output Q; 
endmodule 
module TFFRS (Q,T,CLK,R,S);   // synthesis syn_black_box
input T,CLK,R,S; 
output Q; 
endmodule 
module TFFRSH (Q,T,CLK,R,S);   // synthesis syn_black_box
input T,CLK,R,S; 
output Q; 
endmodule 
module TFFS (Q,T,CLK,S);   // synthesis syn_black_box
input T,CLK,S; 
output Q; 
endmodule 
module TFFSH (Q,T,CLK,S);   // synthesis syn_black_box
input T,CLK,S; 
output Q; 
endmodule 
module XOR2 (O,I0,I1);   // synthesis syn_black_box
input I0,I1; 
output O; 
endmodule 
module XORSOFT (O,I0,I1);   // synthesis syn_black_box
input I0,I1; 
output O; 
endmodule 
//PLL BLOCK cells
//SPLL Software Usage Model 7.09 -QQ
module SPLL(CLK_IN, CLK_OUT);   // synthesis syn_black_box black_box_pad_pin="CLK_IN"
parameter in_freq = "1";
parameter clk_out_to_pin =  "OFF";
parameter wake_on_lock = "OFF";
input  CLK_IN;
output CLK_OUT;
endmodule
//STDPLL Software Usage Model 7.09 -QQ
module STDPLL(CLK_IN, PLL_LOCK, CLK_OUT);   // synthesis syn_black_box black_box_pad_pin="CLK_IN"
parameter in_freq = "1";
parameter mult = "1";
parameter div = "1";
parameter post = "1";
parameter pll_dly = "1";
parameter clk_out_to_pin = "OFF";
parameter wake_on_lock = "OFF";
input  CLK_IN;
output CLK_OUT;
output PLL_LOCK;
endmodule
//STDPLLX Software Usage Model 7.09 -QQ
module STDPLLX(CLK_IN, PLL_FBK, PLL_RST, PLL_LOCK, SEC_OUT, CLK_OUT);   // synthesis syn_black_box black_box_pad_pin="CLK_IN"
parameter in_freq = "1";
parameter mult = "1";
parameter div = "1";
parameter post = "1";
parameter pll_dly = "1";
parameter secdiv = "1";
parameter clk_out_to_pin = "ON";
parameter wake_on_lock = "OFF";
input  CLK_IN;	
input  PLL_FBK;		 
input  PLL_RST;		
output CLK_OUT;
output PLL_LOCK;
output SEC_OUT;
endmodule
//LVDS BLOCK cells
module LVDSIN (O, P_IN,N_IN);    // synthesis syn_black_box black_box_pad_pin="P_IN,N_IN"
input P_IN,N_IN; 
output O; 
endmodule 
module LVDSOUT (P_OUT,N_OUT, I);    // synthesis syn_black_box black_box_pad_pin="P_OUT,N_OUT"
input I; 
output P_OUT,N_OUT; 
endmodule 
module LVDSTRI (P_OUT,N_OUT, I,OE);    // synthesis syn_black_box black_box_pad_pin="P_OUT,N_OUT"
input I,OE; 
output P_OUT,N_OUT; 
endmodule 
module LVDSIO (O, P_IO, N_IO, I, OE);    // synthesis syn_black_box black_box_pad_pin="P_IO,N_IO"
input I,OE; 
inout P_IO,N_IO; 
output O;
endmodule 
module BLVDSIN (O, P_IN,N_IN);    // synthesis syn_black_box black_box_pad_pin="P_IN,N_IN"
input P_IN,N_IN; 
output O; 
endmodule 
module BLVDSOUT (P_OUT,N_OUT, I);    // synthesis syn_black_box black_box_pad_pin="P_OUT,N_OUT"
input I; 
output P_OUT,N_OUT; 
endmodule 
module BLVDSTRI (P_OUT,N_OUT, I,OE);    // synthesis syn_black_box black_box_pad_pin="P_OUT,N_OUT"
input I,OE; 
output P_OUT,N_OUT; 
endmodule 
module BLVDSIO (O, P_IO, N_IO, I, OE);    // synthesis syn_black_box black_box_pad_pin="P_IO,N_IO"
input I,OE; 
inout P_IO,N_IO; 
output O;
endmodule 
module CCU_AGB (COUT,A0,B0,CIN);   // synthesis syn_black_box
input A0,B0,CIN; 
output COUT; 
endmodule 
module CCU_AS (S0,COUT,A0,B0,CIN,AS);   // synthesis syn_black_box
input A0,B0,CIN,AS; 
output S0,COUT; 
endmodule 
module CCU_ADD (S0,COUT,A0,B0,CIN);   // synthesis syn_black_box
input A0,B0,CIN; 
output S0,COUT; 
endmodule 
module CCU_SUB (S0,COUT,A0,B0,CIN);   // synthesis syn_black_box
input A0,B0,CIN; 
output S0,COUT; 
endmodule 
module CCU_UDCP (S0,COUT,D, SD, LOAD, UD, CIN);  // synthesis syn_black_box
input D, SD, LOAD, UD, CIN ;
output S0,COUT; 
endmodule 
module CCU_UDC (S0,COUT, D, UD,CIN);   // synthesis syn_black_box
input D, UD, CIN; 
output S0,COUT; 
endmodule 
module CCU_DC (S0,COUT, D, CIN);   // synthesis syn_black_box
input D, CIN; 
output S0,COUT; 
endmodule 
module CCU_UC (S0,COUT, D, CIN);   // synthesis syn_black_box
input D, CIN; 
output S0,COUT; 
endmodule 
module DC_LSB (S0,COUT, D, CIN);   // synthesis syn_black_box
input D, CIN; 
output S0,COUT; 
endmodule 
module UC_LSB (S0,COUT, D, CIN);   // synthesis syn_black_box
input D, CIN; 
output S0,COUT; 
endmodule
module CCU_UCP (S0,COUT,D, SD, LOAD, CIN);  // synthesis syn_black_box
input D, SD, LOAD, CIN ;
output S0,COUT; 
endmodule
module CCU_DCP (S0,COUT,D, SD, LOAD, CIN);  // synthesis syn_black_box
input D, SD, LOAD, CIN ;
output S0,COUT; 
endmodule
//Memory Cells for ispMACH5000MX -- SuperCool
module RAMB16K_X1(CEN, CLK, WR, CS0, CS1, RST, DI0, AD0, AD1, AD2, AD3, AD4, AD5, AD6, AD7, AD8, AD9, AD10, AD11, AD12, AD13, DO0);// synthesis syn_black_box
input CEN;
input CLK;
input WR;
input CS0;
input CS1;
input RST;
input DI0;
input AD0;
input AD1;
input AD2;
input AD3;
input AD4;
input AD5;
input AD6;
input AD7;
input AD8;
input AD9;
input AD10;
input AD11;
input AD12;
input AD13;
output DO0;
endmodule 
module RAMB16K_X2(CEN, CLK, WR, CS0, CS1, RST, DI0, DI1, AD0, AD1, AD2, AD3, AD4, AD5, AD6, AD7, AD8, AD9, AD10, AD11, AD12, DO0, DO1);// synthesis syn_black_box
input CEN;
input CLK;
input WR;
input CS0;
input CS1;
input RST;
input DI0;
input DI1;
input AD0;
input AD1;
input AD2;
input AD3;
input AD4;
input AD5;
input AD6;
input AD7;
input AD8;
input AD9;
input AD10;
input AD11;
input AD12;
output DO0;
output DO1;
endmodule 
module RAMB16K_X4(CEN, CLK, WR, CS0, CS1, RST, DI0, DI1, DI2, DI3, AD0, AD1, AD2, AD3, AD4, AD5, AD6, AD7, AD8, AD9, AD10, AD11, DO0, DO1, DO2, DO3);// synthesis syn_black_box
input CEN;
input CLK;
input WR;
input CS0;
input CS1;
input RST;
input DI0;
input DI1;
input DI2;
input DI3;
input AD0;
input AD1;
input AD2;
input AD3;
input AD4;
input AD5;
input AD6;
input AD7;
input AD8;
input AD9;
input AD10;
input AD11;
output DO0;
output DO1;
output DO2;
output DO3;
endmodule 
module RAMB16K_X8(CEN, CLK, WR, CS0, CS1, RST, DI0, DI1, DI2, DI3, DI4, DI5, DI6, DI7, AD0, AD1, AD2, AD3, AD4, AD5, AD6, AD7, AD8, AD9, AD10, DO0, DO1, DO2, DO3, DO4, DO5, DO6, DO7);// synthesis syn_black_box
input CEN;
input CLK;
input WR;
input CS0;
input CS1;
input RST;
input DI0;
input DI1;
input DI2;
input DI3;
input DI4;
input DI5;
input DI6;
input DI7;
input AD0;
input AD1;
input AD2;
input AD3;
input AD4;
input AD5;
input AD6;
input AD7;
input AD8;
input AD9;
input AD10;
output DO0;
output DO1;
output DO2;
output DO3;
output DO4;
output DO5;
output DO6;
output DO7;
endmodule 
module RAMB16K_X16(CEN, CLK, WR, CS0, CS1, RST, DI0, DI1, DI2, DI3, DI4, DI5, DI6, DI7, DI8, DI9, DI10, DI11, DI12, DI13, DI14, DI15, AD0, AD1, AD2, AD3, AD4, AD5, AD6, AD7, AD8, AD9, DO0, DO1, DO2, DO3, DO4, DO5, DO6, DO7, DO8, DO9, DO10, DO11, DO12, DO13, DO14, DO15);// synthesis syn_black_box
input CEN;
input CLK;
input WR;
input CS0;
input CS1;
input RST;
input DI0;
input DI1;
input DI2;
input DI3;
input DI4;
input DI5;
input DI6;
input DI7;
input DI8;
input DI9;
input DI10;
input DI11;
input DI12;
input DI13;
input DI14;
input DI15;
input AD0;
input AD1;
input AD2;
input AD3;
input AD4;
input AD5;
input AD6;
input AD7;
input AD8;
input AD9;
output DO0;
output DO1;
output DO2;
output DO3;
output DO4;
output DO5;
output DO6;
output DO7;
output DO8;
output DO9;
output DO10;
output DO11;
output DO12;
output DO13;
output DO14;
output DO15;
endmodule 
module RAMB16K_X32(CEN, CLK, WR, CS0, CS1, RST, DI0, DI1, DI2, DI3, DI4, DI5, DI6, DI7, DI8, DI9, DI10, DI11, DI12, DI13, DI14, DI15, DI16, DI17, DI18, DI19, DI20, DI21, DI22, DI23, DI24, DI25, DI26, DI27, DI28, DI29, DI30, DI31, AD0, AD1, AD2, AD3, AD4, AD5, AD6, AD7, AD8, DO0, DO1, DO2, DO3, DO4, DO5, DO6, DO7, DO8, DO9, DO10, DO11, DO12, DO13, DO14, DO15, DO16, DO17, DO18, DO19, DO20, DO21, DO22, DO23, DO24, DO25, DO26, DO27, DO28, DO29, DO30, DO31);// synthesis syn_black_box
input CEN;
input CLK;
input WR;
input CS0;
input CS1;
input RST;
input DI0;
input DI1;
input DI2;
input DI3;
input DI4;
input DI5;
input DI6;
input DI7;
input DI8;
input DI9;
input DI10;
input DI11;
input DI12;
input DI13;
input DI14;
input DI15;
input DI16;
input DI17;
input DI18;
input DI19;
input DI20;
input DI21;
input DI22;
input DI23;
input DI24;
input DI25;
input DI26;
input DI27;
input DI28;
input DI29;
input DI30;
input DI31;
input AD0;
input AD1;
input AD2;
input AD3;
input AD4;
input AD5;
input AD6;
input AD7;
input AD8;
output DO0;
output DO1;
output DO2;
output DO3;
output DO4;
output DO5;
output DO6;
output DO7;
output DO8;
output DO9;
output DO10;
output DO11;
output DO12;
output DO13;
output DO14;
output DO15;
output DO16;
output DO17;
output DO18;
output DO19;
output DO20;
output DO21;
output DO22;
output DO23;
output DO24;
output DO25;
output DO26;
output DO27;
output DO28;
output DO29;
output DO30;
output DO31;
endmodule 
module RAMB16K_RX1_WX1(WCEN, WCLK, WCS0, WCS1, WE, RCEN, RCLK, RST, WD0, WAD0, WAD1, WAD2, WAD3, WAD4, WAD5, WAD6, WAD7, WAD8, WAD9, WAD10, WAD11, WAD12, WAD13, RAD0, RAD1, RAD2, RAD3, RAD4, RAD5, RAD6, RAD7, RAD8, RAD9, RAD10, RAD11, RAD12, RAD13, RD0);// synthesis syn_black_box
input WCEN;
input WCLK;
input WCS0;
input WCS1;
input WE;
input RCEN;
input RCLK;
input RST;
input WD0;
input WAD0;
input WAD1;
input WAD2;
input WAD3;
input WAD4;
input WAD5;
input WAD6;
input WAD7;
input WAD8;
input WAD9;
input WAD10;
input WAD11;
input WAD12;
input WAD13;
input RAD0;
input RAD1;
input RAD2;
input RAD3;
input RAD4;
input RAD5;
input RAD6;
input RAD7;
input RAD8;
input RAD9;
input RAD10;
input RAD11;
input RAD12;
input RAD13;
output RD0;
endmodule 
module RAMB16K_RX1_WX2(WCEN, WCLK, WCS0, WCS1, WE, RCEN, RCLK, RST, WD0, WAD0, WAD1, WAD2, WAD3, WAD4, WAD5, WAD6, WAD7, WAD8, WAD9, WAD10, WAD11, WAD12, WAD13, RAD0, RAD1, RAD2, RAD3, RAD4, RAD5, RAD6, RAD7, RAD8, RAD9, RAD10, RAD11, RAD12, RD0, RD1);// synthesis syn_black_box
input WCEN;
input WCLK;
input WCS0;
input WCS1;
input WE;
input RCEN;
input RCLK;
input RST;
input WD0;
input WAD0;
input WAD1;
input WAD2;
input WAD3;
input WAD4;
input WAD5;
input WAD6;
input WAD7;
input WAD8;
input WAD9;
input WAD10;
input WAD11;
input WAD12;
input WAD13;
input RAD0;
input RAD1;
input RAD2;
input RAD3;
input RAD4;
input RAD5;
input RAD6;
input RAD7;
input RAD8;
input RAD9;
input RAD10;
input RAD11;
input RAD12;
output RD0;
output RD1;
endmodule 
module RAMB16K_RX1_WX4(WCEN, WCLK, WCS0, WCS1, WE, RCEN, RCLK, RST, WD0, WAD0, WAD1, WAD2, WAD3, WAD4, WAD5, WAD6, WAD7, WAD8, WAD9, WAD10, WAD11, WAD12, WAD13, RAD0, RAD1, RAD2, RAD3, RAD4, RAD5, RAD6, RAD7, RAD8, RAD9, RAD10, RAD11, RD0, RD1, RD2, RD3);// synthesis syn_black_box
input WCEN;
input WCLK;
input WCS0;
input WCS1;
input WE;
input RCEN;
input RCLK;
input RST;
input WD0;
input WAD0;
input WAD1;
input WAD2;
input WAD3;
input WAD4;
input WAD5;
input WAD6;
input WAD7;
input WAD8;
input WAD9;
input WAD10;
input WAD11;
input WAD12;
input WAD13;
input RAD0;
input RAD1;
input RAD2;
input RAD3;
input RAD4;
input RAD5;
input RAD6;
input RAD7;
input RAD8;
input RAD9;
input RAD10;
input RAD11;
output RD0;
output RD1;
output RD2;
output RD3;
endmodule 
module RAMB16K_RX1_WX8(WCEN, WCLK, WCS0, WCS1, WE, RCEN, RCLK, RST, WD0, WAD0, WAD1, WAD2, WAD3, WAD4, WAD5, WAD6, WAD7, WAD8, WAD9, WAD10, WAD11, WAD12, WAD13, RAD0, RAD1, RAD2, RAD3, RAD4, RAD5, RAD6, RAD7, RAD8, RAD9, RAD10, RD0, RD1, RD2, RD3, RD4, RD5, RD6, RD7);// synthesis syn_black_box
input WCEN;
input WCLK;
input WCS0;
input WCS1;
input WE;
input RCEN;
input RCLK;
input RST;
input WD0;
input WAD0;
input WAD1;
input WAD2;
input WAD3;
input WAD4;
input WAD5;
input WAD6;
input WAD7;
input WAD8;
input WAD9;
input WAD10;
input WAD11;
input WAD12;
input WAD13;
input RAD0;
input RAD1;
input RAD2;
input RAD3;
input RAD4;
input RAD5;
input RAD6;
input RAD7;
input RAD8;
input RAD9;
input RAD10;
output RD0;
output RD1;
output RD2;
output RD3;
output RD4;
output RD5;
output RD6;
output RD7;
endmodule 
module RAMB16K_RX1_WX16(WCEN, WCLK, WCS0, WCS1, WE, RCEN, RCLK, RST, WD0, WAD0, WAD1, WAD2, WAD3, WAD4, WAD5, WAD6, WAD7, WAD8, WAD9, WAD10, WAD11, WAD12, WAD13, RAD0, RAD1, RAD2, RAD3, RAD4, RAD5, RAD6, RAD7, RAD8, RAD9, RD0, RD1, RD2, RD3, RD4, RD5, RD6, RD7, RD8, RD9, RD10, RD11, RD12, RD13, RD14, RD15);// synthesis syn_black_box
input WCEN;
input WCLK;
input WCS0;
input WCS1;
input WE;
input RCEN;
input RCLK;
input RST;
input WD0;
input WAD0;
input WAD1;
input WAD2;
input WAD3;
input WAD4;
input WAD5;
input WAD6;
input WAD7;
input WAD8;
input WAD9;
input WAD10;
input WAD11;
input WAD12;
input WAD13;
input RAD0;
input RAD1;
input RAD2;
input RAD3;
input RAD4;
input RAD5;
input RAD6;
input RAD7;
input RAD8;
input RAD9;
output RD0;
output RD1;
output RD2;
output RD3;
output RD4;
output RD5;
output RD6;
output RD7;
output RD8;
output RD9;
output RD10;
output RD11;
output RD12;
output RD13;
output RD14;
output RD15;
endmodule 
module RAMB16K_RX1_WX32(WCEN, WCLK, WCS0, WCS1, WE, RCEN, RCLK, RST, WD0, WAD0, WAD1, WAD2, WAD3, WAD4, WAD5, WAD6, WAD7, WAD8, WAD9, WAD10, WAD11, WAD12, WAD13, RAD0, RAD1, RAD2, RAD3, RAD4, RAD5, RAD6, RAD7, RAD8, RD0, RD1, RD2, RD3, RD4, RD5, RD6, RD7, RD8, RD9, RD10, RD11, RD12, RD13, RD14, RD15, RD16, RD17, RD18, RD19, RD20, RD21, RD22, RD23, RD24, RD25, RD26, RD27, RD28, RD29, RD30, RD31);// synthesis syn_black_box
input WCEN;
input WCLK;
input WCS0;
input WCS1;
input WE;
input RCEN;
input RCLK;
input RST;
input WD0;
input WAD0;
input WAD1;
input WAD2;
input WAD3;
input WAD4;
input WAD5;
input WAD6;
input WAD7;
input WAD8;
input WAD9;
input WAD10;
input WAD11;
input WAD12;
input WAD13;
input RAD0;
input RAD1;
input RAD2;
input RAD3;
input RAD4;
input RAD5;
input RAD6;
input RAD7;
input RAD8;
output RD0;
output RD1;
output RD2;
output RD3;
output RD4;
output RD5;
output RD6;
output RD7;
output RD8;
output RD9;
output RD10;
output RD11;
output RD12;
output RD13;
output RD14;
output RD15;
output RD16;
output RD17;
output RD18;
output RD19;
output RD20;
output RD21;
output RD22;
output RD23;
output RD24;
output RD25;
output RD26;
output RD27;
output RD28;
output RD29;
output RD30;
output RD31;
endmodule 
module RAMB16K_RX2_WX2(WCEN, WCLK, WCS0, WCS1, WE, RCEN, RCLK, RST, WD0, WD1, WAD0, WAD1, WAD2, WAD3, WAD4, WAD5, WAD6, WAD7, WAD8, WAD9, WAD10, WAD11, WAD12, RAD0, RAD1, RAD2, RAD3, RAD4, RAD5, RAD6, RAD7, RAD8, RAD9, RAD10, RAD11, RAD12, RD0, RD1);// synthesis syn_black_box
input WCEN;
input WCLK;
input WCS0;
input WCS1;
input WE;
input RCEN;
input RCLK;
input RST;
input WD0;
input WD1;
input WAD0;
input WAD1;
input WAD2;
input WAD3;
input WAD4;
input WAD5;
input WAD6;
input WAD7;
input WAD8;
input WAD9;
input WAD10;
input WAD11;
input WAD12;
input RAD0;
input RAD1;
input RAD2;
input RAD3;
input RAD4;
input RAD5;
input RAD6;
input RAD7;
input RAD8;
input RAD9;
input RAD10;
input RAD11;
input RAD12;
output RD0;
output RD1;
endmodule 
module RAMB16K_RX2_WX4(WCEN, WCLK, WCS0, WCS1, WE, RCEN, RCLK, RST, WD0, WD1, WAD0, WAD1, WAD2, WAD3, WAD4, WAD5, WAD6, WAD7, WAD8, WAD9, WAD10, WAD11, WAD12, RAD0, RAD1, RAD2, RAD3, RAD4, RAD5, RAD6, RAD7, RAD8, RAD9, RAD10, RAD11, RD0, RD1, RD2, RD3);// synthesis syn_black_box
input WCEN;
input WCLK;
input WCS0;
input WCS1;
input WE;
input RCEN;
input RCLK;
input RST;
input WD0;
input WD1;
input WAD0;
input WAD1;
input WAD2;
input WAD3;
input WAD4;
input WAD5;
input WAD6;
input WAD7;
input WAD8;
input WAD9;
input WAD10;
input WAD11;
input WAD12;
input RAD0;
input RAD1;
input RAD2;
input RAD3;
input RAD4;
input RAD5;
input RAD6;
input RAD7;
input RAD8;
input RAD9;
input RAD10;
input RAD11;
output RD0;
output RD1;
output RD2;
output RD3;
endmodule 
module RAMB16K_RX2_WX8(WCEN, WCLK, WCS0, WCS1, WE, RCEN, RCLK, RST, WD0, WD1, WAD0, WAD1, WAD2, WAD3, WAD4, WAD5, WAD6, WAD7, WAD8, WAD9, WAD10, WAD11, WAD12, RAD0, RAD1, RAD2, RAD3, RAD4, RAD5, RAD6, RAD7, RAD8, RAD9, RAD10, RD0, RD1, RD2, RD3, RD4, RD5, RD6, RD7);// synthesis syn_black_box
input WCEN;
input WCLK;
input WCS0;
input WCS1;
input WE;
input RCEN;
input RCLK;
input RST;
input WD0;
input WD1;
input WAD0;
input WAD1;
input WAD2;
input WAD3;
input WAD4;
input WAD5;
input WAD6;
input WAD7;
input WAD8;
input WAD9;
input WAD10;
input WAD11;
input WAD12;
input RAD0;
input RAD1;
input RAD2;
input RAD3;
input RAD4;
input RAD5;
input RAD6;
input RAD7;
input RAD8;
input RAD9;
input RAD10;
output RD0;
output RD1;
output RD2;
output RD3;
output RD4;
output RD5;
output RD6;
output RD7;
endmodule 
module RAMB16K_RX2_WX16(WCEN, WCLK, WCS0, WCS1, WE, RCEN, RCLK, RST, WD0, WD1, WAD0, WAD1, WAD2, WAD3, WAD4, WAD5, WAD6, WAD7, WAD8, WAD9, WAD10, WAD11, WAD12, RAD0, RAD1, RAD2, RAD3, RAD4, RAD5, RAD6, RAD7, RAD8, RAD9, RD0, RD1, RD2, RD3, RD4, RD5, RD6, RD7, RD8, RD9, RD10, RD11, RD12, RD13, RD14, RD15);// synthesis syn_black_box
input WCEN;
input WCLK;
input WCS0;
input WCS1;
input WE;
input RCEN;
input RCLK;
input RST;
input WD0;
input WD1;
input WAD0;
input WAD1;
input WAD2;
input WAD3;
input WAD4;
input WAD5;
input WAD6;
input WAD7;
input WAD8;
input WAD9;
input WAD10;
input WAD11;
input WAD12;
input RAD0;
input RAD1;
input RAD2;
input RAD3;
input RAD4;
input RAD5;
input RAD6;
input RAD7;
input RAD8;
input RAD9;
output RD0;
output RD1;
output RD2;
output RD3;
output RD4;
output RD5;
output RD6;
output RD7;
output RD8;
output RD9;
output RD10;
output RD11;
output RD12;
output RD13;
output RD14;
output RD15;
endmodule 
module RAMB16K_RX2_WX32(WCEN, WCLK, WCS0, WCS1, WE, RCEN, RCLK, RST, WD0, WD1, WAD0, WAD1, WAD2, WAD3, WAD4, WAD5, WAD6, WAD7, WAD8, WAD9, WAD10, WAD11, WAD12, RAD0, RAD1, RAD2, RAD3, RAD4, RAD5, RAD6, RAD7, RAD8, RD0, RD1, RD2, RD3, RD4, RD5, RD6, RD7, RD8, RD9, RD10, RD11, RD12, RD13, RD14, RD15, RD16, RD17, RD18, RD19, RD20, RD21, RD22, RD23, RD24, RD25, RD26, RD27, RD28, RD29, RD30, RD31);// synthesis syn_black_box
input WCEN;
input WCLK;
input WCS0;
input WCS1;
input WE;
input RCEN;
input RCLK;
input RST;
input WD0;
input WD1;
input WAD0;
input WAD1;
input WAD2;
input WAD3;
input WAD4;
input WAD5;
input WAD6;
input WAD7;
input WAD8;
input WAD9;
input WAD10;
input WAD11;
input WAD12;
input RAD0;
input RAD1;
input RAD2;
input RAD3;
input RAD4;
input RAD5;
input RAD6;
input RAD7;
input RAD8;
output RD0;
output RD1;
output RD2;
output RD3;
output RD4;
output RD5;
output RD6;
output RD7;
output RD8;
output RD9;
output RD10;
output RD11;
output RD12;
output RD13;
output RD14;
output RD15;
output RD16;
output RD17;
output RD18;
output RD19;
output RD20;
output RD21;
output RD22;
output RD23;
output RD24;
output RD25;
output RD26;
output RD27;
output RD28;
output RD29;
output RD30;
output RD31;
endmodule 
module RAMB16K_RX4_WX4(WCEN, WCLK, WCS0, WCS1, WE, RCEN, RCLK, RST, WD0, WD1, WD2, WD3, WAD0, WAD1, WAD2, WAD3, WAD4, WAD5, WAD6, WAD7, WAD8, WAD9, WAD10, WAD11, RAD0, RAD1, RAD2, RAD3, RAD4, RAD5, RAD6, RAD7, RAD8, RAD9, RAD10, RAD11, RD0, RD1, RD2, RD3);// synthesis syn_black_box
input WCEN;
input WCLK;
input WCS0;
input WCS1;
input WE;
input RCEN;
input RCLK;
input RST;
input WD0;
input WD1;
input WD2;
input WD3;
input WAD0;
input WAD1;
input WAD2;
input WAD3;
input WAD4;
input WAD5;
input WAD6;
input WAD7;
input WAD8;
input WAD9;
input WAD10;
input WAD11;
input RAD0;
input RAD1;
input RAD2;
input RAD3;
input RAD4;
input RAD5;
input RAD6;
input RAD7;
input RAD8;
input RAD9;
input RAD10;
input RAD11;
output RD0;
output RD1;
output RD2;
output RD3;
endmodule 
module RAMB16K_RX4_WX8(WCEN, WCLK, WCS0, WCS1, WE, RCEN, RCLK, RST, WD0, WD1, WD2, WD3, WAD0, WAD1, WAD2, WAD3, WAD4, WAD5, WAD6, WAD7, WAD8, WAD9, WAD10, WAD11, RAD0, RAD1, RAD2, RAD3, RAD4, RAD5, RAD6, RAD7, RAD8, RAD9, RAD10, RD0, RD1, RD2, RD3, RD4, RD5, RD6, RD7);// synthesis syn_black_box
input WCEN;
input WCLK;
input WCS0;
input WCS1;
input WE;
input RCEN;
input RCLK;
input RST;
input WD0;
input WD1;
input WD2;
input WD3;
input WAD0;
input WAD1;
input WAD2;
input WAD3;
input WAD4;
input WAD5;
input WAD6;
input WAD7;
input WAD8;
input WAD9;
input WAD10;
input WAD11;
input RAD0;
input RAD1;
input RAD2;
input RAD3;
input RAD4;
input RAD5;
input RAD6;
input RAD7;
input RAD8;
input RAD9;
input RAD10;
output RD0;
output RD1;
output RD2;
output RD3;
output RD4;
output RD5;
output RD6;
output RD7;
endmodule 
//////////////////////////
module RAMB16K_RX4_WX16(WCEN, WCLK, WCS0, WCS1, WE, RCEN, RCLK, RST, WD0, WD1, WD2, WD3, WAD0, WAD1, WAD2, WAD3, WAD4, WAD5, WAD6, WAD7, WAD8, WAD9, WAD10, WAD11, RAD0, RAD1, RAD2, RAD3, RAD4, RAD5, RAD6, RAD7, RAD8, RAD9, RD0, RD1, RD2, RD3, RD4, RD5, RD6, RD7, RD8, RD9, RD10, RD11, RD12, RD13, RD14, RD15);// synthesis syn_black_box
input WCEN;
input WCLK;
input WCS0;
input WCS1;
input WE;
input RCEN;
input RCLK;
input RST;
input WD0;
input WD1;
input WD2;
input WD3;
input WAD0;
input WAD1;
input WAD2;
input WAD3;
input WAD4;
input WAD5;
input WAD6;
input WAD7;
input WAD8;
input WAD9;
input WAD10;
input WAD11;
input RAD0;
input RAD1;
input RAD2;
input RAD3;
input RAD4;
input RAD5;
input RAD6;
input RAD7;
input RAD8;
input RAD9;
output RD0;
output RD1;
output RD2;
output RD3;
output RD4;
output RD5;
output RD6;
output RD7;
output RD8;
output RD9;
output RD10;
output RD11;
output RD12;
output RD13;
output RD14;
output RD15;
endmodule
module RAMB16K_RX4_WX32(WCEN, WCLK, WCS0, WCS1, WE, RCEN, RCLK, RST, WD0, WD1, WD2, WD3, WAD0, WAD1, WAD2, WAD3, WAD4, WAD5, WAD6, WAD7, WAD8, WAD9, WAD10, WAD11, RAD0, RAD1, RAD2, RAD3, RAD4, RAD5, RAD6, RAD7, RAD8, RD0, RD1, RD2, RD3, RD4, RD5, RD6, RD7, RD8, RD9, RD10, RD11, RD12, RD13, RD14, RD15, RD16, RD17, RD18, RD19, RD20, RD21, RD22, RD23, RD24, RD25, RD26, RD27, RD28, RD29, RD30, RD31);// synthesis syn_black_box
input WCEN;
input WCLK;
input WCS0;
input WCS1;
input WE;
input RCEN;
input RCLK;
input RST;
input WD0;
input WD1;
input WD2;
input WD3;
input WAD0;
input WAD1;
input WAD2;
input WAD3;
input WAD4;
input WAD5;
input WAD6;
input WAD7;
input WAD8;
input WAD9;
input WAD10;
input WAD11;
input RAD0;
input RAD1;
input RAD2;
input RAD3;
input RAD4;
input RAD5;
input RAD6;
input RAD7;
input RAD8;
output RD0;
output RD1;
output RD2;
output RD3;
output RD4;
output RD5;
output RD6;
output RD7;
output RD8;
output RD9;
output RD10;
output RD11;
output RD12;
output RD13;
output RD14;
output RD15;
output RD16;
output RD17;
output RD18;
output RD19;
output RD20;
output RD21;
output RD22;
output RD23;
output RD24;
output RD25;
output RD26;
output RD27;
output RD28;
output RD29;
output RD30;
output RD31;
endmodule  
module RAMB16K_RX8_WX8(WCEN, WCLK, WCS0, WCS1, WE, RCEN, RCLK, RST, WD0, WD1, WD2, WD3, WD4, WD5, WD6, WD7, WAD0, WAD1, WAD2, WAD3, WAD4, WAD5, WAD6, WAD7, WAD8, WAD9, WAD10, RAD0, RAD1, RAD2, RAD3, RAD4, RAD5, RAD6, RAD7, RAD8, RAD9, RAD10, RD0, RD1, RD2, RD3, RD4, RD5, RD6, RD7);// synthesis syn_black_box
input WCEN;
input WCLK;
input WCS0;
input WCS1;
input WE;
input RCEN;
input RCLK;
input RST;
input WD0;
input WD1;
input WD2;
input WD3;
input WD4;
input WD5;
input WD6;
input WD7;
input WAD0;
input WAD1;
input WAD2;
input WAD3;
input WAD4;
input WAD5;
input WAD6;
input WAD7;
input WAD8;
input WAD9;
input WAD10;
input RAD0;
input RAD1;
input RAD2;
input RAD3;
input RAD4;
input RAD5;
input RAD6;
input RAD7;
input RAD8;
input RAD9;
input RAD10;
output RD0;
output RD1;
output RD2;
output RD3;
output RD4;
output RD5;
output RD6;
output RD7;
endmodule 
module RAMB16K_RX8_WX16(WCEN, WCLK, WCS0, WCS1, WE, RCEN, RCLK, RST, WD0, WD1, WD2, WD3, WD4, WD5, WD6, WD7, WAD0, WAD1, WAD2, WAD3, WAD4, WAD5, WAD6, WAD7, WAD8, WAD9, WAD10, RAD0, RAD1, RAD2, RAD3, RAD4, RAD5, RAD6, RAD7, RAD8, RAD9, RD0, RD1, RD2, RD3, RD4, RD5, RD6, RD7, RD8, RD9, RD10, RD11, RD12, RD13, RD14, RD15);// synthesis syn_black_box
input WCEN;
input WCLK;
input WCS0;
input WCS1;
input WE;
input RCEN;
input RCLK;
input RST;
input WD0;
input WD1;
input WD2;
input WD3;
input WD4;
input WD5;
input WD6;
input WD7;
input WAD0;
input WAD1;
input WAD2;
input WAD3;
input WAD4;
input WAD5;
input WAD6;
input WAD7;
input WAD8;
input WAD9;
input WAD10;
input RAD0;
input RAD1;
input RAD2;
input RAD3;
input RAD4;
input RAD5;
input RAD6;
input RAD7;
input RAD8;
input RAD9;
output RD0;
output RD1;
output RD2;
output RD3;
output RD4;
output RD5;
output RD6;
output RD7;
output RD8;
output RD9;
output RD10;
output RD11;
output RD12;
output RD13;
output RD14;
output RD15;
endmodule
module RAMB16K_RX8_WX32(WCEN, WCLK, WCS0, WCS1, WE, RCEN, RCLK, RST, WD0, WD1, WD2, WD3, WD4, WD5, WD6, WD7, WAD0, WAD1, WAD2, WAD3, WAD4, WAD5, WAD6, WAD7, WAD8, WAD9, WAD10, RAD0, RAD1, RAD2, RAD3, RAD4, RAD5, RAD6, RAD7, RAD8, RD0, RD1, RD2, RD3, RD4, RD5, RD6, RD7, RD8, RD9, RD10, RD11, RD12, RD13, RD14, RD15, RD16, RD17, RD18, RD19, RD20, RD21, RD22, RD23, RD24, RD25, RD26, RD27, RD28, RD29, RD30, RD31);// synthesis syn_black_box
input WCEN;
input WCLK;
input WCS0;
input WCS1;
input WE;
input RCEN;
input RCLK;
input RST;
input WD0;
input WD1;
input WD2;
input WD3;
input WD4;
input WD5;
input WD6;
input WD7;
input WAD0;
input WAD1;
input WAD2;
input WAD3;
input WAD4;
input WAD5;
input WAD6;
input WAD7;
input WAD8;
input WAD9;
input WAD10;
input RAD0;
input RAD1;
input RAD2;
input RAD3;
input RAD4;
input RAD5;
input RAD6;
input RAD7;
input RAD8;
output RD0;
output RD1;
output RD2;
output RD3;
output RD4;
output RD5;
output RD6;
output RD7;
output RD8;
output RD9;
output RD10;
output RD11;
output RD12;
output RD13;
output RD14;
output RD15;
output RD16;
output RD17;
output RD18;
output RD19;
output RD20;
output RD21;
output RD22;
output RD23;
output RD24;
output RD25;
output RD26;
output RD27;
output RD28;
output RD29;
output RD30;
output RD31;
endmodule  
module RAMB16K_RX16_WX16(WCEN, WCLK, WCS0, WCS1, WE, RCEN, RCLK, RST, WD0, WD1, WD2, WD3, WD4, WD5, WD6, WD7, WD8, WD9, WD10, WD11, WD12, WD13, WD14, WD15, WAD0, WAD1, WAD2, WAD3, WAD4, WAD5, WAD6, WAD7, WAD8, WAD9, RAD0, RAD1, RAD2, RAD3, RAD4, RAD5, RAD6, RAD7, RAD8, RAD9, RD0, RD1, RD2, RD3, RD4, RD5, RD6, RD7, RD8, RD9, RD10, RD11, RD12, RD13, RD14, RD15);// synthesis syn_black_box
input WCEN;
input WCLK;
input WCS0;
input WCS1;
input WE;
input RCEN;
input RCLK;
input RST;
input WD0;
input WD1;
input WD2;
input WD3;
input WD4;
input WD5;
input WD6;
input WD7;
input WD8;
input WD9;
input WD10;
input WD11;
input WD12;
input WD13;
input WD14;
input WD15;
input WAD0;
input WAD1;
input WAD2;
input WAD3;
input WAD4;
input WAD5;
input WAD6;
input WAD7;
input WAD8;
input WAD9;
input RAD0;
input RAD1;
input RAD2;
input RAD3;
input RAD4;
input RAD5;
input RAD6;
input RAD7;
input RAD8;
input RAD9;
output RD0;
output RD1;
output RD2;
output RD3;
output RD4;
output RD5;
output RD6;
output RD7;
output RD8;
output RD9;
output RD10;
output RD11;
output RD12;
output RD13;
output RD14;
output RD15;
endmodule
module RAMB16K_RX16_WX32(WCEN, WCLK, WCS0, WCS1, WE, RCEN, RCLK, RST, WD0, WD1, WD2, WD3, WD4, WD5, WD6, WD7, WD8, WD9, WD10, WD11, WD12, WD13, WD14, WD15, WAD0, WAD1, WAD2, WAD3, WAD4, WAD5, WAD6, WAD7, WAD8, WAD9, RAD0, RAD1, RAD2, RAD3, RAD4, RAD5, RAD6, RAD7, RAD8, RD0, RD1, RD2, RD3, RD4, RD5, RD6, RD7, RD8, RD9, RD10, RD11, RD12, RD13, RD14, RD15, RD16, RD17, RD18, RD19, RD20, RD21, RD22, RD23, RD24, RD25, RD26, RD27, RD28, RD29, RD30, RD31);// synthesis syn_black_box
input WCEN;
input WCLK;
input WCS0;
input WCS1;
input WE;
input RCEN;
input RCLK;
input RST;
input WD0;
input WD1;
input WD2;
input WD3;
input WD4;
input WD5;
input WD6;
input WD7;
input WD8;
input WD9;
input WD10;
input WD11;
input WD12;
input WD13;
input WD14;
input WD15;
input WAD0;
input WAD1;
input WAD2;
input WAD3;
input WAD4;
input WAD5;
input WAD6;
input WAD7;
input WAD8;
input WAD9;
input RAD0;
input RAD1;
input RAD2;
input RAD3;
input RAD4;
input RAD5;
input RAD6;
input RAD7;
input RAD8;
output RD0;
output RD1;
output RD2;
output RD3;
output RD4;
output RD5;
output RD6;
output RD7;
output RD8;
output RD9;
output RD10;
output RD11;
output RD12;
output RD13;
output RD14;
output RD15;
output RD16;
output RD17;
output RD18;
output RD19;
output RD20;
output RD21;
output RD22;
output RD23;
output RD24;
output RD25;
output RD26;
output RD27;
output RD28;
output RD29;
output RD30;
output RD31;
endmodule  
module RAMB16K_RX32_WX32(WCEN, WCLK, WCS0, WCS1, WE, RCEN, RCLK, RST, WD0, WD1, WD2, WD3, WD4, WD5, WD6, WD7, WD8, WD9, WD10, WD11, WD12, WD13, WD14, WD15, WD16, WD17, WD18, WD19, WD20, WD21, WD22, WD23, WD24, WD25, WD26, WD27, WD28, WD29, WD30, WD31, WAD0, WAD1, WAD2, WAD3, WAD4, WAD5, WAD6, WAD7, WAD8, RAD0, RAD1, RAD2, RAD3, RAD4, RAD5, RAD6, RAD7, RAD8, RD0, RD1, RD2, RD3, RD4, RD5, RD6, RD7, RD8, RD9, RD10, RD11, RD12, RD13, RD14, RD15, RD16, RD17, RD18, RD19, RD20, RD21, RD22, RD23, RD24, RD25, RD26, RD27, RD28, RD29, RD30, RD31);// synthesis syn_black_box
input WCEN;
input WCLK;
input WCS0;
input WCS1;
input WE;
input RCEN;
input RCLK;
input RST;
input WD0;
input WD1;
input WD2;
input WD3;
input WD4;
input WD5;
input WD6;
input WD7;
input WD8;
input WD9;
input WD10;
input WD11;
input WD12;
input WD13;
input WD14;
input WD15;
input WD16;
input WD17;
input WD18;
input WD19;
input WD20;
input WD21;
input WD22;
input WD23;
input WD24;
input WD25;
input WD26;
input WD27;
input WD28;
input WD29;
input WD30;
input WD31;
input WAD0;
input WAD1;
input WAD2;
input WAD3;
input WAD4;
input WAD5;
input WAD6;
input WAD7;
input WAD8;
input RAD0;
input RAD1;
input RAD2;
input RAD3;
input RAD4;
input RAD5;
input RAD6;
input RAD7;
input RAD8;
output RD0;
output RD1;
output RD2;
output RD3;
output RD4;
output RD5;
output RD6;
output RD7;
output RD8;
output RD9;
output RD10;
output RD11;
output RD12;
output RD13;
output RD14;
output RD15;
output RD16;
output RD17;
output RD18;
output RD19;
output RD20;
output RD21;
output RD22;
output RD23;
output RD24;
output RD25;
output RD26;
output RD27;
output RD28;
output RD29;
output RD30;
output RD31;
endmodule  
module RAMB8K_X1_X1(CENA, CLKA, WRA, CSA0, CSA1, RSTA, CENB, CLKB, WRB, CSB0, CSB1, RSTB, DIA0, ADA0, ADA1, ADA2, ADA3, ADA4, ADA5, ADA6, ADA7, ADA8, ADA9, ADA10, ADA11, ADA12, DIB0, ADB0, ADB1, ADB2, ADB3, ADB4, ADB5, ADB6, ADB7, ADB8, ADB9, ADB10, ADB11, ADB12, DOA0, DOB0);// synthesis syn_black_box
input CENA;
input CLKA;
input WRA;
input CSA0;
input CSA1;
input RSTA;
input CENB;
input CLKB;
input WRB;
input CSB0;
input CSB1;
input RSTB;
input DIA0;
input ADA0;
input ADA1;
input ADA2;
input ADA3;
input ADA4;
input ADA5;
input ADA6;
input ADA7;
input ADA8;
input ADA9;
input ADA10;
input ADA11;
input ADA12;
input DIB0;
input ADB0;
input ADB1;
input ADB2;
input ADB3;
input ADB4;
input ADB5;
input ADB6;
input ADB7;
input ADB8;
input ADB9;
input ADB10;
input ADB11;
input ADB12;
output DOA0;
output DOB0;
endmodule 
module RAMB8K_X1_X2(CENA, CLKA, WRA, CSA0, CSA1, RSTA, CENB, CLKB, WRB, CSB0, CSB1, RSTB, DIA0, ADA0, ADA1, ADA2, ADA3, ADA4, ADA5, ADA6, ADA7, ADA8, ADA9, ADA10, ADA11, ADA12, DIB0, DIB1, ADB0, ADB1, ADB2, ADB3, ADB4, ADB5, ADB6, ADB7, ADB8, ADB9, ADB10, ADB11, DOA0, DOB0, DOB1);// synthesis syn_black_box
input CENA;
input CLKA;
input WRA;
input CSA0;
input CSA1;
input RSTA;
input CENB;
input CLKB;
input WRB;
input CSB0;
input CSB1;
input RSTB;
input DIA0;
input ADA0;
input ADA1;
input ADA2;
input ADA3;
input ADA4;
input ADA5;
input ADA6;
input ADA7;
input ADA8;
input ADA9;
input ADA10;
input ADA11;
input ADA12;
input DIB0;
input DIB1;
input ADB0;
input ADB1;
input ADB2;
input ADB3;
input ADB4;
input ADB5;
input ADB6;
input ADB7;
input ADB8;
input ADB9;
input ADB10;
input ADB11;
output DOA0;
output DOB0;
output DOB1;
endmodule 
module RAMB8K_X1_X4(CENA, CLKA, WRA, CSA0, CSA1, RSTA, CENB, CLKB, WRB, CSB0, CSB1, RSTB, DIA0, ADA0, ADA1, ADA2, ADA3, ADA4, ADA5, ADA6, ADA7, ADA8, ADA9, ADA10, ADA11, ADA12, DIB0, DIB1, DIB2, DIB3, ADB0, ADB1, ADB2, ADB3, ADB4, ADB5, ADB6, ADB7, ADB8, ADB9, ADB10, DOA0, DOB0, DOB1, DOB2, DOB3);// synthesis syn_black_box
input CENA;
input CLKA;
input WRA;
input CSA0;
input CSA1;
input RSTA;
input CENB;
input CLKB;
input WRB;
input CSB0;
input CSB1;
input RSTB;
input DIA0;
input ADA0;
input ADA1;
input ADA2;
input ADA3;
input ADA4;
input ADA5;
input ADA6;
input ADA7;
input ADA8;
input ADA9;
input ADA10;
input ADA11;
input ADA12;
input DIB0;
input DIB1;
input DIB2;
input DIB3;
input ADB0;
input ADB1;
input ADB2;
input ADB3;
input ADB4;
input ADB5;
input ADB6;
input ADB7;
input ADB8;
input ADB9;
input ADB10;
output DOA0;
output DOB0;
output DOB1;
output DOB2;
output DOB3;
endmodule 
module RAMB8K_X1_X8(CENA, CLKA, WRA, CSA0, CSA1, RSTA, CENB, CLKB, WRB, CSB0, CSB1, RSTB, DIA0, ADA0, ADA1, ADA2, ADA3, ADA4, ADA5, ADA6, ADA7, ADA8, ADA9, ADA10, ADA11, ADA12, DIB0, DIB1, DIB2, DIB3, DIB4, DIB5, DIB6, DIB7, ADB0, ADB1, ADB2, ADB3, ADB4, ADB5, ADB6, ADB7, ADB8, ADB9, DOA0, DOB0, DOB1, DOB2, DOB3, DOB4, DOB5, DOB6, DOB7);// synthesis syn_black_box
input CENA;
input CLKA;
input WRA;
input CSA0;
input CSA1;
input RSTA;
input CENB;
input CLKB;
input WRB;
input CSB0;
input CSB1;
input RSTB;
input DIA0;
input ADA0;
input ADA1;
input ADA2;
input ADA3;
input ADA4;
input ADA5;
input ADA6;
input ADA7;
input ADA8;
input ADA9;
input ADA10;
input ADA11;
input ADA12;
input DIB0;
input DIB1;
input DIB2;
input DIB3;
input DIB4;
input DIB5;
input DIB6;
input DIB7;
input ADB0;
input ADB1;
input ADB2;
input ADB3;
input ADB4;
input ADB5;
input ADB6;
input ADB7;
input ADB8;
input ADB9;
output DOA0;
output DOB0;
output DOB1;
output DOB2;
output DOB3;
output DOB4;
output DOB5;
output DOB6;
output DOB7;
endmodule 
module RAMB8K_X1_X16(CENA, CLKA, WRA, CSA0, CSA1, RSTA, CENB, CLKB, WRB, CSB0, CSB1, RSTB, DIA0, ADA0, ADA1, ADA2, ADA3, ADA4, ADA5, ADA6, ADA7, ADA8, ADA9, ADA10, ADA11, ADA12, DIB0, DIB1, DIB2, DIB3, DIB4, DIB5, DIB6, DIB7, DIB8, DIB9, DIB10, DIB11, DIB12, DIB13, DIB14, DIB15, ADB0, ADB1, ADB2, ADB3, ADB4, ADB5, ADB6, ADB7, ADB8, DOA0, DOB0, DOB1, DOB2, DOB3, DOB4, DOB5, DOB6, DOB7, DOB8, DOB9, DOB10, DOB11, DOB12, DOB13, DOB14, DOB15);// synthesis syn_black_box
input CENA;
input CLKA;
input WRA;
input CSA0;
input CSA1;
input RSTA;
input CENB;
input CLKB;
input WRB;
input CSB0;
input CSB1;
input RSTB;
input DIA0;
input ADA0;
input ADA1;
input ADA2;
input ADA3;
input ADA4;
input ADA5;
input ADA6;
input ADA7;
input ADA8;
input ADA9;
input ADA10;
input ADA11;
input ADA12;
input DIB0;
input DIB1;
input DIB2;
input DIB3;
input DIB4;
input DIB5;
input DIB6;
input DIB7;
input DIB8;
input DIB9;
input DIB10;
input DIB11;
input DIB12;
input DIB13;
input DIB14;
input DIB15;
input ADB0;
input ADB1;
input ADB2;
input ADB3;
input ADB4;
input ADB5;
input ADB6;
input ADB7;
input ADB8;
output DOA0;
output DOB0;
output DOB1;
output DOB2;
output DOB3;
output DOB4;
output DOB5;
output DOB6;
output DOB7;
output DOB8;
output DOB9;
output DOB10;
output DOB11;
output DOB12;
output DOB13;
output DOB14;
output DOB15;
endmodule 
module RAMB8K_X2_X2(CENA, CLKA, WRA, CSA0, CSA1, RSTA, CENB, CLKB, WRB, CSB0, CSB1, RSTB, DIA0, DIA1, ADA0, ADA1, ADA2, ADA3, ADA4, ADA5, ADA6, ADA7, ADA8, ADA9, ADA10, ADA11, DIB0, DIB1, ADB0, ADB1, ADB2, ADB3, ADB4, ADB5, ADB6, ADB7, ADB8, ADB9, ADB10, ADB11, DOA0, DOA1, DOB0, DOB1);// synthesis syn_black_box
input CENA;
input CLKA;
input WRA;
input CSA0;
input CSA1;
input RSTA;
input CENB;
input CLKB;
input WRB;
input CSB0;
input CSB1;
input RSTB;
input DIA0;
input DIA1;
input ADA0;
input ADA1;
input ADA2;
input ADA3;
input ADA4;
input ADA5;
input ADA6;
input ADA7;
input ADA8;
input ADA9;
input ADA10;
input ADA11;
input DIB0;
input DIB1;
input ADB0;
input ADB1;
input ADB2;
input ADB3;
input ADB4;
input ADB5;
input ADB6;
input ADB7;
input ADB8;
input ADB9;
input ADB10;
input ADB11;
output DOA0;
output DOA1;
output DOB0;
output DOB1;
endmodule 
module RAMB8K_X2_X4(CENA, CLKA, WRA, CSA0, CSA1, RSTA, CENB, CLKB, WRB, CSB0, CSB1, RSTB, DIA0, DIA1, ADA0, ADA1, ADA2, ADA3, ADA4, ADA5, ADA6, ADA7, ADA8, ADA9, ADA10, ADA11, DIB0, DIB1, DIB2, DIB3, ADB0, ADB1, ADB2, ADB3, ADB4, ADB5, ADB6, ADB7, ADB8, ADB9, ADB10, DOA0, DOA1, DOB0, DOB1, DOB2, DOB3);// synthesis syn_black_box
input CENA;
input CLKA;
input WRA;
input CSA0;
input CSA1;
input RSTA;
input CENB;
input CLKB;
input WRB;
input CSB0;
input CSB1;
input RSTB;
input DIA0;
input DIA1;
input ADA0;
input ADA1;
input ADA2;
input ADA3;
input ADA4;
input ADA5;
input ADA6;
input ADA7;
input ADA8;
input ADA9;
input ADA10;
input ADA11;
input DIB0;
input DIB1;
input DIB2;
input DIB3;
input ADB0;
input ADB1;
input ADB2;
input ADB3;
input ADB4;
input ADB5;
input ADB6;
input ADB7;
input ADB8;
input ADB9;
input ADB10;
output DOA0;
output DOA1;
output DOB0;
output DOB1;
output DOB2;
output DOB3;
endmodule 
module RAMB8K_X2_X8(CENA, CLKA, WRA, CSA0, CSA1, RSTA, CENB, CLKB, WRB, CSB0, CSB1, RSTB, DIA0, DIA1, ADA0, ADA1, ADA2, ADA3, ADA4, ADA5, ADA6, ADA7, ADA8, ADA9, ADA10, ADA11, DIB0, DIB1, DIB2, DIB3, DIB4, DIB5, DIB6, DIB7, ADB0, ADB1, ADB2, ADB3, ADB4, ADB5, ADB6, ADB7, ADB8, ADB9, DOA0, DOA1, DOB0, DOB1, DOB2, DOB3, DOB4, DOB5, DOB6, DOB7);// synthesis syn_black_box
input CENA;
input CLKA;
input WRA;
input CSA0;
input CSA1;
input RSTA;
input CENB;
input CLKB;
input WRB;
input CSB0;
input CSB1;
input RSTB;
input DIA0;
input DIA1;
input ADA0;
input ADA1;
input ADA2;
input ADA3;
input ADA4;
input ADA5;
input ADA6;
input ADA7;
input ADA8;
input ADA9;
input ADA10;
input ADA11;
input DIB0;
input DIB1;
input DIB2;
input DIB3;
input DIB4;
input DIB5;
input DIB6;
input DIB7;
input ADB0;
input ADB1;
input ADB2;
input ADB3;
input ADB4;
input ADB5;
input ADB6;
input ADB7;
input ADB8;
input ADB9;
output DOA0;
output DOA1;
output DOB0;
output DOB1;
output DOB2;
output DOB3;
output DOB4;
output DOB5;
output DOB6;
output DOB7;
endmodule 
module RAMB8K_X2_X16(CENA, CLKA, WRA, CSA0, CSA1, RSTA, CENB, CLKB, WRB, CSB0, CSB1, RSTB, DIA0, DIA1, ADA0, ADA1, ADA2, ADA3, ADA4, ADA5, ADA6, ADA7, ADA8, ADA9, ADA10, ADA11, DIB0, DIB1, DIB2, DIB3, DIB4, DIB5, DIB6, DIB7, DIB8, DIB9, DIB10, DIB11, DIB12, DIB13, DIB14, DIB15, ADB0, ADB1, ADB2, ADB3, ADB4, ADB5, ADB6, ADB7, ADB8, DOA0, DOA1, DOB0, DOB1, DOB2, DOB3, DOB4, DOB5, DOB6, DOB7, DOB8, DOB9, DOB10, DOB11, DOB12, DOB13, DOB14, DOB15);// synthesis syn_black_box
input CENA;
input CLKA;
input WRA;
input CSA0;
input CSA1;
input RSTA;
input CENB;
input CLKB;
input WRB;
input CSB0;
input CSB1;
input RSTB;
input DIA0;
input DIA1;
input ADA0;
input ADA1;
input ADA2;
input ADA3;
input ADA4;
input ADA5;
input ADA6;
input ADA7;
input ADA8;
input ADA9;
input ADA10;
input ADA11;
input DIB0;
input DIB1;
input DIB2;
input DIB3;
input DIB4;
input DIB5;
input DIB6;
input DIB7;
input DIB8;
input DIB9;
input DIB10;
input DIB11;
input DIB12;
input DIB13;
input DIB14;
input DIB15;
input ADB0;
input ADB1;
input ADB2;
input ADB3;
input ADB4;
input ADB5;
input ADB6;
input ADB7;
input ADB8;
output DOA0;
output DOA1;
output DOB0;
output DOB1;
output DOB2;
output DOB3;
output DOB4;
output DOB5;
output DOB6;
output DOB7;
output DOB8;
output DOB9;
output DOB10;
output DOB11;
output DOB12;
output DOB13;
output DOB14;
output DOB15;
endmodule 
module RAMB8K_X4_X4(CENA, CLKA, WRA, CSA0, CSA1, RSTA, CENB, CLKB, WRB, CSB0, CSB1, RSTB, DIA0, DIA1, DIA2, DIA3, ADA0, ADA1, ADA2, ADA3, ADA4, ADA5, ADA6, ADA7, ADA8, ADA9, ADA10, DIB0, DIB1, DIB2, DIB3, ADB0, ADB1, ADB2, ADB3, ADB4, ADB5, ADB6, ADB7, ADB8, ADB9, ADB10, DOA0, DOA1, DOA2, DOA3, DOB0, DOB1, DOB2, DOB3);// synthesis syn_black_box
input CENA;
input CLKA;
input WRA;
input CSA0;
input CSA1;
input RSTA;
input CENB;
input CLKB;
input WRB;
input CSB0;
input CSB1;
input RSTB;
input DIA0;
input DIA1;
input DIA2;
input DIA3;
input ADA0;
input ADA1;
input ADA2;
input ADA3;
input ADA4;
input ADA5;
input ADA6;
input ADA7;
input ADA8;
input ADA9;
input ADA10;
input DIB0;
input DIB1;
input DIB2;
input DIB3;
input ADB0;
input ADB1;
input ADB2;
input ADB3;
input ADB4;
input ADB5;
input ADB6;
input ADB7;
input ADB8;
input ADB9;
input ADB10;
output DOA0;
output DOA1;
output DOA2;
output DOA3;
output DOB0;
output DOB1;
output DOB2;
output DOB3;
endmodule 
module RAMB8K_X4_X8(CENA, CLKA, WRA, CSA0, CSA1, RSTA, CENB, CLKB, WRB, CSB0, CSB1, RSTB, DIA0, DIA1, DIA2, DIA3, ADA0, ADA1, ADA2, ADA3, ADA4, ADA5, ADA6, ADA7, ADA8, ADA9, ADA10, DIB0, DIB1, DIB2, DIB3, DIB4, DIB5, DIB6, DIB7, ADB0, ADB1, ADB2, ADB3, ADB4, ADB5, ADB6, ADB7, ADB8, ADB9, DOA0, DOA1, DOA2, DOA3, DOB0, DOB1, DOB2, DOB3, DOB4, DOB5, DOB6, DOB7);// synthesis syn_black_box
input CENA;
input CLKA;
input WRA;
input CSA0;
input CSA1;
input RSTA;
input CENB;
input CLKB;
input WRB;
input CSB0;
input CSB1;
input RSTB;
input DIA0;
input DIA1;
input DIA2;
input DIA3;
input ADA0;
input ADA1;
input ADA2;
input ADA3;
input ADA4;
input ADA5;
input ADA6;
input ADA7;
input ADA8;
input ADA9;
input ADA10;
input DIB0;
input DIB1;
input DIB2;
input DIB3;
input DIB4;
input DIB5;
input DIB6;
input DIB7;
input ADB0;
input ADB1;
input ADB2;
input ADB3;
input ADB4;
input ADB5;
input ADB6;
input ADB7;
input ADB8;
input ADB9;
output DOA0;
output DOA1;
output DOA2;
output DOA3;
output DOB0;
output DOB1;
output DOB2;
output DOB3;
output DOB4;
output DOB5;
output DOB6;
output DOB7;
endmodule 
module RAMB8K_X4_X16(CENA, CLKA, WRA, CSA0, CSA1, RSTA, CENB, CLKB, WRB, CSB0, CSB1, RSTB, DIA0, DIA1, DIA2, DIA3, ADA0, ADA1, ADA2, ADA3, ADA4, ADA5, ADA6, ADA7, ADA8, ADA9, ADA10, DIB0, DIB1, DIB2, DIB3, DIB4, DIB5, DIB6, DIB7, DIB8, DIB9, DIB10, DIB11, DIB12, DIB13, DIB14, DIB15, ADB0, ADB1, ADB2, ADB3, ADB4, ADB5, ADB6, ADB7, ADB8, DOA0, DOA1, DOA2, DOA3, DOB0, DOB1, DOB2, DOB3, DOB4, DOB5, DOB6, DOB7, DOB8, DOB9, DOB10, DOB11, DOB12, DOB13, DOB14, DOB15);// synthesis syn_black_box
input CENA;
input CLKA;
input WRA;
input CSA0;
input CSA1;
input RSTA;
input CENB;
input CLKB;
input WRB;
input CSB0;
input CSB1;
input RSTB;
input DIA0;
input DIA1;
input DIA2;
input DIA3;
input ADA0;
input ADA1;
input ADA2;
input ADA3;
input ADA4;
input ADA5;
input ADA6;
input ADA7;
input ADA8;
input ADA9;
input ADA10;
input DIB0;
input DIB1;
input DIB2;
input DIB3;
input DIB4;
input DIB5;
input DIB6;
input DIB7;
input DIB8;
input DIB9;
input DIB10;
input DIB11;
input DIB12;
input DIB13;
input DIB14;
input DIB15;
input ADB0;
input ADB1;
input ADB2;
input ADB3;
input ADB4;
input ADB5;
input ADB6;
input ADB7;
input ADB8;
output DOA0;
output DOA1;
output DOA2;
output DOA3;
output DOB0;
output DOB1;
output DOB2;
output DOB3;
output DOB4;
output DOB5;
output DOB6;
output DOB7;
output DOB8;
output DOB9;
output DOB10;
output DOB11;
output DOB12;
output DOB13;
output DOB14;
output DOB15;
endmodule 
module RAMB8K_X8_X8(CENA, CLKA, WRA, CSA0, CSA1, RSTA, CENB, CLKB, WRB, CSB0, CSB1, RSTB, DIA0, DIA1, DIA2, DIA3, DIA4, DIA5, DIA6, DIA7, ADA0, ADA1, ADA2, ADA3, ADA4, ADA5, ADA6, ADA7, ADA8, ADA9, DIB0, DIB1, DIB2, DIB3, DIB4, DIB5, DIB6, DIB7, ADB0, ADB1, ADB2, ADB3, ADB4, ADB5, ADB6, ADB7, ADB8, ADB9, DOA0, DOA1, DOA2, DOA3, DOA4, DOA5, DOA6, DOA7, DOB0, DOB1, DOB2, DOB3, DOB4, DOB5, DOB6, DOB7);// synthesis syn_black_box
input CENA;
input CLKA;
input WRA;
input CSA0;
input CSA1;
input RSTA;
input CENB;
input CLKB;
input WRB;
input CSB0;
input CSB1;
input RSTB;
input DIA0;
input DIA1;
input DIA2;
input DIA3;
input DIA4;
input DIA5;
input DIA6;
input DIA7;
input ADA0;
input ADA1;
input ADA2;
input ADA3;
input ADA4;
input ADA5;
input ADA6;
input ADA7;
input ADA8;
input ADA9;
input DIB0;
input DIB1;
input DIB2;
input DIB3;
input DIB4;
input DIB5;
input DIB6;
input DIB7;
input ADB0;
input ADB1;
input ADB2;
input ADB3;
input ADB4;
input ADB5;
input ADB6;
input ADB7;
input ADB8;
input ADB9;
output DOA0;
output DOA1;
output DOA2;
output DOA3;
output DOA4;
output DOA5;
output DOA6;
output DOA7;
output DOB0;
output DOB1;
output DOB2;
output DOB3;
output DOB4;
output DOB5;
output DOB6;
output DOB7;
endmodule 
module RAMB8K_X8_X16(CENA, CLKA, WRA, CSA0, CSA1, RSTA, CENB, CLKB, WRB, CSB0, CSB1, RSTB, DIA0, DIA1, DIA2, DIA3, DIA4, DIA5, DIA6, DIA7, ADA0, ADA1, ADA2, ADA3, ADA4, ADA5, ADA6, ADA7, ADA8, ADA9, DIB0, DIB1, DIB2, DIB3, DIB4, DIB5, DIB6, DIB7, DIB8, DIB9, DIB10, DIB11, DIB12, DIB13, DIB14, DIB15, ADB0, ADB1, ADB2, ADB3, ADB4, ADB5, ADB6, ADB7, ADB8, DOA0, DOA1, DOA2, DOA3, DOA4, DOA5, DOA6, DOA7, DOB0, DOB1, DOB2, DOB3, DOB4, DOB5, DOB6, DOB7, DOB8, DOB9, DOB10, DOB11, DOB12, DOB13, DOB14, DOB15);// synthesis syn_black_box
input CENA;
input CLKA;
input WRA;
input CSA0;
input CSA1;
input RSTA;
input CENB;
input CLKB;
input WRB;
input CSB0;
input CSB1;
input RSTB;
input DIA0;
input DIA1;
input DIA2;
input DIA3;
input DIA4;
input DIA5;
input DIA6;
input DIA7;
input ADA0;
input ADA1;
input ADA2;
input ADA3;
input ADA4;
input ADA5;
input ADA6;
input ADA7;
input ADA8;
input ADA9;
input DIB0;
input DIB1;
input DIB2;
input DIB3;
input DIB4;
input DIB5;
input DIB6;
input DIB7;
input DIB8;
input DIB9;
input DIB10;
input DIB11;
input DIB12;
input DIB13;
input DIB14;
input DIB15;
input ADB0;
input ADB1;
input ADB2;
input ADB3;
input ADB4;
input ADB5;
input ADB6;
input ADB7;
input ADB8;
output DOA0;
output DOA1;
output DOA2;
output DOA3;
output DOA4;
output DOA5;
output DOA6;
output DOA7;
output DOB0;
output DOB1;
output DOB2;
output DOB3;
output DOB4;
output DOB5;
output DOB6;
output DOB7;
output DOB8;
output DOB9;
output DOB10;
output DOB11;
output DOB12;
output DOB13;
output DOB14;
output DOB15;
endmodule 
module RAMB8K_X16_X16(CENA, CLKA, WRA, CSA0, CSA1, RSTA, CENB, CLKB, WRB, CSB0, CSB1, RSTB, DIA0, DIA1, DIA2, DIA3, DIA4, DIA5, DIA6, DIA7, DIA8, DIA9, DIA10, DIA11, DIA12, DIA13, DIA14, DIA15, ADA0, ADA1, ADA2, ADA3, ADA4, ADA5, ADA6, ADA7, ADA8, DIB0, DIB1, DIB2, DIB3, DIB4, DIB5, DIB6, DIB7, DIB8, DIB9, DIB10, DIB11, DIB12, DIB13, DIB14, DIB15, ADB0, ADB1, ADB2, ADB3, ADB4, ADB5, ADB6, ADB7, ADB8, DOA0, DOA1, DOA2, DOA3, DOA4, DOA5, DOA6, DOA7, DOA8, DOA9, DOA10, DOA11, DOA12, DOA13, DOA14, DOA15, DOB0, DOB1, DOB2, DOB3, DOB4, DOB5, DOB6, DOB7, DOB8, DOB9, DOB10, DOB11, DOB12, DOB13, DOB14, DOB15);// synthesis syn_black_box
input CENA;
input CLKA;
input WRA;
input CSA0;
input CSA1;
input RSTA;
input CENB;
input CLKB;
input WRB;
input CSB0;
input CSB1;
input RSTB;
input DIA0;
input DIA1;
input DIA2;
input DIA3;
input DIA4;
input DIA5;
input DIA6;
input DIA7;
input DIA8;
input DIA9;
input DIA10;
input DIA11;
input DIA12;
input DIA13;
input DIA14;
input DIA15;
input ADA0;
input ADA1;
input ADA2;
input ADA3;
input ADA4;
input ADA5;
input ADA6;
input ADA7;
input ADA8;
input DIB0;
input DIB1;
input DIB2;
input DIB3;
input DIB4;
input DIB5;
input DIB6;
input DIB7;
input DIB8;
input DIB9;
input DIB10;
input DIB11;
input DIB12;
input DIB13;
input DIB14;
input DIB15;
input ADB0;
input ADB1;
input ADB2;
input ADB3;
input ADB4;
input ADB5;
input ADB6;
input ADB7;
input ADB8;
output DOA0;
output DOA1;
output DOA2;
output DOA3;
output DOA4;
output DOA5;
output DOA6;
output DOA7;
output DOA8;
output DOA9;
output DOA10;
output DOA11;
output DOA12;
output DOA13;
output DOA14;
output DOA15;
output DOB0;
output DOB1;
output DOB2;
output DOB3;
output DOB4;
output DOB5;
output DOB6;
output DOB7;
output DOB8;
output DOB9;
output DOB10;
output DOB11;
output DOB12;
output DOB13;
output DOB14;
output DOB15;
endmodule 
module RAMBFIFO512X32A(WE, WCLK, RST, FULLIN, RE, RCLK, EMPTYIN, RPRST, DI0, DI1, DI2, DI3, DI4, DI5, DI6, DI7, DI8, DI9, DI10, DI11, DI12, DI13, DI14, DI15, DI16, DI17, DI18, DI19, DI20, DI21, DI22, DI23, DI24, DI25, DI26, DI27, DI28, DI29, DI30, DI31, DO0, DO1, DO2, DO3, DO4, DO5, DO6, DO7, DO8, DO9, DO10, DO11, DO12, DO13, DO14, DO15, DO16, DO17, DO18, DO19, DO20, DO21, DO22, DO23, DO24, DO25, DO26, DO27, DO28, DO29, DO30, DO31, FULL, AMFULL, EMPTY, AMEMPTY);// synthesis syn_black_box
input WE;
input WCLK;
input RST;
input FULLIN;
input RE;
input RCLK;
input EMPTYIN;
input RPRST;
input DI0;
input DI1;
input DI2;
input DI3;
input DI4;
input DI5;
input DI6;
input DI7;
input DI8;
input DI9;
input DI10;
input DI11;
input DI12;
input DI13;
input DI14;
input DI15;
input DI16;
input DI17;
input DI18;
input DI19;
input DI20;
input DI21;
input DI22;
input DI23;
input DI24;
input DI25;
input DI26;
input DI27;
input DI28;
input DI29;
input DI30;
input DI31;
output DO0;
output DO1;
output DO2;
output DO3;
output DO4;
output DO5;
output DO6;
output DO7;
output DO8;
output DO9;
output DO10;
output DO11;
output DO12;
output DO13;
output DO14;
output DO15;
output DO16;
output DO17;
output DO18;
output DO19;
output DO20;
output DO21;
output DO22;
output DO23;
output DO24;
output DO25;
output DO26;
output DO27;
output DO28;
output DO29;
output DO30;
output DO31;
output FULL;
output AMFULL;
output EMPTY;
output AMEMPTY;
endmodule 
module RAMBFIFO1KX16A(WE, WCLK, RST, FULLIN, RE, RCLK, EMPTYIN, RPRST, DI0, DI1, DI2, DI3, DI4, DI5, DI6, DI7, DI8, DI9, DI10, DI11, DI12, DI13, DI14, DI15, DO0, DO1, DO2, DO3, DO4, DO5, DO6, DO7, DO8, DO9, DO10, DO11, DO12, DO13, DO14, DO15, FULL, AMFULL, EMPTY, AMEMPTY);// synthesis syn_black_box
input WE;
input WCLK;
input RST;
input FULLIN;
input RE;
input RCLK;
input EMPTYIN;
input RPRST;
input DI0;
input DI1;
input DI2;
input DI3;
input DI4;
input DI5;
input DI6;
input DI7;
input DI8;
input DI9;
input DI10;
input DI11;
input DI12;
input DI13;
input DI14;
input DI15;
output DO0;
output DO1;
output DO2;
output DO3;
output DO4;
output DO5;
output DO6;
output DO7;
output DO8;
output DO9;
output DO10;
output DO11;
output DO12;
output DO13;
output DO14;
output DO15;
output FULL;
output AMFULL;
output EMPTY;
output AMEMPTY;
endmodule 
module RAMBFIFO2KX8A(WE, WCLK, RST, FULLIN, RE, RCLK, EMPTYIN, RPRST, DI0, DI1, DI2, DI3, DI4, DI5, DI6, DI7, DO0, DO1, DO2, DO3, DO4, DO5, DO6, DO7, FULL, AMFULL, EMPTY, AMEMPTY);// synthesis syn_black_box
input WE;
input WCLK;
input RST;
input FULLIN;
input RE;
input RCLK;
input EMPTYIN;
input RPRST;
input DI0;
input DI1;
input DI2;
input DI3;
input DI4;
input DI5;
input DI6;
input DI7;
output DO0;
output DO1;
output DO2;
output DO3;
output DO4;
output DO5;
output DO6;
output DO7;
output FULL;
output AMFULL;
output EMPTY;
output AMEMPTY;
endmodule 
module RAMBFIFO4KX4A(WE, WCLK, RST, FULLIN, RE, RCLK, EMPTYIN, RPRST, DI0, DI1, DI2, DI3, DO0, DO1, DO2, DO3, FULL, AMFULL, EMPTY, AMEMPTY);// synthesis syn_black_box
input WE;
input WCLK;
input RST;
input FULLIN;
input RE;
input RCLK;
input EMPTYIN;
input RPRST;
input DI0;
input DI1;
input DI2;
input DI3;
output DO0;
output DO1;
output DO2;
output DO3;
output FULL;
output AMFULL;
output EMPTY;
output AMEMPTY;
endmodule 
module RAMBFIFO8KX2A(WE, WCLK, RST, FULLIN, RE, RCLK, EMPTYIN, RPRST, DI0, DI1, DO0, DO1, FULL, AMFULL, EMPTY, AMEMPTY);// synthesis syn_black_box
input WE;
input WCLK;
input RST;
input FULLIN;
input RE;
input RCLK;
input EMPTYIN;
input RPRST;
input DI0;
input DI1;
output DO0;
output DO1;
output FULL;
output AMFULL;
output EMPTY;
output AMEMPTY;
endmodule 
module RAMBFIFO16KX1A(WE, WCLK, RST, FULLIN, RE, RCLK, EMPTYIN, RPRST, DI0, DO0, FULL, AMFULL, EMPTY, AMEMPTY);// synthesis syn_black_box
input WE;
input WCLK;
input RST;
input FULLIN;
input RE;
input RCLK;
input EMPTYIN;
input RPRST;
input DI0;
output DO0;
output FULL;
output AMFULL;
output EMPTY;
output AMEMPTY;
endmodule 
module CAM128X48(CE, WE, CLK, EN_MASK, WR_MASK, WR_DC, RST, CS0, CS1, WAD0, WAD1, WAD2, WAD3, WAD4, WAD5, WAD6, WD0, WD1, WD2, WD3, WD4, WD5, WD6, WD7, WD8, WD9, WD10, WD11, WD12, WD13, WD14, WD15, WD16, WD17, WD18, WD19, WD20, WD21, WD22, WD23, WD24, WD25, WD26, WD27, WD28, WD29, WD30, WD31, WD32, WD33, WD34, WD35, WD36, WD37, WD38, WD39, WD40, WD41, WD42, WD43, WD44, WD45, WD46, WD47, CO0, CO1, CO2, CO3, CO4, CO5, CO6, MATCH, MUL_MATCH);// synthesis syn_black_box
input CE;
input WE;
input CLK;
input EN_MASK;
input WR_MASK;
input WR_DC;
input RST;
input CS0;
input CS1;
input WAD0;
input WAD1;
input WAD2;
input WAD3;
input WAD4;
input WAD5;
input WAD6;
input WD0;
input WD1;
input WD2;
input WD3;
input WD4;
input WD5;
input WD6;
input WD7;
input WD8;
input WD9;
input WD10;
input WD11;
input WD12;
input WD13;
input WD14;
input WD15;
input WD16;
input WD17;
input WD18;
input WD19;
input WD20;
input WD21;
input WD22;
input WD23;
input WD24;
input WD25;
input WD26;
input WD27;
input WD28;
input WD29;
input WD30;
input WD31;
input WD32;
input WD33;
input WD34;
input WD35;
input WD36;
input WD37;
input WD38;
input WD39;
input WD40;
input WD41;
input WD42;
input WD43;
input WD44;
input WD45;
input WD46;
input WD47;
output CO0;
output CO1;
output CO2;
output CO3;
output CO4;
output CO5;
output CO6;
output MATCH;
output MUL_MATCH;
endmodule 
module CAM128X48CL(CE, WE, CLK, EN_MASK, WR_MASK, WR_DC, RST, CS0, CS1, WAD0, WAD1, WAD2, WAD3, WAD4, WAD5, WAD6, WD0, WD1, WD2, WD3, WD4, WD5, WD6, WD7, WD8, WD9, WD10, WD11, WD12, WD13, WD14, WD15, WD16, WD17, WD18, WD19, WD20, WD21, WD22, WD23, WD24, WD25, WD26, WD27, WD28, WD29, WD30, WD31, WD32, WD33, WD34, WD35, WD36, WD37, WD38, WD39, WD40, WD41, WD42, WD43, WD44, WD45, WD46, WD47, CMO);// synthesis syn_black_box
input CE;
input WE;
input CLK;
input EN_MASK;
input WR_MASK;
input WR_DC;
input RST;
input CS0;
input CS1;
input WAD0;
input WAD1;
input WAD2;
input WAD3;
input WAD4;
input WAD5;
input WAD6;
input WD0;
input WD1;
input WD2;
input WD3;
input WD4;
input WD5;
input WD6;
input WD7;
input WD8;
input WD9;
input WD10;
input WD11;
input WD12;
input WD13;
input WD14;
input WD15;
input WD16;
input WD17;
input WD18;
input WD19;
input WD20;
input WD21;
input WD22;
input WD23;
input WD24;
input WD25;
input WD26;
input WD27;
input WD28;
input WD29;
input WD30;
input WD31;
input WD32;
input WD33;
input WD34;
input WD35;
input WD36;
input WD37;
input WD38;
input WD39;
input WD40;
input WD41;
input WD42;
input WD43;
input WD44;
input WD45;
input WD46;
input WD47;
output [127:0] CMO;
endmodule 
module CAM128X48CM(CE, WE, CLK, EN_MASK, WR_MASK, WR_DC, RST, CS0, CS1, WAD0, WAD1, WAD2, WAD3, WAD4, WAD5, WAD6, WD0, WD1, WD2, WD3, WD4, WD5, WD6, WD7, WD8, WD9, WD10, WD11, WD12, WD13, WD14, WD15, WD16, WD17, WD18, WD19, WD20, WD21, WD22, WD23, WD24, WD25, WD26, WD27, WD28, WD29, WD30, WD31, WD32, WD33, WD34, WD35, WD36, WD37, WD38, WD39, WD40, WD41, WD42, WD43, WD44, WD45, WD46, WD47, CMI, CMO);// synthesis syn_black_box
input CE;
input WE;
input CLK;
input EN_MASK;
input WR_MASK;
input WR_DC;
input RST;
input CS0;
input CS1;
input WAD0;
input WAD1;
input WAD2;
input WAD3;
input WAD4;
input WAD5;
input WAD6;
input WD0;
input WD1;
input WD2;
input WD3;
input WD4;
input WD5;
input WD6;
input WD7;
input WD8;
input WD9;
input WD10;
input WD11;
input WD12;
input WD13;
input WD14;
input WD15;
input WD16;
input WD17;
input WD18;
input WD19;
input WD20;
input WD21;
input WD22;
input WD23;
input WD24;
input WD25;
input WD26;
input WD27;
input WD28;
input WD29;
input WD30;
input WD31;
input WD32;
input WD33;
input WD34;
input WD35;
input WD36;
input WD37;
input WD38;
input WD39;
input WD40;
input WD41;
input WD42;
input WD43;
input WD44;
input WD45;
input WD46;
input WD47;
input [127:0] CMI;
output [127:0] CMO;
endmodule 
module CAM128X48CR(CE, WE, CLK, EN_MASK, WR_MASK, WR_DC, RST, CS0, CS1, WAD0, WAD1, WAD2, WAD3, WAD4, WAD5, WAD6, WD0, WD1, WD2, WD3, WD4, WD5, WD6, WD7, WD8, WD9, WD10, WD11, WD12, WD13, WD14, WD15, WD16, WD17, WD18, WD19, WD20, WD21, WD22, WD23, WD24, WD25, WD26, WD27, WD28, WD29, WD30, WD31, WD32, WD33, WD34, WD35, WD36, WD37, WD38, WD39, WD40, WD41, WD42, WD43, WD44, WD45, WD46, WD47, CMI, CO0, CO1, CO2, CO3, CO4, CO5, CO6, MATCH, MUL_MATCH);// synthesis syn_black_box
input CE;
input WE;
input CLK;
input EN_MASK;
input WR_MASK;
input WR_DC;
input RST;
input CS0;
input CS1;
input WAD0;
input WAD1;
input WAD2;
input WAD3;
input WAD4;
input WAD5;
input WAD6;
input WD0;
input WD1;
input WD2;
input WD3;
input WD4;
input WD5;
input WD6;
input WD7;
input WD8;
input WD9;
input WD10;
input WD11;
input WD12;
input WD13;
input WD14;
input WD15;
input WD16;
input WD17;
input WD18;
input WD19;
input WD20;
input WD21;
input WD22;
input WD23;
input WD24;
input WD25;
input WD26;
input WD27;
input WD28;
input WD29;
input WD30;
input WD31;
input WD32;
input WD33;
input WD34;
input WD35;
input WD36;
input WD37;
input WD38;
input WD39;
input WD40;
input WD41;
input WD42;
input WD43;
input WD44;
input WD45;
input WD46;
input WD47;
input [127:0] CMI;
output CO0;
output CO1;
output CO2;
output CO3;
output CO4;
output CO5;
output CO6;
output MATCH;
output MUL_MATCH;
endmodule 
