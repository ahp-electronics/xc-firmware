--
@ER--RbBF$osHE50RO42RgRgg1b$MDHHO0R$,Q3MO
R--RDqDRosHER0#sCC#s8PC3-
-
R--#CCDOF0HMCR#0CR8VHHM0MHF3WRRCHRIDCDRP0CMkDND$8RN8DRLF_O	sRFl0
FF-N-RsDOEHR#0=CR#D0CO_lsF

---f-R]8CNCRs:/$/#MHbDO$H0/blND.N0jJ4U./b4lbNbC/s#GHHDMDG/HoL/CsMCHoO/CoM_CsMCH/O.s3FlPyE84
Rf-
-
DsHLNRs$HCCC;k

#HCRC3CC#_08DHFoO4_4nNc3D
D;kR#CHCCC38#0_oDFHNO_sEH03DND;#
kCCRHC#C30D8_FOoH_#kMHCoM8D3NDk;
#ICRF3s	obCMNNO	oNC3D
D;
LDHs$NsRHkM#;Hl
Ck#RHkM#3HlPlOFbCFMM30#N;DD
M
C0$H0Rv)m_#LNC#RH
CSoMHCsO
R5SISSHE80RH:RMo0CC:sR=;Rc
SSSNs88I0H8ERR:HCM0oRCs:(=R;S
SSIDFNs88RH:RMo0CC:sR=;Rj
SSSEEHoNs88RH:RMo0CC:sR=UR(;S
SSL0ND:CRRlsF0DNLCS;
SVS8D:0RRlsFI8Fs
;S2
FSbs50R
SSSq)77RH:RM0R#8F_Do_HOP0COF5sRNs88I0H8ERR-4FR8IFM0R;j2
SSS7amzRF:Rk#0R0D8_FOoH_OPC0RFs58IH0-ERR84RF0IMF2Rj
2SS;N
S0H0sLCk0RQQhaRR:#H0sM
o;S0N0skHL0\CR3MsN	:\RR0HMCsoC;R
RR0RN0LsHkR0C\C3slCFP__MFIMNs\RR:HCM0o;Cs
8CMR0CMHR0$)_mvLCN#;N

sHOE00COkRsC#CCDO)0_mFvRVmR)vN_L#HCR##
Sk$L0bsCRFklF0#RHR8#0_oDFHPO_CFO0sH5I8-0E4FR8IFM0R;j2
S--ObFlFMMC0zRvX
wn-S-Sb0FsR-5
-SSSSRmR:kRF00R#8F_Do;HO
S--SQSSjRR:H#MR0D8_FOoH;-
-SSSSQ:4RRRHM#_08DHFoO-;
-SSSSR1R:MRHR8#0_oDFH-O
-SSS2-;
-MSC8FROlMbFC;M0SS

O#FM00NMRGECR#:R0MsHoR5j04FR6:2R=jR"4c.d6Un(gBqA7" w;S

VOkM0MHFRlsF0DNLCNsC8N50LRDC:FRslL0NDRC;IL,R,CRDMRR:HCM0o2CsR0sCkRsM#H0sM=oR>sR"FNl0LsDCC"N8;S

VOkM0MHFRMVkODPN50LF0DFlH_MCVD,RF8IN8Vs_,HREo8EN8Vs_,HRL0M,RL#H0RH:RMo0CCRs2skC0s#MR0MsHo#RH
OSSF0M#NRM00RFb:MRH0CCos=R:R0LF0DFlH_MCVRR+M0LH#RR-4S;
SsPNHDNLC,RHRR[,PL,RbRF#:MRH0CCosS;
SMOF#M0N0FR0bNOEsRR:HCM0oRCs:M=RL#H0Rc/RR4-R;S
SPHNsNCLDRVLkR#:R0MsHoF50bNOEsFR8IFM0R;j2
CSLo
HMSVSH50LF0DFlH_MCVRR<DNFI8_8sVsRFRb0FRE>RHNoE8_8sV02RE
CMS[SSRR:=jS;
SRSP:j=R;S
SSFLb#=R:R
j;SVSSFHsRRRHML0F0FHlDMVC_RR0F0RFbRFDFbS
SSVSHR<HRRIDFNs88_FVRsRRH>HREo8EN8Vs_RC0EMS
SSHSSVVR8DL05HR02=4R''ER0CSM
SSSSS:PR=RRP+*R.*
[;SSSSS8CMR;HV
SSSS#CDCS
SSHSSVNR0L5DCHL25HR02=4R''ER0CSM
SSSSS:PR=RRP+*R.*
[;SSSSS8CMR;HV
SSSS8CMR;HV
SSSS:[R=RR[+;R4RRRR-M-RkClLsVRFR0LH#FRODODC0RC8
SSSS5HV[RR=c02RERCM-C-RP$CsRIcRCkR8lHbRMR0FNERONOsN0
CsSSSSS:[R=;Rj
SSSSkSLVb5LFR#2:E=RCPG52S;
SSSSL#bFRR:=L#bFR4+R;S
SSPSSRR:=jS;
SCSSMH8RVS;
SMSC8FRDF
b;SsSSCs0kMkRLVS;
S#CDCS
SS0sCkRsMs0FlNCLDs8CN5L0NDRC,L0F0FHlDMVC_,HRL0M,RL#H02S;
S8CMR;HV
MSC8kRVMHO0FVMRkPMON
D;
FSOMN#0ML0RFF00lMpHCRR:HCM0oRCs:5=RDNFI8/8s4*n24
n;SMOF#M0N0FRL0l0FdH.pM:CRR0HMCsoCRR:=5IDFNs88/2d.*;d.
FSOMN#0ME0RHpoEHRMC:MRH0CCos=R:RH5Eo8EN84s/n42*nS;
O#FM00NMRoEHEpd.HRMC:MRH0CCos=R:RH5Eo8EN8ds/.d2*.S;
O#FM00NMRoEHEsAF8RCs:MRH0CCos=R:RoEHEMpHCRR+4;6R
FSOMN#0M00Rs0H#N_0CHRR:HCM0oRCs:5=REEHoA8FsC4s+-0LF0pFlH2MC/R4n;0
S$RbC0RNLHN#Rs$sNRE55HdoE.MpHCRR-L0F0F.ldpCHM2./d+84RF0IMF2RjRRFVsFFlk;0R
HS#oDMNRz1map,RmRza:NR0LS;
#MHoN7DRm_zaN,kGRz7mak_NG:.RR8#0_oDFHPO_CFO0sH5I8-0E4FR8IFM0R;j2
oLCHRM
RRRRV_FsbCHb:FRVsRRHHjMRRR0FI0H8ER-4oCCMsCN0
NSS0H0sLCk0Rs\3N\M	RRFVs#CoRD:RNDLCRRH#4R;
RRRRRNRR0H0sLCk0Rs\3CPlFCF_M_sINMF\RVCRso:#RRLDNCHDR#;R4
LSRCMoH
RSSs#Co:HRbbkCLVS
SSFRbsl0RN
b5SRRRSSSSRRRQ=7>Rm_zaN5kGH
2,SRRRSSSSRRRm=7>Rm5zaHS2
SSSSR
2;SMRC8CRoMNCs0VCRFbs_H;bC
H
SVn_4#H:RVER5HdoE.MpHCRR>L0F0F.ldpCHM2CRoMNCs0SC
SoLCHSM
S_HV4:nLRRHV50LF0pFlHRMC=FRL0l0FdH.pMRC2oCCMsCN0
SSSLV:RFLsRHH0RMRRj0IFRHE80R4-RRMoCC0sNCS
SS0SN0LsHkR0CQahQRRFV) mv6RR:DCNLD#RHRMVkODPN50LF0pFlH,MCRIDFNs88,HREo8EN8Rs,L,H0R2d.;S
SSoLCHSM
S)SSm6v R):Rm.vdXS4
SSSSSsbF0NRlbRR5RRqj=q>R757)j
2,SSSSSSSSSRq4=q>R757)4
2,SSSSSSSSSRq.=q>R757).
2,SSSSSSSSSRqd=q>R757)d
2,SSSSSSSSSRqc=q>R757)c
2,SSSSSSSSSRmR=1>Rm5zajL25H
02SSSSSSSSS
2;SCSSMo8RCsMCNR0CLS;
S8CMRMoCC0sNCVRH_L4n;S
SH4V_nRL:H5VRL0F0FHlpM>CRR0LF0dFl.MpHCo2RCsMCN
0CSLSS:FRVsHRL0MRHR0jRFHRI8R0E-RR4oCCMsCN0
SSSS0N0skHL0QCRhRQaF)VRmcv RD:RNDLCRRH#VOkMP5NDL0F0FHlpMRC,DNFI8,8sRoEHE8N8sL,RHR0,4;n2
SSSLHCoMS
SSmS)vR c:mR)vX4n4S
SSSSSb0FsRblNRR5Rq=jR>7Rq7j)52S,
SSSSSSSSq=4R>7Rq74)52S,
SSSSSSSSq=.R>7Rq7.)52S,
SSSSSSSSq=dR>7Rq7d)52S,
SSSSSSSSm=RR>mR1zja52H5L0S2
SSSSSSSS2S;
SMSC8CRoMNCs0LCR;S
SCRM8oCCMsCN0R_HV4;nL
MSC8CRoMNCs0HCRVn_4#
;
S_HVd:.#RRHV5oEHEpd.HRMC=FRL0l0FdH.pMRC2oCCMsCN0
HSSVn_4OH:RVLR5FF00lMpHCRR=L0F0F.ldpCHM2CRoMNCs0SC
S:SLRsVFR0LHRRHMjFR0R8IH0-ERRo4RCsMCN
0CSSSSH4V_:VRHR85N8HsI8R0E=2R4RMoCC0sNCS
SSNSS0H0sLCk0RQQhaVRFRv)m :4RRLDNCHDR#kRVMNOPDF5L0l0FpCHM,FRDI8N8sE,RHNoE8,8sR0LH,nR42S;
SLSSCMoH
SSSSmS)vR 4:mR)vX4n4S
SSSSSSsbF0NRlbRR5RRqj=q>R757)j
2,SSSSSSSSS4SqRR=>',j'
SSSSSSSSqSS.>R=R''j,S
SSSSSSSSSq=dR>jR''S,
SSSSSSSSSRmR=1>Rm5zajL25H
02SSSSSSSSS
2;SSSSCRM8oCCMsCN0R_HV4S;
SHSSV:_.RRHV58N8s8IH0=ERRR.2oCCMsCN0
SSSS0SN0LsHkR0CQahQRRFV) mv.RR:DCNLD#RHRMVkODPN50LF0pFlH,MCRIDFNs88,HREo8EN8Rs,L,H0R24n;S
SSCSLo
HMSSSSSv)m :.RRv)m44nX
SSSSSSSb0FsRblNRR5Rq=jR>7Rq7j)52S,
SSSSSSSSSRq4=q>R757)4
2,SSSSSSSSS.SqRR=>',j'
SSSSSSSSqSSd>R=R''j,S
SSSSSSSSSm=RR>mR1zja52H5L0S2
SSSSSSSS2S;
SCSSMo8RCsMCNR0CH.V_;S
SSVSH_Rd:H5VRNs88I0H8ERR=do2RCsMCN
0CSSSSS0N0skHL0QCRhRQaF)VRmdv RD:RNDLCRRH#VOkMP5NDL0F0FHlpMRC,DNFI8,8sRoEHE8N8sL,RHR0,4;n2
SSSSoLCHSM
SSSS) mvdRR:)4mvn
X4SSSSSbSSFRs0lRNb5qRRj>R=R7q7)25j,S
SSSSSSSSSq=4R>7Rq74)52S,
SSSSSSSSSRq.=q>R757).
2,SSSSSSSSSdSqRR=>',j'
SSSSSSSSmSSR>R=Rz1ma25j50LH2S
SSSSSS
2;SSSSCRM8oCCMsCN0R_HVdS;
SHSSV:_cRRHV5H5Eo8EN8Ls-FF00lMpHCRR<4Rn2NRM858N8s8IH0>ER=2Rc2CRoMNCs0SC
SSSSNs00H0LkChRQQFaRVmR)vR c:NRDLRCDHV#RkPMONLD5FF00lMpHCD,RF8IN8Rs,EEHoNs88,HRL04,Rn
2;SSSSLHCoMS
SS)SSmcv R):Rmnv4XS4
SSSSSFSbsl0RN5bRRjRqRR=>q)775,j2
SSSSSSSSqSS4>R=R7q7)254,S
SSSSSSSSSq=.R>7Rq7.)52S,
SSSSSSSSSRqd=q>R757)d
2,SSSSSSSSSRSmRR=>1amz55j2L2H0
SSSSSSSS;S2
SSSS8CMRMoCC0sNCVRH_
c;SSSSH6V_:VRHRN558I8sHE80RR>=6N2RM58REEHoNs88RL-RFF00lMpHC=R>R24n2CRoMNCs0SC
SSSSNs00H0LkChRQQFaRVmR)vR 6:NRDLRCDHV#RkPMONLD5FF00lMpHCD,RF8IN8Rs,EEHoNs88,HRL0d,R.
2;SSSSLHCoMS
SS)SSm6v R):Rm.vdXS4
SSSSSFSbsl0RN5bRRjRqRR=>q)775,j2
SSSSSSSSqSS4>R=R7q7)254,S
SSSSSSSSSq=.R>7Rq7.)52S,
SSSSSSSSSRqd=q>R757)d
2,SSSSSSSSScSqRR=>q)775,c2
SSSSSSSSmSSR>R=Rz1ma25j50LH2S
SSSSSS2SS;S
SSMSC8CRoMNCs0HCRV;_6
SSSCRM8oCCMsCN0R
L;SMSC8CRoMNCs0HCRVn_4OS;
S_HV4:n8RRHV50LF0pFlHRMC>FRL0l0FdH.pMRC2oCCMsCN0
SSSHNV_8HsI8:0ERRHV58N8s8IH0>ERRRc2oCCMsCN0
SSSSRL:VRFsLRH0HjMRRR0FI0H8ERR-4CRoMNCs0SC
SSSSHcV_:VRHRE55HNoE8-8sL0F0FHlDM<CRR24nR8NMR85N8HsI8R0E>c=R2o2RCsMCN
0CSSSSS0SN0LsHkR0CQahQRRFV) mvcRR:DCNLD#RHRMVkODPN50LF0pFlH,MCRIDFNs88,HREo8EN8Rs,L,H0R24n;S
SSLSSCMoH
SSSS)SSmcv R):Rmnv4XS4
SSSSSbSSFRs0lRNb5jRqRR=>q)775,j2
SSSSSSSSSSSq=4R>7Rq74)52S,
SSSSSSSSS.SqRR=>q)775,.2
SSSSSSSSSSSq=dR>7Rq7d)52S,
SSSSSSSSSRSm=1>Rm5zajL25H
02SSSSSSSSS2SS;S
SSCSSMo8RCsMCNR0CHcV_;S
SSMSC8CRoMNCs0LCR;S
SS8CMRMoCC0sNCVRH_sN8I0H8ES;
SVSH_8N8s8IH0RE:H5VRNs88I0H8E=R<RRc2oCCMsCN0
SSSSRL:VRFsLRH0HjMRRR0FI0H8ERR-4CRoMNCs0SC
SSSSH4V_:VRHR85N8HsI8R0E=2R4RMoCC0sNCS
SSSSSNs00H0LkChRQQFaRVmR)vR 4:NRDLRCDHV#RkPMONLD5FF00lMpHCD,RF8IN8Rs,EEHoNs88,HRL04,Rn
2;SSSSSoLCHSM
SSSSSv)m :4RRv)m44nX
SSSSSSSSsbF0NRlbRR5RRqj=q>R757)j
2,SSSSSSSSSqSS4>R=R''j,S
SSSSSSSSSSRq.='>Rj
',SSSSSSSSSqSSd>R=R''j,S
SSSSSSSSSSRmR=1>Rm5zajL25H
02SSSSSSSSS;S2
SSSSMSC8CRoMNCs0HCRV;_4
SSSSVSH_R.:H5VRNs88I0H8ERR=.o2RCsMCN
0CSSSSS0SN0LsHkR0CQahQRRFV) mv.RR:DCNLD#RHRMVkODPN50LF0pFlH,MCRIDFNs88,HREo8EN8Rs,L,H0R24n;S
SSLSSCMoH
SSSS)SSm.v R):Rmnv4XS4
SSSSSbSSFRs0lRNb5qRRj>R=R7q7)25j,S
SSSSSSSSSSRq4=q>R757)4
2,SSSSSSSSSqSS.>R=R''j,S
SSSSSSSSSSRqd='>Rj
',SSSSSSSSSmSSR>R=Rz1ma25j50LH2S
SSSSSSSSS2S;
SSSSCRM8oCCMsCN0R_HV.S;
SSSSHdV_:VRHR85N8HsI8R0E=2RdRMoCC0sNCS
SSSSSNs00H0LkChRQQFaRVmR)vR d:NRDLRCDHV#RkPMONLD5FF00lMpHCD,RF8IN8Rs,EEHoNs88,HRL04,Rn
2;SSSSSoLCHSM
SSSSSv)m :dRRv)m44nX
SSSSSSSSsbF0NRlbRR5RRqj=q>R757)j
2,SSSSSSSSSqSS4>R=R7q7)254,S
SSSSSSSSSSRq.=q>R757).
2,SSSSSSSSSqSSd>R=R''j,S
SSSSSSSSSSRmR=1>Rm5zajL25H
02SSSSSSSS2S;
SSSSCRM8oCCMsCN0R_HVdS;
SSSSHcV_:VRHRE55HNoE8-8sL0F0FHlDM<CRR24nR8NMR85N8HsI8R0E>c=R2o2RCsMCN
0CSSSSS0SN0LsHkR0CQahQRRFV) mvcRR:DCNLD#RHRMVkODPN50LF0pFlH,MCRIDFNs88,HREo8EN8Rs,L,H0R24n;S
SSLSSCMoH
SSSS)SSmcv R):Rmnv4XS4
SSSSSbSSFRs0lRNb5qRRj>R=R7q7)25j,S
SSSSSSSSSSRq4=q>R757)4
2,SSSSSSSSSqSS.>R=R7q7)25.,S
SSSSSSSSSSRqd=q>R757)d
2,SSSSSSSSSmSSR>R=Rz1ma25j50LH2S
SSSSSS;S2
SSSSMSC8CRoMNCs0HCRV;_c
SSSS8CMRMoCC0sNC;RL
SSSCRM8oCCMsCN0R_HVNs88I0H8ES;
S8CMRMoCC0sNCVRH_84n;C
SMo8RCsMCNR0CHdV_.
#;
4SL:FRVsRRIH4MRRR0F5oEHEpd.HRMC-FRL0l0FdH.pMdC-.d2/.CRoMNCs0SC
SRL:VRFsLRH0HjMRRR0FI0H8ERR-4CRoMNCs0SC
S0SN0LsHkR0CQahQRRFV) mv6RR:DCNLD#RHRMVkODPN5dI*.F+L0l0FdH.pMRC,DNFI8,8sRoEHE8N8sL,RHR0,d;.2
SSS#MHoNbDRH_bC80Fk#RR:#_08DHFoOS;
SoLCHSM
SmS)vR 6:mR)vXd.4S
SSbSSFRs0lRNb5qRRj>R=R7q7)25j,S
SSSSSS4SqRR=>q)775,42
SSSSSSSSRq.=q>R757).
2,SSSSSSSSq=dR>7Rq7d)52S,
SSSSSqSSc>R=R7q7)25c,S
SSSSSSRSmRR=>1amz55I2L2H0
SSSSSSS2S;
S8CMRMoCC0sNC;RL
MSC8CRoMNCs0LCR4
;
S_HV4:nFRRHV5H5Eo.EdpCHMRR=REEHopCHM2MRN8ER5HdoE.MpHCRR>L0F0F.ldpCHM2o2RCsMCN
0CS:SLRsVFR0LHRRHMjFR0R8IH0-ERRo4RCsMCN
0CS#SSHNoMDkRF0M_C8RR:#_08DHFoOS;
S0SN0LsHkR0CQahQRRFV) mvcRR:DCNLD#RHRMVkODPN5oEHEsAF8-Cs4R6,EEHoA8FsC4s-6E,RHNoE8,8sR0LH,nR42S;
SoLCHSM
SmS)vR c:mR)vX4n4S
SSbSSFRs0lRNb5jRqR>R=R7q7)25j,S
SSSSSS4SqRR=>q)775,42
SSSSSSSSRq.=q>R757).
2,SSSSSSSSq=dR>7Rq7d)52S,
SSSSSmSSR>R=Rz1maE55HdoE.MpHCF-L0l0FdH.pMdC-.d2/.2+450LH2S
SSSSSS
2;SMSC8CRoMNCs0LCR;C
SMo8RCsMCNR0CH4V_n
F;S_HV4:n#RRHV5H5Eo.EdpCHMRR<REEHopCHM2MRN8ER5HdoE.MpHCRR>L0F0F.ldpCHM2o2RCsMCN
0CS:SLRsVFR0LHRRHMjFR0R8IH0-ERRo4RCsMCN
0CS#SSHNoMDkRF0M_C8RR:#_08DHFoOS;
S0SN0LsHkR0CQahQRRFV) mv6RR:DCNLD#RHRMVkODPN5oEHEsAF8-CsdR4,EEHoA8FsCds-4E,RHNoE8,8sR0LH,.Rd2S;
SoLCHSM
SmS)vR 6:mR)vXd.4S
SSbSSFRs0lRNb5qRRj>R=R7q7)25j,S
SSSSSS4SqRR=>q)775,42
SSSSSSSSRq.=q>R757).
2,SSSSSSSSq=dR>7Rq7d)52S,
SSSSSqSSc>R=R7q7)25c,S
SSSSSSRSmRR=>1amz5H5Eo.EdpCHM-0LF0dFl.MpHCd2/.L25H
02SSSSS2SS;S
SCRM8oCCMsCN0R
L;S8CMRMoCC0sNCVRH_#4n;R

RHRRVH_I8:0ERRHV5H0s#00NCR_H<2R6RMoCC0sNCR
RRRRRRVRH_0FkjH:RVER5HdoE.MpHCRR=L0F0F.ldpCHM2CRoMNCs0RC
RRRRRRRRRmRpzja52=R<Rz1ma25j;R
RRRRRRMRC8CRoMNCs0HCRVk_F0
j;RRRRRRRRHFV_k:04RRHV5oEHEpd.HRMC>FRL0l0FdH.pMRC2oCCMsCN0
RRRRRRRRRRRHOV_N4#C:VRHRF5L0l0FpCHMRL=RFF00lpd.H2MCRMoCC0sNC-
-SHS#oDMNRV8HVRR:#_08DHFoOS;
RLRRCMoH
R--RRRRRRRRRRRRRV8HV=R<R''jRCIEM7Rq7<)R=mRBh1e_ap7_mBtQ_Be a5m)dL4+FF00lMpHCN,R8I8sHE802-R
-RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRDRC#'CR4
';-R-SRRRRRsVF_8IH0RE:VRFsHMRHR0jRFHRI8-0E4CRoMNCs0-C
-RSRRRRRRlRRksG0C:CRRXvzw-n
-SSSb0FsRblNR-5
-SSSSmRRR>R=Rzpma25j5,H2
S--SRSSRRQj=1>Rm5zajH252-,
-SSSSQRR4>R=Rz1ma2545,H2
S--SRSSRR1R=8>RH
VV-S-SS
2;-R-RRRRRRRRRRRRRCRM8oCCMsCN0RsVF_8IH0
E;RRRRRRRRRRRRRmRpzja52=R<Rz1ma25jRCIEM7Rq7<)R=mRBh1e_ap7_mBtQ_Be a5m)dL4+FF00lMpHCN,R8I8sHE802RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRCCD#Rz1ma254;R
RRRRRRRRRR8CMRMoCC0sNCVRH_#ONC
4;RRRRRRRRRHRRVN_O#:C.RRHV50LF0pFlHRMC>FRL0l0FdH.pMRC2oCCMsCN0
S--So#HMRND8VHVjRR:#_08DHFoOS;
RRRRLHCoM-
-RRRRRRRRRRRRRHR8VRVj<'=RjI'RERCMq)77RR<=Bemh_71a_tpmQeB_ mBa)654+0LF0pFlH,MCR8N8s8IH0RE2
R--RRRRRRRRRRRRRRRRRRRRRRRRRRRRRCRRDR#C';4'
S--RRRRRFRVsH_I8j0E:FRVsRRHHjMRRR0FI0H8ER-4oCCMsCN0
S--RRRRRRRRRGlk0CsCRv:RznXw
S--SFSbsl0RN5bR
S--SRSSRRmR=p>Rm5zajH252-,
-SSSSQRRj>R=Rz1ma25j5,H2
S--SRSSRRQ4=1>Rm5za4H252-,
-SSSS1RRR>R=RV8HV-j
-SSS2-;
-RRRRRRRRRRRRCRRMo8RCsMCNR0CV_FsI0H8E
j;RRRRRRRRRRRRRmRpzja52=R<Rz1ma25jRCIEM7Rq7<)R=mRBh1e_ap7_mBtQ_Be a5m)4L6+FF00lMpHCN,R8I8sHE802RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRCCD#Rz1ma254;R
RRRRRRRRRR8CMRMoCC0sNCVRH_#ONC
.;RRRRRRRRCRM8oCCMsCN0R_HVF4k0;R
RRRRRR:RNRsVFRHIRMRR405FREEHodH.pM-CRR0LF0dFl.MpHC.-d2./d-o4RCsMCN
0C-S-S#MHoN8DRH4VVR#:R0D8_FOoH_OPC05Fs5oEHEpd.HRMC-FRL0l0FdH.pMdC-.d2/.R-48MFI04FR2S;
RRRRLHCoM-
-RRRRRRRRRRRRRHR8V5V4I<2R=jR''ERICqMR7R7)<mRBh1e_ap7_mBtQ_Be a5m)d5.*I2+4+0LF0dFl.MpHCN,R8I8sHE802-
-RRRRRRRRRRRRRRRRRRRRRRRRRRRRR#CDC4R''-;
-RSRRRRRV_FsI0H8ER4:VRFsHMRHR0jRFHRI8-0E4CRoMNCs0-C
-RSRRRRRRlRRksG0C:CRRXvzw-n
-SSSb0FsRblNR-5
-SSSSmRRR>R=Rzpma25I5,H2
S--SRSSRRQj=p>Rm5zaI2-45,H2
S--SRSSRRQ4=1>Rm5zaI2+45,H2
S--SRSSRR1R=8>RH4VV5
I2-S-SS
2;-R-RRRRRRRRRRRRRCRM8oCCMsCN0RsVF_8IH0;E4
RRRRRRRRRRRRpRRm5zaI<2R=mRpzIa5-R42IMECR7q7)RR<Bemh_71a_tpmQeB_ mBa).5d*+5I4L2+FF00lpd.H,MCR8N8s8IH0
E2RRRRRRRRRRRRRRRRRRRRRRRRRRRRR#CDCmR1zIa5+;42
RRRRRRRR8CMRMoCC0sNC;RN
RRRR
RRRRRRRRRRHDV_N4#0nH:RV5R5EEHodH.pM=CRRoEHEMpHCN2RM58REEHodH.pM-CRR0LF0dFl.MpHCRR>n2d2RMoCC0sNC-
-SHS#oDMNRV8HV:.RR8#0_oDFH
O;SRRRRoLCH-M
-RRRRRRRRRRRR8RRH.VVRR<='Rj'IMECR7q7)RR<Bemh_71a_tpmQeB_ mBa)H5EoFEAss8C-,46R8N8s8IH0RE2
R--RRRRRRRRRRRRRRRRRRRRRRRRRRRRCCD#R''4;-
-SRRRRVRRFIs_HE80.V:RFHsRRRHMjFR0R8IH04E-RMoCC0sNC-
-SRRRRRRRRkRlGC0sCRR:vwzXn-
-SbSSFRs0lRNb5-
-SSSSRRRmRR=>pamz5H5Eo.EdpCHM-0LF0dFl.MpHC.-d2./d225H,-
-SSSSRjRQRR=>pamz5H5Eo.EdpCHM-0LF0dFl.MpHC.-d2./d-542H
2,-S-SSRSRQ=4R>mR1z5a5EEHodH.pMLC-FF00lpd.H2MC/2d.5,H2
S--SRSSRR1R=8>RH.VV
S--S;S2
R--RRRRRRRRRRRRR8CMRMoCC0sNCFRVsH_I8.0E;R
RRRRRRRRRRmRpz5a5EEHodH.pMLC-FF00lpd.H-MCd/.2dR.2<p=Rm5za5oEHEpd.H-MCL0F0F.ldpCHM-2d./-d.4
2RSSSSSCIEM7Rq7<)RRhBmea_17m_pt_QBea BmE)5HAoEFCs8s6-4,8RN8HsI820E
RRRRRRRRRRRRRRRRRRRR#CDCmR1z5a5EEHodH.pMLC-FF00lpd.H2MC/2d.;R
RRRRRRMRC8CRoMNCs0HCRVN_D#n04;R

RRRRRHRRVN_D#.0d:VRHRE55HdoE.MpHCRR<RoEHEMpHCN2RM58REEHodH.pM-CRR0LF0dFl.MpHCRR>n2d2RMoCC0sNC-
-SHS#oDMNRV8HV:dRR8#0_oDFH
O;SRRRRoLCH-M
-RRRRRRRRRRRR8RRHdVVRR<='Rj'IMECR7q7)RR<Bemh_71a_tpmQeB_ mBa)H5EoFEAss8C-,d4R8N8s8IH0RE2
R--RRRRRRRRRRRRRRRRRRRRRRRRRRRRCCD#R''4;-
-SRRRRVRRFIs_HE80dV:RFHsRRRHMjFR0R8IH04E-RMoCC0sNC-
-SRRRRRRRRkRlGC0sCRR:vwzXn-
-SbSSFRs0lRNb5-
-SSSSRRRmRR=>pamz5H5Eo.EdpCHM-0LF0dFl.MpHC.-d2./d225H,-
-SSSSRjRQRR=>pamz5H5Eo.EdpCHM-0LF0dFl.MpHC.-d2./d-542H
2,-S-SSRSRQ=4R>mR1z5a5EEHodH.pMLC-FF00lpd.H2MC/2d.5,H2
S--SRSSRR1R=8>RHdVV
S--S;S2
R--RRRRRRRRRRRRR8CMRMoCC0sNCFRVsH_I8d0E;R
RRRRRRRRRRmRpz5a5EEHodH.pMLC-FF00lpd.H-MCd/.2dR.2<p=Rm5za5oEHEpd.H-MCL0F0F.ldpCHM-2d./-d.4
2RSSSSSCIEM7Rq7<)RRhBmea_17m_pt_QBea BmE)5HAoEFCs8s4-d,8RN8HsI820E
RRRRRRRRRRRRRRRRRRRR#CDCmR1z5a5EEHodH.pMLC-FF00lpd.H2MC/2d.;R
RRRRRRMRC8CRoMNCs0HCRVN_D#.0d;R

RRRRRHRRVk_F0R.:H5VREEHoA8FsC-sRR0LF0pFlHRMC<cRn2CRoMNCs0RC
RRRRRRRRRRRRRz7mak_NG=R<RD8V0ERIC5MRRRRR57q7)RR>Bemh_71a_tpmQeB_ mBa)H5EoFEAss8C,8RN8HsI820E2R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRFRRsqR57R7)<mRBh1e_ap7_mBtQ_Be a5m)L0F0FHlpMRC,Ns88I0H8E222
RRRRRRRRRRRRRRRRRRRRRRRRRRRCCD#Rzpma25j;R
RRRRRRMRC8CRoMNCs0HCRVk_F0
.;RRRRRRRRHFV_k:0dRRHV5oEHEsAF8RCs-FRL0l0FpCHMRn>Rdo2RCsMCN
0CRRRRRRRRRRRRRmR7zNa_k<GR=VR8DI0RERCM5RRRR75q7>)RRhBmea_17m_pt_QBea BmE)5HAoEFCs8sN,R8I8sHE802R2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRFs57q7)RR<Bemh_71a_tpmQeB_ mBa)F5L0l0FpCHM,8RN8HsI820E2R2
RRRRRRRRRRRRRRRRRRRRRRRRRDRC#pCRm5za5oEHEpd.H-MCL0F0F.ldpCHM-2d./2d.;R
RRRRRRMRC8CRoMNCs0HCRVk_F0
d;RRRRR8CMRMoCC0sNCVRH_8IH0
E;R
RRRRRRR_HVI0H8ERj:H5VR0#sH0CN0_>HR=2R6RMoCC0sNCR
RRRRRRVRH_#ONCR4:H5VRL0F0FHlpM=CRR0LF0dFl.MpHCo2RCsMCN
0CRRRRRRRRR7RRm_zaNRkG<1=Rm5zajI2RERCM5RRRR75q7<)R=mRBh1e_ap7_mBtQ_Be a5m)dL4+FF00lMpHCN,R8I8sHE802
2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR8NMR75q7>)R=mRBh1e_ap7_mBtQ_Be a5m)L0F0FHlpMRC,Ns88I0H8E222
RRRRRRRRRRRRRRRRRRRRRRRRRRRCCD#RlsFF'k05EF0CRs#='>RZ;'2
RRRRRRRR8CMRMoCC0sNCVRH_#ONC
4;RRRRRRRRHOV_N.#C:VRHRF5L0l0FpCHMRL>RFF00lpd.H2MCRMoCC0sNCR
RRRRRRRRRRz7mak_NG=R<Rz1ma25jRCIEMRR5R5RRq)77RR<=Bemh_71a_tpmQeB_ mBa)654+0LF0pFlH,MCR8N8s8IH02E2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRSRRR8NMR75q7>)R=mRBh1e_ap7_mBtQ_Be a5m)L0F0FHlpMRC,Ns88I0H8E222
RRRRRRRRRRRRRRRRRRRRRRRRRRRCCD#RlsFF'k05EF0CRs#='>RZ;'2
RRRRRRRR8CMRMoCC0sNCVRH_#ONC
.;RRRRRRRRNRj:VRFsIMRHR04RFER5HdoE.MpHCF-L0l0FdH.pMdC-.d2/.CRoMNCs0RC
RRRRRRRRRRRRRz7mak_NG=R<Rz1ma25IRCIEMRR5R5RRq)77RR<=Bemh_71a_tpmQeB_ mBa).5d*+5I4R2+L0F0F.ldpCHM-R4,Ns88I0H8E
22RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRNRM857q7)=R>RhBmea_17m_pt_QBea Bmd)5.+*IL0F0F.ldpCHM,8RN8HsI820E2R2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR#CDCFRsl0Fk'05FE#CsRR=>'2Z';R
RRRRRRMRC8CRoMNCs0NCRjR;
RRRRRHRRVk_#b:d.RRHV5H5Eo.EdpCHMRR=REEHopCHM2MRN8ER5HdoE.MpHCRR-L0F0F.ldpCHMRn>RdR22oCCMsCN0
RRRRRRRRRRRR7RRm_zaNRkG<1=Rm5za5oEHEpd.H-MCL0F0F.ldpCHM2./d2SR
SRSRSSSSIMECRR5RRqR57R7)<B=Rm_he1_a7pQmtB _eB)am5oEHEsAF8,CsR8N8s8IH02E2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRNRRM58Rq)77RR>=Bemh_71a_tpmQeB_ mBa)H5EoFEAss8C-,46R8N8s8IH02E22R
RRRRRRRRRRRRRRRRRRRRRRRRRRDRC#sCRFklF0F'50sEC#>R=R''Z2R;
RRRRRCRRMo8RCsMCNR0CH#V_k.bd;R
RRRRRRVRH_b#k4Rn:H5VR5oEHEpd.HRMC<ERRHpoEH2MCR8NMRH5Eo.EdpCHMRL-RFF00lpd.HRMC>dRn2o2RCsMCN
0CRRRRRRRRRRRRRmR7zNa_k<GR=mR1z5a5EEHodH.pMLC-FF00lpd.H2MC/2d.RS
SSSRRSISSERCM5RRRR75q7<)R=mRBh1e_ap7_mBtQ_Be a5m)EEHoA8FsCRs,Ns88I0H8E
22RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRMRN8qR57R7)>B=Rm_he1_a7pQmtB _eB)am5oEHEsAF8-CsdR4,Ns88I0H8E222
RRRRRRRRRRRRRRRRRRRRRRRRRRRR#CDCFRsl0Fk'05FE#CsRR=>'2Z';R
RRRRRRMRC8CRoMNCs0HCRVk_#b;4n
RRRRRRRR_HVD:FIRRHV50LF0pFlHRMC>2RjRMoCC0sNCR
RRRRRRRRRRz7mak_NG=R<RD8V0ERIC5MRR5RRq)77RB<Rm_he1_a7pQmtB _eB)am50LF0pFlH,MCR8N8s8IH02E2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRSRRRsRFR75q7>)RRhBmea_17m_pt_QBea BmE)5HAoEFCs8sN,R8I8sHE802
22RRRRRRRRRRRRRRRRRRRRRRRRCCD#RlsFF'k05EF0CRs#='>RZ;'2
RRRRRRRR8CMRMoCC0sNCVRH_IDF;R
RRRRRRVRH_IDFjH:RVLR5FF00lMpHCRR<4o2RCsMCN
0CRRRRRRRRR7RRm_zaNRkG<8=RVRD0IMECR75q7>)RRhBmea_17m_pt_QBea BmE)5HAoEFCs8sN,R8I8sHE802R2
RRRRRRRRRRRRRRRRRRRRRCRRDR#CsFFlk50'FC0Es=#R>ZR''
2;RRRRRRRRCRM8oCCMsCN0R_HVDjFI;R
RRCRRMo8RCsMCNR0CHIV_HE80j
;
CRM8NEsOHO0C0CksRD#CC_O0);mv
H
DLssN$CRHC
C;kR#CHCCC38#0_oDFH4O_43ncN;DD
Ck#RCHCC03#8F_Do_HON0sHED3NDk;
#HCRC3CC#_08DHFoOM_k#MHoCN83D
D;kR#CI	Fs3MoCb	NON3oCN;DD
H
DLssN$MRkHl#H;#
kCMRkHl#H3FPOlMbFC#M03DND;C

M00H$mR)v#RH
CSoMHCsO
R5SVSSNDlH$RR:#H0sM:oR=NR"M;$"
SSSI0H8ERR:HCM0oRCs:c=R;S
SS8N8s8IH0:ERR0HMCsoCRR:=(S;
SFSDI8N8sRR:HCM0oRCs:j=R;S
SSoEHE8N8sRR:HCM0oRCs:(=RUS;
SNS0LRDC:FRslL0ND
C;S8SSVRD0:FRslsIF82
S;b
SFRs05S
SS7q7)RR:H#MR0D8_FOoH_OPC0RFs58N8s8IH0-ERR84RF0IMF2Rj;S
SSz7maRR:FRk0#_08DHFoOC_POs0FRH5I8R0E-RR48MFI0jFR2S
S2
;
S0N0skHL0\CR3MsN	:\RR0HMCsoC;R
RR0RN0LsHkR0C\C3slCFP__MFIMNs\RR:HCM0o;Cs
8CMR0CMHR0$);mv
s
NO0EHCkO0s#CRCODC0m_)vVRFRv)mR
H#SlOFbCFMM)0RmLv_N
#CSCSoMHCsO
R5SSSSI0H8ERR:HCM0o;Cs
SSSS8N8s8IH0:ERR0HMCsoC;S
SSFSDI8N8sRR:HCM0o;Cs
SSSSoEHE8N8sRR:HCM0o;Cs
SSSSL0ND:CRRlsF0DNLCS;
S8SSVRD0:FRslsIF8S
S2S;
SsbF0
R5SSSSq)77RH:RM0R#8F_Do_HOP0COF5sRNs88I0H8ERR-4FR8IFM0R;j2
SSSSz7maRR:FRk0#_08DHFoOC_POs0FRH5I8R0E-RR48MFI0jFR2S
SS
2;S8CMRlOFbCFMM
0;
FSOMN#0MM0R0:LRR0HMCsoCRR:=4
n;
kSVMHO0F#MR00Ns)pFlHRMCskC0sHMRMo0CCHsR#S
SPHNsNCLDRx#HCRR:HCM0o;Cs
OSSF0M#NRM0LODF	x#HCRR:HCM0oRCs:M=R0*LRR;nc
CSLo
HMSVSHRF5DI8N8sFRl8DRLF#O	H2xCRR=RjER0CSM
SCSs0MksRIDFNs88RL+RD	FO#CHx;S
SCCD#
SSSskC0s5MR5IDFNs88RL+RD	FO#CHxR4-R2RR/LODF	x#HC*2RRFLDOH	#x
C;SMSC8VRH;C
SMV8Rk0MOHRFM#s0N0l)FpCHM;S

O#FM00NMRFLDOH	#x:CRR0HMCsoCRR:=n*cRRLM0;O
SF0M#NRM0DqHl8R8s:MRH0CCos=R:RN#0sF0)lMpHC
;RSMOF#M0N0LRM_lsF_NVsORR:HCM0oRCs:5=REEHoNs88RD-RH8lq8+sRR/42RFLDOH	#x
C;SMOF#M0N0CRDVs0_FVl_sRNO:MRH0CCos=R:RH5Eo8EN8-sRRlDHqs88R4+R2FRl8DRLF#O	H;xC
0
S$RbC0DNLCF_8kH0R#sRNsRN$5_MLs_FlVOsN+84RF0IMF2RjRRFVsIFlF;s8
#
SHNoMDFR8ks0_F:lRRL0ND8C_F;k0
oLCH
M
S_HVL)HomRv:H5VREEHoNs88RD-RF8IN8+sRR>4RRFLDOH	#xRC2oCCMsCN0
#SSHNoMDFR8kV0_H0s#,mR7zNa_k:GRRlsFI8Fs;S
S#MHoNqDR7_7)N,kGR7q7)R_V:0R#8F_Do_HOP0COF5sRNs88I0H8ERR-4FR8IFM0R;j2
CSLo
HM
VSSFbs_H:bCRsVFRHHRMRRj0NFR8I8sHE80-o4RCsMCN
0CSNSS0H0sLCk0Rs\3N\M	RRFVs#CoqRR:DCNLD#RHR
j;SNSS0H0sLCk0Rs\3N\M	RRFVs#CoARR:DCNLD#RHR
4;RRRRRRRRRRRRNs00H0LkC3R\sFClPMC_FN_IsRM\FsVRCqo#RD:RNDLCRRH#4R;
RRRRRRRRRNRR0H0sLCk0Rs\3CPlFCF_M_sINMF\RVCRsoR#A:NRDLRCDH4#R;S
SLHCoMS
SSosC#Rq:bCHbL
kVSbSSFRs0l5Nb
SSSSQSRRR=>q)775,H2
SSSSRRSm>R=R7q7)5_VHS2
SSSS2
;
SsSSCAo#:HRbbkCLVS
SSsbF0NRlbS5
SSSSR=QR>7Rq7V)_5,H2
SSSSRRSm>R=R7q7)k_NG25H
SSSS;S2
CSSMo8RCsMCNR0CV_FsbCHb;S

Sv)m R4(:mR)vN_L#SC
SCSoMHCsONRlbS5
SISSHE80R=SS>HRI8,0E
SSSS8N8s8IH0RERSR=>Ns88I0H8E
,RSSSSDNFI8R8sR=RS>FRDI8N8sS,
SESSHNoE8R8sR=RS>HRDl8q8s,-4
SSSSL0NDRCRR>S=RL0ND
C,SSSS80VDRSRRSR=>80VD
SSS2S
SSsbF0NRlbRR5R7q7)>R=R7q7),_VRS
SSSSS7amzRR=>80Fk_sVH#S0
SSSS2
;S
8SSF_k0s5Flj<2R=FR8kV0_H0s#RCIEMqR57_7)NRkG>B=Rm_he1_a7pQmtB _eB)am5IDFNs88,8RN8HsI820E2S
SSSSSSRSRR#CDCVR8D
0;
VSSFDs_F:FbRsVFRHHRMRR40MFRLF_sls_VNoORCsMCN
0CS#SSHNoMDFR8k#0_0CNoRs:RFFlIs
8;SCSLo
HMS)SSm6v R):RmLv_N
#CSoSSCsMCHlORN
b5SSSSI0H8ESRS=I>RHE80,S
SS8SN8HsI8R0ER>S=R8N8s8IH0RE,
SSSSIDFNs88RSRR=D>RH8lq8+sRR-5H4L2*D	FO#CHx,S
SSHSEo8EN8RsRR>S=RlDHqs88RH+R*FLDOH	#x4C-,SR
S0SSNCLDRSRR=0>RNCLD,S
SSVS8DR0RR=SS>VR8DS0
S
S2SbSSFRs0lRNb5qRR7R7)=q>R7_7)V
,RSSSSSmS7z=aR>FR8k#0_0CNo
SSSS;S2SS

SFS8ks0_FHl52=R<Rk8F00_#NRoCIMECR75q7N)_k>GR=mRBh1e_ap7_mBtQ_Be a5m)DqHl8+8s54H-2D*LF#O	H,xCR8N8s8IH02E2
SSSSSSSSRRRCCD#Rk8F0F_sl-5H4
2;SMSC8CRoMNCs0VCRFDs_F;Fb
SS
S_HV#CHx:VRHRC5DVs0_FVl_sRNO>2RjRMoCC0sNCS
SSo#HMRND80Fk_N#0o:CRRlsFI8Fs;S
SLHCoMS
SSv)m :6RRv)m_#LNCS
SSMoCCOsHRblN5S
SSHSI8R0ES>S=R8IH0
E,SSSSNs88I0H8ESRR=N>R8I8sHE80,SR
SDSSF8IN8RsRR>S=RlDHqs88RM+RLF_sls_VNLO*D	FO#CHx,S
SSHSEo8EN8RsRR>S=RoEHE8N8s
,RSSSS0DNLCRRRSR=>0DNLCS,
S8SSVRD0RSRS=8>RV
D0S2SS
SSSb0FsRblNRR5Rq)77RR=>q)77_RV,
SSSS7SSmRza=8>RF_k0#o0NCS
SS2SS;SS

SSS80Fk_lsF5_MLs_FlVOsN+R42<8=RF_k0s5FlMsL_FVl_s2NO
SSSSSSSSSSSIMECR75q7N)_k<GRRhBmea_17m_pt_QBea BmD)5H8lq8Ms+LF_sls_VNLO*D	FO#CHx,8RN8HsI820E2S
SSSSSSRSRRRSSRCRRDR#C80Fk_N#0o
C;SS
SSz7mak_NG=R<RD8V0ERIC5MRq)77_GNkRB>Rm_he1_a7pQmtB _eB)am5oEHE8N8sN,R8I8sHE802S2
SSSSSCSRDR#C80Fk_lsF5_MLs_FlVOsN+;42
CSSMo8RCsMCNR0CH#V_H;xC
SS
S_HVMx#HCH:RVDR5C_V0s_FlVOsNRj=R2CRoMNCs0SC
SmS7zNa_k<GR=VR8DI0RERCM57q7)k_NGRR>Bemh_71a_tpmQeB_ mBa)H5Eo8EN8Rs,Ns88I0H8E
22SSSSSRSSCCD#Rk8F0F_slL5M_lsF_NVsO
2;SMSC8CRoMNCs0HCRV#_MH;xC
S
SV_FsbCHb:FRVsRRHHjMRRR0FI0H8ER-4oCCMsCN0
SSSNs00H0LkC3R\s	NM\VRFRosC#RR:DCNLD#RHR
.;RRRRRRRRRRRRNs00H0LkC3R\sFClPMC_FN_IsRM\FsVRCRo#:NRDLRCDH4#R;S
SRoLCHSM
SsSRC:o#RbbHCVLk
SSSSFRbsl0RN
b5SRSRRSSSSQRRRR=>7amz_GNk5,H2
RSSRSRSSRSRm>R=Rz7ma25H
SSSSRSS2S;
SMRC8CRoMNCs0VCRFbs_H;bC
C
SMo8RCsMCNR0CHLV_Hmo)v
;
S_HV#DlNDv)m:VRHRH5Eo8EN8-sRRIDFNs88R4+RRR<=LODF	x#HCo2RCsMCN
0CSHS#oDMNR7q7)R_V:0R#8F_Do_HOP0COF5sRNs88I0H8ERR-4FR8IFM0R;j2
CSLo
HMSFSVsH_bbRC:VRFsHMRHR0jRF8RN8HsI8-0E4CRoMNCs0SC
S0N0skHL0\CR3MsN	F\RVCRsoR#q:NRDLRCDHj#R;S
SNs00H0LkC3R\sFClPMC_FN_IsRM\FsVRCqo#RD:RNDLCRRH#4S;
SoLCHSM
SCSso:#qRbbHCVLk
SSSSsbF0NRlbS5
SSSSQ>R=R7q7)25H,S
SSmSSRR=>q)77_HV52S
SS;S2
CSSMo8RCsMCNR0CV_FsbCHb;S

) mv6RR:)_mvLCN#
SSSSMoCCOsHRblN5S
SSSSSS8IH0SERSR=>I0H8ER,
RSSSSSSSNs88I0H8ERRR=N>R8I8sHE80,SR
SSSSSFSDI8N8sRRRSR=>DNFI8,8s
SSSSSSSEEHoNs88RSRR=E>RHNoE8,8s
SSSSSSS0DNLCRRRSR=>0DNLCS,
SSSSSVS8DR0RR=SS>VR8DS0
SSSSS
S2SSSSb0FsRblNRR5Rq)77RR=>q)77_RV,
SSSSSSS7amzRR=>7amz
SSSS2SS;
S
S8CMRMoCC0sNCVRH_N#lDmD)v
;
CRM8NEsOHO0C0CksRD#CC_O0);mv
