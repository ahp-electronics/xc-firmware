----------------------------------------------------------------------------
--
-- Dummy package for backward compatibility of the designs
-- All the procedures defined herein are already part of
-- the Vhdl 2008 IEEE std_logic_1164 package, so available 
-- to designers. This file is only to stub out the use 
-- clauses made in the old designs.
-- 
----------------------------------------------------------------------------

package std_logic_textio is
end std_logic_textio;

package body std_logic_textio is

end std_logic_textio;
