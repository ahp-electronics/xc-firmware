--
@ER--B$FbsEHo0OR52gR4g-cRRj.jd$R1MHbDO$H0ROQM
R--fN]C8:CsR#//$DMbH0OH$N/lb0DN.Uj4J4.b/blNb#Cs/DGHH/MGD/HLoCCMs/HOo_CMoCCMs.HO/lsNMI_s38PEyf4R

--

-----
-HR1lCbDRv)qR0IHEHR#MCoDR7q7)1 1RsVFR0LFECRsNN8RMI8RsCH0
R--aoNsC:0RRDXHH
MG
LDHs$NsRCHCC
;
kR#CHCCC38#0_oDFH4O_43ncN;DD
Ck#RCHCC03#8F_Do_HO#MHoCN83D
D;DsHLNRs$k#MHH
l;kR#Ck#MHHPl3ObFlFMMC0N#3D
D;CHM00)$Rq_vh)HWR#R
RRCRoMHCsO
R5RRRRRRRRVHNlD:$RRs#0HRMo:"=RMCFM"R;
RRRRRIRRHE80RH:RMo0CC:sR=jR4;RR
RRRRRNRR8I8sHE80RH:RMo0CC:sR=dR4;RRRRRRRRR--LRHoCkMFoVERF8sRCEb0
RRRRRRRRb8C0:ERR0HMCsoCRR:=U.4g;R
RRRRRRFR8ks0_C:oRRFLFDMCNRR:=V#NDCR;RR-RR-NRE#kRF00bkRosC
RRRRRRRRM8H_osCRL:RFCFDN:MR=NRVD;#CRRRRR-R-R#ENR08NNMRHbRk0s
CoSRRRR0s#_08NNRR:#H0sM
o;SsSI_8lFCRR:#H0sM:oR=WR") Qa_)wQ1;a"
RRRRRRRR8N8sC_soRR:LDFFCRNM:0=RsRkCRRRRRR--ERN8Ns88CR##s
CoRRRRRRRR2R;
RbRRFRs05R
RRRRRRmR7zRa:FRk0#_08DHFoOC_POs0F58IH04E-RI8FMR0Fj
2;RRRRRRRR7RQhRH:RM0R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj;R
RRRRRR7Rq7:)RRRHM#_08DHFoOC_POs0F58N8s8IH04E-RI8FMR0Fj
2;RRRRRRRRWR R:MRHR8#0_oDFHRO;RRRRR-R-RHIs0CCRMDNLCFRVsNRslR
RRRRRRpRBiRR:H#MR0D8_FOoH;RRRRRRR-O-RD	FORsVFRlsN,8RN8Rs,8
HMSBSmp:iRRRHM#_08DHFoOS;
Sa)1RH:RM0R#8F_Do;HORRRRR-RR-CRs#RC0FFMRkk0b0CRsoS
S :hRRRHM#_08DHFoORSSRR--CbMRHFMRVDRLFRO	s
NlS;S2
8CMR0CMHR0$)hqv_;)W
s
NO0EHCkO0sLCRD	FO_lsNRRFV)hqv_R)WHV#
k0MOHRFMVOkM_HHM0R5L:FRLFNDCMs2RCs0kM0R#soHMR
H#LHCoMR
RH5VRL02RE
CMRRRRskC0s"M5"
2;RDRC#RC
RsRRCs0kMB5"F8kDR0MFRbHlDCClMA0RD	FORv)q3#RQRC0ERNsC88RN8#sC#CRso0H#C8sCRHk#M0oRE#CRNRlCOODF	#RNRC0ERv)q?;"2
CRRMH8RVC;
MV8Rk_MOH0MH;0
N0LsHkR0CoCCMsFN0sC_sb0FsR#:R0MsHo-;
-0N0skHL0oCRCsMCNs0F_bsCFRs0FLVRD	FO_lsNRN:RsHOE00COkRsCHV#Rk_MOH0MH5k8F0C_so
2;VOkM0MHFRs#0H.Mo#5DPNRR:#H0sMRo2skC0s#MR0D8_FOoH_OPC0RFsHP#
NNsHLRDC#RDP:0R#8F_Do_HOP0COFNs5'oEHE'-NDRFI8MFI0jFR2P;
NNsHLRDCHRR:HCM0o;Cs
oLCHRM
RsVFRHHRMRRj0#FRDEP'HRoEDbFF
RRRRRHV5NN5'oEHE2-HR'=R4R'20MEC
RSR#5DPH:2R=4R''S;
CCD#
RSR#5DPH:2R=jR''S;
CRM8H
V;RMRC8FRDF
b;RCRs0MksRP#D;M
C80R#soHM.P#D;k
VMHO0F#MRD#P.0MsHoR5N:0R#8F_Do_HOP0COFRs2skC0s#MR0MsHo#RH
sPNHDNLCRR#:0R#soHM5EN'H-oENF'DIR+48MFI04FR2P;
NNsHLRDCHRR:HCM0o;Cs
oLCHRM
RsVFRHHRM'RNDRFI0NFR'oEHEFRDFRb
RHRRVNR55RH2=4R''02RE
CMS#RR5NH-'IDF+R42:'=R4
';S#CDCR
SRH#5-DN'F4I+2=R:R''j;C
SMH8RVR;
R8CMRFDFbR;
R0sCkRsM#C;
M#8RD#P.0MsHoN;
0H0sLCk0R_GObbsF#RR:#H0sM
o;-F-OMN#0M#0RsDPNR#:R0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2=R:Rs#0H.Mo#5DPs_#08NN02-;
-CRLoRHMLODF	NRsllRHblDCCNM00MHFRo#HM#ND
MVkOF0HMCRo0E_OFCHO_8IH0IE5HE80RH:RMo0CCRs2skC0sHMRMo0CCHsR#N
PsLHNDPCRN:DRR0HMCsoCRR:=jP;
NNsHLRDC8dHP.8,RHnP4,HR8PRU,8cHP,HR8PR.,84HPRH:RMo0CC
s;LHCoMR
R8dHP.=R:RH5I8-0E4d2/nR;
RP8H4:nR=IR5HE80-/424
U;RHR8P:UR=IR5HE80-/42gR;
RP8Hc=R:RH5I8-0E4c2/;R
R8.HPRR:=58IH04E-2;/.
8RRHRP4:5=RI0H8E2-4;R
RH5VR84HPRj>R2ER0CRM
RPRRN:DR=NRPDRR+4R;
R8CMR;HV
HRRV8R5HRP.>2RjRC0EMR
RRNRPD=R:RDPNR4+R;R
RCRM8H
V;RVRHRH58P>cRRRj20MEC
RRRRDPNRR:=PRND+;R4
CRRMH8RVR;
RRHV5P8HURR>j02RE
CMRRRRPRND:P=RN+DRR
4;RMRC8VRH;R
RH5VR84HPnRR>j02RE
CMRRRRPRND:P=RN+DRR
4;RMRC8VRH;-
-RVRHRH58PRd.>2RjRC0EM-
-RRRRPRND:P=RN+DRR
4;-R-RCRM8H
V;RVRHRN5PDRR>.02RE
CMRRRRskC0s5MR.*R*RDPNR.+RRR**5DPNRd-R2
2;RDRC#RC
RsRRCs0kM.R5RR**P2ND;R
RCRM8HRV;RRRRRCR
Mo8RCO0_EOFHCH_I8;0E
MVkOF0HMCRo0E_OFCHO_b8C08E5CEb0RH:RMo0CCRs2skC0sHMRMo0CCHsR#N
PsLHND8CR_FOEH_OC80CbERR:HCM0oRCs:j=R;C
Lo
HMRVRHRC58bR0E>4RUgR.20MEC
RRRRO8_EOFHCC_8bR0E:4=RncdU;R
RCHD#V8R5CEb0RR<=U.4gR8NMRb8C0>ERRgcjnRR20MEC
RRRRO8_EOFHCC_8bR0E:U=R4;g.
CRRDV#HRC58bR0E<c=RjRgnNRM880CbERR>.Ujc2ER0CRM
R8RR_FOEH_OC80CbE=R:RgcjnR;
R#CDH5VR80CbE=R<Rc.jUMRN8CR8bR0E>jR4.2cRRC0EMR
RR_R8OHEFO8C_CEb0RR:=.Ujc;R
RCHD#V8R5CEb0RR<=4cj.R8NMRb8C0>ERR.642ER0CRM
R8RR_FOEH_OC80CbE=R:R.4jcR;
R#CDH5VR80CbE=R<R.642ER0CRM
R8RR_FOEH_OC80CbE=R:R.64;R
RCRM8H
V;RCRs0MksRO8_EOFHCC_8b;0E
8CMR0oC_FOEH_OC80CbEV;
k0MOHRFMo_C0I0H8EF_l85_UOHEFOIC_8RR:HCM0o2CsR0sCkRsMHCM0oRCsHP#
NNsHLRDCI0H8EF_l8R_U:MRH0CCosL;
CMoH
HRRVOR5EOFHC8_IRU>R2ER0CRM
RIRRHE80_8lF_:UR=EROFCHO_RI8-OR5EOFHC8_IR8lFR;U2
CRRD
#CRRRRI0H8EF_l8R_U:O=REOFHC8_I;R
RCRM8H
V;RCRs0MksR8IH0lE_FU8_;M
C8CRo0H_I8_0El_F8U
;
O#FM00NMROI_EOFHCH_I8R0E:MRH0CCos=R:R0oC_FOEH_OCI0H8EH5I820E;F
OMN#0MI0R_FOEH_OC80CbERR:HCM0oRCs:4=RncdU/0oC_8IH0lE_FU8_5OI_EOFHCH_I820E;F
OMN#0M80R_FOEH_OC80CbERR:HCM0oRCs:o=RCO0_EOFHCC_8b50E80CbE
2;O#FM00NMRO8_EOFHCH_I8R0E:MRH0CCos=R:Rn54d/Uc8E_OFCHO_b8C0RE2+5R54Undc_/8OHEFO8C_CEb02RR/U
2;
MVkOF0HMCRo0k_MlC_OD5D#I:8RR0HMCsoC;FOEH_OCI:8RR0HMCsoC2CRs0MksR0HMCsoCR
H#PHNsNCLDRlMk_DOCD:#RR0HMCsoC;C
Lo
HMRkRMlC_ODRD#:5=RI48-2E/OFCHO_RI8+;R4
sRRCs0kMkRMlC_OD;D#
8CMR0oC_lMk_DOCD
#;
MVkOF0HMCRo0H_#xIC5M:ORR0HMCsoC;MR8ORR:HCM0o2CsR0sCkRsMHCM0oRCsHL#
CMoH
RRRskC0sIMRM*ORRO8M;M
C8CRo0H_#x
C;
MVkOF0HMCRo0F_LF5D88H_#x:CRR0HMCsoC;_RI#CHxRH:RMo0CCRs;8I_ORH:RMo0CCRs;II_ORH:RMo0CCRs2skC0sHMRMo0CCHsR#C
Lo
HMH5VR8H_#x<CR=_RI#CHx2ER0CRM
R0sCkRsM8I_O;D
C#RC
R0sCkRsMII_O;M
C8VRH;M
C8CRo0F_LF;D8
MVkOF0HMCRo0M_C8C_8b50E#CHxRH:RMo0CC;sRRb8C0:ERR0HMCsoC2CRs0MksR0HMCsoCR
H#PHNsNCLDRMlH_x#HCRR:HCM0oRCs:j=R;C
Lo
HMRHRlMH_#x:CR=CR8b;0E
HRRV#R5HRxC<CR8b20ERC0EMR
RRHRlMH_#x:CR=HR#x
C;RMRC8VRH;R
RskC0slMRH#M_H;xC
8CMR0oC_8CM_b8C0
E;
MOF#M0N0EROFCHO_8IH0:ERR0HMCsoCRR:=o_C0LDFF8C5o0H_#xoC5CM0_kOl_C#DD58IH0RE,8E_OFCHO_8IH0,E2o_C0M_klODCD#C58b,0ERO8_EOFHCC_8b20E2R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRo_C0#CHx50oC_lMk_DOCDI#5HE80,_RIOHEFOIC_HE802C,o0k_MlC_OD5D#80CbEI,R_FOEH_OC80CbE,22
SSSSSSSSSSSRO8_EOFHCH_I8,0EROI_EOFHCH_I820E;F
OMN#0MI0RHE80_lMk_DOCD:#RR0HMCsoCRR:=o_C0LDFF8C5o0H_#xoC5CM0_kOl_C#DD58IH0RE,8E_OFCHO_8IH0,E2o_C0M_klODCD#C58b,0ERO8_EOFHCC_8b20E2R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRoRRC#0_H5xCo_C0M_klODCD#H5I8,0EROI_EOFHCH_I820E,0oC_lMk_DOCD8#5CEb0,_RIOHEFO8C_CEb02
2,SSSSSSSSSRSSR5RRI0H8E2-4/O8_EOFHCH_I8,0ERH5I8-0E4I2/_FOEH_OCI0H8E+2RR
4;O#FM00NMRb8C0ME_kOl_C#DDRH:RMo0CC:sR=CRo0F_LF5D8o_C0#CHx50oC_lMk_DOCDI#5HE80,_R8OHEFOIC_HE802C,o0k_MlC_OD5D#80CbE8,R_FOEH_OC80CbE,22
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRo_C0#CHx50oC_lMk_DOCDI#5HE80,_RIOHEFOIC_HE802C,o0k_MlC_OD5D#80CbEI,R_FOEH_OC80CbE,22
SSSSSSSSRSSR8R5CEb0-/428E_OFCHO_b8C0RE,5b8C04E-2_/IOHEFO8C_CEb02RR+4R;S
MOF#M0N0CRxs:FRR8#0_oDFHPO_CFO0sE5OFCHO_8IH0IE*HE80_lMk_DOCDI#-HE80-84RF0IMF2RjRR:=5EF0CRs#='>Rj;'2
MOF#M0N0sR#P_ND#RDP:0R#8F_Do_HOP0COFOs5EOFHCH_I8*0EI0H8Ek_MlC_OD-D#4FR8IFM0RRj2:x=RCRsF&0R#soHM.P#D50s#_08NN
2;O#FM00NMRP#sN:DRRs#0H5MoOHEFOIC_HE80*8IH0ME_kOl_C#DDRI8FMR0F4:2R=DR#P0.#soHM5P#sN#D_D;P2
#--HNoMDV#RFMsRFDM-#bENCL8RD	FORlsN#$
0bFCRkL0_k_#40C$bRRH#NNss$8R5CEb0_lMk_DOCD4#-RI8FMR0FjI,RHE80_lMk_DOCD4#-RI8FMR0FjF2RV0R#8F_Do;HO
o#HMRNDF_k0L4k#RF:RkL0_k_#40C$b;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFV80FkRM5HbRk000FRs#H-0CN0#02
$RbCF_k0L.k#_b0$C#RHRsNsN5$R80CbEk_MlC_OD-D#4FR8IFM0RRj,.H*I8_0EM_klODCD#R+48MFI0jFR2VRFR8#0_oDFH
O;#MHoNFDRkL0_kR#.:kRF0k_L#0._$;bCRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$F8VRFRk05bHMk00RFsR0H0-#N#0C2$
0bFCRkL0_k_#c0C$bRRH#NNss$8R5CEb0_lMk_DOCD4#-RI8FMR0Fjc,R*8IH0ME_kOl_C#DD+8dRF0IMF2RjRRFV#_08DHFoO#;
HNoMDkRF0k_L#:cRR0Fk_#Lkc$_0bRC;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RVFR8k50RHkMb0FR0RH0s-N#002C#
b0$CkRF0k_L#0U_$RbCHN#Rs$sNRC58b_0EM_klODCD#R-48MFI0jFR,*RUI0H8Ek_MlC_OD+D#(FR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNR0Fk_#LkURR:F_k0LUk#_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFRk8F0HR5M0bkRR0F0-sH#00NC
#20C$bRsbNH_0$LUk#_b0$C#RHRsNsN5$R80CbEk_MlC_OD-D#4FR8IFM0RRj,I0H8Ek_MlC_OD-D#4FR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNRsbNH_0$LUk#Rb:RN0sH$k_L#0U_$;bCRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFRk8F0HR5M0bkRR0F0-sH#00NC
#20C$bR0Fk_#Lk40n_$RbCHN#Rs$sNRC58b_0EM_klODCD#R-48MFI0jFR,nR4*8IH0ME_kOl_C#DD+R468MFI0jFR2VRFR8#0_oDFH
O;#MHoNFDRkL0_kn#4RF:RkL0_kn#4_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$F8VRFRk05bHMk00RFsR0H0-#N#0C2$
0bbCRN0sH$k_L#_4n0C$bRRH#NNss$8R5CEb0_lMk_DOCD4#-RI8FMR0Fj.,R*8IH0ME_kOl_C#DD+84RF0IMF2RjRRFV#_08DHFoO#;
HNoMDNRbs$H0_#Lk4:nRRsbNH_0$L4k#n$_0bRC;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RVFR8k50RHkMb0FR0RH0s-N#002C#
b0$CkRF0k_L#_d.0C$bRRH#NNss$8R5CEb0_lMk_DOCD4#-RI8FMR0Fjd,R.H*I8_0EM_klODCD#4+dRI8FMR0FjF2RV0R#8F_Do;HO
o#HMRNDF_k0Ldk#.RR:F_k0Ldk#.$_0bRC;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFV80FkRM5HbRk000FRs#H-0CN0#02
$RbCbHNs0L$_k.#d_b0$C#RHRsNsN5$R80CbEk_MlC_OD-D#4FR8IFM0RRj,cH*I8_0EM_klODCD#R+d8MFI0jFR2VRFR8#0_oDFH
O;#MHoNbDRN0sH$k_L#Rd.:NRbs$H0_#Lkd0._$;bCRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$F8VRFRk05bHMk00RFsR0H0-#N#0C2H
#oDMNR0Fk_RCM:0R#8F_Do_HOP0COF8s5CEb0_lMk_DOCD4#-RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-C-RMDNLCV#RF0sRs#H-0CN0#H
#oDMNR0Is_RCM:0R#8F_Do_HOP0COF8s5CEb0_lMk_DOCD4#-RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-I-RsCH0RNCML#DCRsVFROCNEFRsIVRFRv)qRDOCD##
HNoMDMRH_osCR#:R0D8_FOoH_OPC05FsI0H8E6+dRI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RCk#8FR0RosCHC#0sQR7h#R
HNoMDkRF0C_soRR:#_08DHFoOC_POs0F58IH0dE+6FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RCk#8FR0RosCHC#0smR7z#a
HNoMD8RN_osCR#:R0D8_FOoH_OPC05FsNs88I0H8ER-48MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--k8#CRR0FsHCo#s0CR7q7)H
#oDMNRIDF_8N8sRR:#_08DHFoOC_POs0F5R4d8MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--Ns88R0LH#MRHbRk00)FRqOvRC#DDRR5cL#H0RJsCkCHs8#2
HNoMD8RNsRCo:0R#8F_Do_HOP0COFNs58I8sHE80-84RF0IMF2Rj;-R-RR0FsHCo#s0CRC0ERD#CCRO0#MHoNFDRVsR0HN#00-C
-MRC8DRLFRO	sRNlHDlbCMlC0HN0F#MRHNoMDN#
0H0sLCk0Rs\3NFl_VCV#0:\RRs#0H;Mo
C
Lo
HMRRR
R-RR-VRQR8N8s8IH0<ERRFOEH_OCI0H8E#RN#MHoR''jRR0Fk#MkCL8RH
0#RRRRzRjR:VRHR85N8HsI8R0E=2R4RMoCC0sNCR
SRDRRFNI_8R8s<"=Rjjjjjjjjjjjjj&"RR_N8s5Coj
2;S8CMRMoCC0sNCjRz;R
RR4RzRRR:H5VRNs88I0H8ERR=.o2RCsMCN
0CSRRRRIDF_8N8s=R<Rj"jjjjjjjjjjRj"&8RN_osC584RF0IMF2Rj;C
SMo8RCsMCNR0Cz
4;RRRRzR.R:VRHR85N8HsI8R0E=2RdRMoCC0sNCR
SRDRRFNI_8R8s<"=Rjjjjjjjjj"jjRN&R8C_soR5.8MFI0jFR2S;
CRM8oCCMsCN0R;z.
RRRRRzdRH:RVNR58I8sHE80Rc=R2CRoMNCs0SC
RRRRD_FINs88RR<="jjjjjjjj"jjRN&R8C_soR5d8MFI0jFR2S;
CRM8oCCMsCN0R;zd
RRRRRzcRH:RVNR58I8sHE80R6=R2CRoMNCs0SC
RRRRD_FINs88RR<="jjjjjjjjRj"&8RN_osC58cRF0IMF2Rj;C
SMo8RCsMCNR0Cz
c;RRRRzR6R:VRHR85N8HsI8R0E=2RnRMoCC0sNCR
SRDRRFNI_8R8s<"=Rjjjjjjjj"RR&Ns8_C6o5RI8FMR0Fj
2;S8CMRMoCC0sNC6Rz;R
RRnRzRRR:H5VRNs88I0H8ERR=(o2RCsMCN
0CSRRRRIDF_8N8s=R<Rj"jjjjjj&"RR_N8s5ConFR8IFM0R;j2
MSC8CRoMNCs0zCRnR;
RzRR(:RRRRHV58N8s8IH0=ERRRU2oCCMsCN0
RSRRFRDI8_N8<sR=jR"jjjjj&"RR_N8s5Co(FR8IFM0R;j2
MSC8CRoMNCs0zCR(R;
RzRRU:RRRRHV58N8s8IH0=ERRRg2oCCMsCN0
RSRRFRDI8_N8<sR=jR"jjjj"RR&Ns8_CUo5RI8FMR0Fj
2;S8CMRMoCC0sNCURz;R
RRgRzRRR:H5VRNs88I0H8ERR=4Rj2oCCMsCN0
RSRRFRDI8_N8<sR=jR"j"jjRN&R8C_soR5g8MFI0jFR2S;
CRM8oCCMsCN0R;zg
RRRRjz4RRR:H5VRNs88I0H8ERR=4R42oCCMsCN0
RSRRFRDI8_N8<sR=jR"jRj"&8RN_osC5R4j8MFI0jFR2S;
CRM8oCCMsCN0Rjz4;R
RR4Rz4:RRRRHV58N8s8IH0=ERR24.RMoCC0sNCR
SRDRRFNI_8R8s<"=RjRj"&8RN_osC5R448MFI0jFR2S;
CRM8oCCMsCN0R4z4;R
RR4Rz.:RRRRHV58N8s8IH0=ERR24dRMoCC0sNCR
SRDRRFNI_8R8s<'=Rj&'RR_N8s5Co48.RF0IMF2Rj;C
SMo8RCsMCNR0Cz;4.
RRRRdz4RRR:H5VRNs88I0H8ERR>4Rd2oCCMsCN0
RSRRFRDI8_N8<sR=8RN_osC5R4d8MFI0jFR2S;
CRM8oCCMsCN0Rdz4;R

R-RR-VRQRH58MC_sos2RC#oH0RCs7RQhkM#HopRBiR
RR4Rzc:RRRRHV5M8H_osC2CRoMNCs0RC
RRRRRbRRsCFO#5#RB,piRh7Q2CRLo
HMRRRRRRRRRRRRH5VRBRpi=4R''MRN8pRBiP'CC2M0RC0EMR
RRRRRRRRRRRRRRMRH_osCRR<=5j"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjRj"&QR7h
2;RRRRRRRRRRRRCRM8H
V;RRRRRRRRCRM8bOsFC;##
MSC8CRoMNCs0zCR4
c;RRRRzR46RH:RVMR5F80RHsM_CRo2oCCMsCN0
RRRRRRRRRRRR_HMsRCo<5=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj&"RRh7Q2S;
CRM8oCCMsCN0R6z4;R

R7RRmRza<F=Rks0_CIo5HE80-84RF0IMF2Rj;R

RNRR8C_so=R<R7q7)R;
R-RR-CRtMNCs00CRE)CRqOvRC#DDR8NMRD#CCRO0DHFoOFRVsqR)vnA4__141R4
RzRR4:URRRHV5FOEH_OCI0H8ERR=4o2RCsMCN
0CSzRRORE	:VRHRN5R8I8sHE80R4>RcRR2oCCMsCN0
RRRRRRRRDzO	b:RsCFO#5#RB2pi
RSRRRRRLHCoMR
SRRRRRVRHRp5BiP'CCRM0NRM8BRpi=4R''02RE
CMSRRRRRRRRNRR8osC58N8s8IH04E-RI8FMR0F4Rc2<N=R8C_so85N8HsI8-0E4FR8IFM0R24c;S
SRCRRMH8RVS;
S8CMRFbsO#C#RDkO	S;
RMRC8CRoMNCs0zCRO;E	
RRRRRRRRgz4RV:RFHsRRRHM5b8C0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CRRRR-Q-RVNR58I8sHE80R4>RcM2RCRC80OFRs0CNCsRIHR0CCLMNDNCRMF8Rkk0b0MRCNCLDRD#CCRO0DHFoOR
RRRRRRzRS.:jRRRHV58N8s8IH0>ERR24cRMoCC0sNC-
S-HRVGFRVsNROD4DRd(UU,CR#D0CORRFV0#sH0CN0R0MFRHLCMsoRC#oH0CCs8R
RRRRRRRRRRRRRRkRF0M_C5RH2<'=R4I'RERCM5sN8CNo58I8sHE80-84RF0IMFcR42RR=HC2RDR#C';j'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RWRCIEMNR58C_so85N8HsI8-0E4FR8IFM0R24cRH=R2DRC#'CRj
';RRRRRRRRS8CMRMoCC0sNC.RzjR;
R-RR-VRQR85N8HsI8R0E<4=R.M2RFsRIHR0CCLMNDFCRskRF00bkRNCMLRDC#CCDOD0RFOoHRCMC8
C8RRRRRRRRRRRRzR.4:VRHR85N8HsI8R0E<4=Rco2RCsMCN
0CRRRRRRRRRRRRRRRRF_k0CHM52=R<R''4;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R R;
RRRRRRRRRCRRMo8RCsMCNR0Cz;.4
RRRRR--tCCMsCN0RC0ERv)qRDOCDN#RM08Rs#H-0CN0#R
RRRRRRzRS.:.RRsVFRH[RMIR5HE80_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNCS
SS0N0skHL0GCROs_bFRb#FAVR)_qv4UndcRX4:NRDLRCDH"#R1q)epR="&sR#P5ND[2+4R"&R,)RWQ_a v m7=&"RR_IslCF8;R
RRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqA)vn_4dXUc4RR:DCNLD#RHR1"Aa&"RR0HMCsoC'NHloIC5HE802RR&"R7"&MRH0CCosl'HN5oCHn*4d2UcR"&RW&"RR0HMCsoC'NHlo[C52RR&"R "&MRH0CCosl'HN5oCo_C0C_M880CbEH55R4+R2n*4d,UcRb8C02E2R"&RX&"RR0HMCsoC'NHlo[C5+;42
SSSLHCoMR
RRRRRRRRRRARS)_qv4UndcRX4:qR)vnA4_
14SRRRRRRRRRRRRsbF0NRlb7R5Q25jRR=>HsM_C[o52q,R7R7)=D>RFNI_858s48dRF0IMF2Rj,hR RR=> Rh,1R1)=)>R1
a,SSSSW= R>sRI0M_C5,H2RiBpRR=>B,piR57mj=2R>kRF0k_L#H45,2[2;R
RRRRRRRRRRRRRRkRF0C_so25[RR<=F_k0L4k#5[H,2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRSRRCRM8oCCMsCN0R.z.;R
RRRRRRMRC8CRoMNCs0zCR4
g;RRRRCRM8oCCMsCN0RUz4;RRRRR
RRRRR
RRRRR--tCCMsCN0RC0ERv)qRDOCDN#RM#8RCODC0FRDoRHOVRFs)Aqv41n_.z
S.:dRRRHV5FOEH_OCI0H8ERR=.o2RCsMCN
0CS-S-RGVHRsVFRDONDdR4U,U(RD#CCRO0F0VRs0H#NR0CMRF0LMCHoCRso0H#C8sC
RSRz	OERH:RVRR5Ns88I0H8ERR>4Rd2oCCMsCN0
RRRRRRRRDzO	b:RsCFO#5#RB2pi
RSRRRRRLHCoMR
SRRRRRVRHRp5BiP'CCRM0NRM8BRpi=4R''02RE
CMSRRRRRRRRNRR8osC58N8s8IH04E-RI8FMR0F4Rd2<N=R8C_so85N8HsI8-0E4FR8IFM0R24d;S
SRCRRMH8RVS;
S8CMRFbsO#C#RDkO	S;
RMRC8CRoMNCs0zCRO;E	
RRRR.SzcRR:VRFsHMRHRC58b_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
-S-RRQV58N8s8IH0>ERR24dRCMC8FR0RCOsNR0CI0sHCMRCNCLDR8NMR0FkbRk0CLMND#CRCODC0FRDo
HORRRRRRRRS6z.RH:RVNR58I8sHE80R4>Rdo2RCsMCN
0CSR--VRHGVRFsODNDRU4dUR(,#CCDOF0RVsR0HN#00MCRFL0RCoHMRosCHC#0s
C8RRRRRRRRRRRRRRRRF_k0CHM52=R<R''4RCIEMNR58osC58N8s8IH04E-RI8FMR0F4Rd2=2RHR#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=WI RERCM5_N8s5CoNs88I0H8ER-48MFI04FRd=2RRRH2CCD#R''j;R
RRRRRRCRSMo8RCsMCNR0Cz;.6
-S-RRQV58N8s8IH0<ER=dR42FRMRHIs0CCRMDNLCsRFR0FkbRk0CLMND#CRCODC0FRDoRHOM8CCCR8
SRRRR.SznRR:H5VRNs88I0H8E=R<R24dRMoCC0sNCR
SRRRRRRRRRFRRkC0_M25HRR<=';4'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RW;R
RRRRRRCRSMo8RCsMCNR0Cz;.n
-S-RMtCC0sNCER0CqR)vCRODRD#NRM80-sH#00NCR#
RRRRRSRRzR.(:FRVsRR[H5MRI0H8Ek_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0SC
S0SN0LsHkR0CGbO_s#FbRRFVAv)q_gU4.RX.:NRDLRCDH"#R1q)epR="&sR#P5ND.+*[.FR8IFM0R[.*+R42&,R"RQW)av _m=7 "RR&Ils_F;8C
RRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVAv)q_gU4.RX.:NRDLRCDH"#RA"1aRH&RMo0CCHs'lCNo58IH0RE2&7R""RR&HCM0o'CsHolNC*5HU.4g2RR&"RW"&MRH0CCosl'HN5oC[2*.R"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05R5H+2R4*gU4.8,RCEb02&2RR""XRH&RMo0CCHs'lCNo5+5[4.2*2S;
SCSLo
HMRRRRRRRRRRRRSqA)v4_Ug..XR):Rq4vAn._1
RRRRRRRRRRRRRRRRbRRFRs0lRNb5R7Q=H>RMC_so*5.[R+48MFI0.FR*,[2R7q7)>R=RIDF_8N8s.54RI8FMR0FjR2, =hR>hR ,1R1)>R=Ra)1,R
RRRRRRRRRRRRRRRRRRRRRRRRRR RWRR=>I_s0CHM52B,Rp=iR>pRBi7,Rm254RR=>F_k0L.k#5.H,*4[+27,Rm25jRR=>F_k0L.k#5RH,.2*[2R;
RRRRRRRRRRRRRFRRks0_C.o5*R[2<F=RkL0_k5#.H*,.[I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co.+*[4<2R=kRF0k_L#H.5,[.*+R42IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRMSC8CRoMNCs0zCR.
(;RRRRRMSC8CRoMNCs0zCR.
c;RRRRCRM8oCCMsCN0Rdz.;
RR
RSRR-R-RMtCC0sNCER0CqR)vCRODRD#NRM8#CCDOD0RFOoHRsVFRv)qA_4n1Sc
zR.U:VRHRE5OFCHO_8IH0=ERRRc2oCCMsCN0
-SS-HRVGFRVsNROD4DRd(UU,CR#D0CORRFV0#sH0CN0R0MFRHLCMsoRC#oH0CCs8R
SREzO	RR:H5VRNs88I0H8ERR>4R.2oCCMsCN0
RRRRRRRRDzO	b:RsCFO#5#RB2pi
RSRRRRRLHCoMR
SRRRRRVRHRp5BiP'CCRM0NRM8BRpi=4R''02RE
CMSRRRRRRRRNRR8osC58N8s8IH04E-RI8FMR0F4R.2<N=R8C_so85N8HsI8-0E4FR8IFM0R24.;S
SRCRRMH8RVS;
S8CMRFbsO#C#RDkO	S;
RMRC8CRoMNCs0zCRO;E	
RRRR.SzgRR:VRFsHMRHRC58b_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
-S-RRQV58N8s8IH0>ERR24.RCMC8FR0RCOsNR0CI0sHCMRCNCLDR8NMR0FkbRk0CLMND#CRCODC0FRDo
HORRRRRRRRSjzdRH:RVNR58I8sHE80R4>R.o2RCsMCN
0CSR--VRHGVRFsODNDRU4dUR(,#CCDOF0RVsR0HN#00MCRFL0RCoHMRosCHC#0s
C8RRRRRRRRRRRRRRRRF_k0CHM52=R<R''4RCIEMNR58osC58N8s8IH04E-RI8FMR0F4R.2=2RHR#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=WI RERCM5_N8s5CoNs88I0H8ER-48MFI04FR.=2RRRH2CCD#R''j;R
RRRRRRCRSMo8RCsMCNR0Cz;dj
-S-RRQV58N8s8IH0<ER=.R42FRMRHIs0CCRMDNLCsRFR0FkbRk0CLMND#CRCODC0FRDoRHOM8CCCR8
SRRRRdSz4RR:H5VRNs88I0H8E=R<R24.RMoCC0sNCR
SRRRRRRRRRFRRkC0_M25HRR<=';4'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RW;R
RRRRRRCRSMo8RCsMCNR0Cz;d4
-S-RMtCC0sNCER0CqR)vCRODRD#NRM80-sH#00NCR#
RRRRRSRRzRd.:FRVsRR[H5MRI0H8Ek_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0SC
S0SN0LsHkR0CGbO_s#FbRRFVAv)q_gcjnRXc:NRDLRCDH"#R1q)epR="&sR#P5NDc+*[cFR8IFM0R[c*+R42&,R"RQW)av _m=7 "RR&Ils_F;8C
RRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVAv)q_gcjnRXc:NRDLRCDH"#RA"1aRH&RMo0CCHs'lCNo58IH0RE2&7R""RR&HCM0o'CsHolNC*5Hcnjg2RR&"RW"&MRH0CCosl'HN5oC[2*cR"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05R5H+2R4*gcjn8,RCEb02&2RR""XRH&RMo0CCHs'lCNo5+5[4c2*2S;
SCSLo
HMRRRRRRRRRRRRSqA)vj_cgcnXR):Rq4vAnc_1
RSRRRRRRRRRRFRbsl0RN5bR7=QR>MRH_osC5[c*+8dRF0IMF*Rc[R2,q)77RR=>D_FINs885R448MFI0jFR2 ,Rh>R=R, hR)11RR=>),1aRS
SS SWRR=>I_s0CHM52B,Rp=iR>pRBi7,Rm25dRR=>F_k0Lck#5RH,c+*[dR2,7.m52>R=R0Fk_#Lkc,5Hc+*[.R2,
SSSS57m4=2R>kRF0k_L#Hc5,[c*+,42R57mj=2R>kRF0k_L#Hc5,*Rc[;22
RRRRRRRRRRRRRRRR0Fk_osC5[c*2=R<R0Fk_#Lkc,5Hc2*[RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so*5c[2+4RR<=F_k0Lck#5cH,*4[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cco5*.[+2=R<R0Fk_#Lkc,5Hc+*[.I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Coc+*[d<2R=kRF0k_L#Hc5,[c*+Rd2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRMSC8CRoMNCs0zCRd
.;RRRRRMSC8CRoMNCs0zCR.
g;RRRRCRM8oCCMsCN0RUz.;S

RRRR-t-RCsMCNR0C0REC)RqvODCD#MRN8CR#D0CORoDFHVORF)sRq4vAng_1
dSzdRR:H5VROHEFOIC_HE80Rg=R2CRoMNCs0SC
SR--VRHGVRFsODNDRU4dUR(,#CCDOF0RVsR0HN#00MCRFL0RCoHMRosCHC#0s
C8SzRRORE	:VRHRN5R8I8sHE80R4>R4o2RCsMCN
0CRRRRRRRRz	OD:sRbF#OC#BR5p
i2SRRRRLRRCMoH
RSRRRRRRRHV5iBp'CCPMN0RMB8Rp=iRR''42ER0CSM
RRRRRRRRR8RNs5CoNs88I0H8ER-48MFI04FR4<2R=8RN_osC58N8s8IH04E-RI8FMR0F4;42
RSSRMRC8VRH;S
SCRM8bOsFCR##k	OD;R
SR8CMRMoCC0sNCORzE
	;RRRRSczdRV:RFHsRRRHM5b8C0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CSR--Q5VRNs88I0H8ERR>4R42M8CCRR0FONsC0ICRsCH0RNCMLRDCNRM8Fbk0kC0RMDNLCCR#D0CORoDFHRO
RRRRRSRRzRd6:VRHR85N8HsI8R0E>4R42CRoMNCs0SC
-V-RHVGRFOsRNRDD4UdU(#,RCODC0VRFRH0s#00NCFRM0CRLHRMosHCo#s0CCR8
RRRRRRRRRRRRRFRRkC0_M25HRR<='R4'IMECR85Ns5CoNs88I0H8ER-48MFI04FR4=2RRRH2CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R ERIC5MRNs8_CNo58I8sHE80-84RF0IMF4R42RR=HC2RDR#C';j'
RRRRRRRRMSC8CRoMNCs0zCRd
6;SR--Q5VRNs88I0H8E=R<R244RRMFI0sHCMRCNCLDRRFsFbk0kC0RMDNLCCR#D0CORoDFHMORCCC88S
RRRRRSnzdRH:RVNR58I8sHE80RR<=4R42oCCMsCN0
RSRRRRRRRRRRkRF0M_C5RH2<'=R4
';RRRRRRRRRRRRRRRRI_s0CHM52=R<R;W 
RRRRRRRRMSC8CRoMNCs0zCRd
n;SR--tCCMsCN0RC0ERv)qRDOCDN#RM08Rs#H-0CN0#R
RRRRRRzRSd:(RRsVFRH[RMIR5HE80_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNCS
SS0N0skHL0GCROs_bFRb#FAVR)_qv.UjcX:URRLDNCHDR#1R")peq=&"RRP#sNgD5*g[+RI8FMR0Fg+*[4&2RRR",Wa)Q m_v7" =RI&RsF_l8
C;RRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FAVR)_qv.UjcX:URRLDNCHDR#AR"1Ra"&MRH0CCosl'HN5oCI0H8E&2RR""7RH&RMo0CCHs'lCNo5.H*j2cUR"&RW&"RR0HMCsoC'NHlo[C5*Rg2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50E5+HRR*42.Ujc,CR8b20E2RR&"RX"&MRH0CCosl'HN5oC54[+22*g;S
SSoLCHRM
RRRRRRRRRSRRAv)q_c.jURXU:qR)vnA4_
1gSRRRRRRRRRRRRsbF0NRlb7R5Q>R=R_HMs5Cog+*[(FR8IFM0R[g*2q,R7R7)=D>RFNI_858s48jRF0IMF2Rj,hR RR=> Rh,1R1)=)>R1Ra,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRWRR >R=R0Is_5CMHR2,BRpi=B>RpRi,7(m52>R=R0Fk_#LkU,5HU+*[(R2,7nm52>R=R0Fk_#LkU,5HU+*[nR2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRm256RR=>F_k0LUk#5UH,*6[+27,Rm25cRR=>F_k0LUk#5UH,*c[+27,Rm25dRR=>F_k0LUk#5UH,*d[+2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR75R.2=F>RkL0_k5#UH*,U[2+.,mR75R42=F>RkL0_k5#UH*,U[2+4,mR75Rj2=F>RkL0_k5#UH*,U[R2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRQju52>R=R_HMs5Cog+*[UR2,75muj=2R>NRbs$H0_#LkU,5H[;22
RRRRRRRRRRRRRRRR0Fk_osC5[g*2=R<R0Fk_#LkU,5HU2*[RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so*5g[2+4RR<=F_k0LUk#5UH,*4[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cgo5*.[+2=R<R0Fk_#LkU,5HU+*[.I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cog+*[d<2R=kRF0k_L#HU5,[U*+Rd2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5[g*+Rc2<F=RkL0_k5#UH*,U[2+cRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so*5g[2+6RR<=F_k0LUk#5UH,*6[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cgo5*n[+2=R<R0Fk_#LkU,5HU+*[nI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cog+*[(<2R=kRF0k_L#HU5,[U*+R(2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5[g*+RU2<b=RN0sH$k_L#HU5,R[2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRMSC8CRoMNCs0zCRd
(;RRRRRMSC8CRoMNCs0zCRd
c;RRRRCRM8oCCMsCN0Rdzd;S

RRRR-t-RCsMCNR0C0REC)RqvODCD#MRN8CR#D0CORoDFHVORF)sRq4vAn4_1Uz
Sd:URRRHV5FOEH_OCI0H8ERR=4RU2oCCMsCN0
-SS-HRVGFRVsNROD4DRd(UU,CR#D0CORRFV0#sH0CN0R0MFRHLCMsoRC#oH0CCs8R
SREzO	RR:H5VRR8N8s8IH0>ERRR4j2CRoMNCs0RC
RRRRRzRRO:D	RFbsO#C#Rp5BiS2
RRRRRCRLo
HMSRRRRRRRH5VRB'piCMPC0MRN8pRBiRR='24'RC0EMR
SRRRRRRRRRsN8CNo58I8sHE80-84RF0IMFjR42=R<R_N8s5CoNs88I0H8ER-48MFI04FRj
2;SRSRR8CMR;HV
CSSMb8RsCFO#k#RO;D	
RSRCRM8oCCMsCN0REzO	R;
RSRRzRdg:FRVsRRHH5MR80CbEk_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0SC
-Q-RVNR58I8sHE80R4>RjM2RCRC80OFRs0CNCsRIHR0CCLMNDNCRMF8Rkk0b0MRCNCLDRD#CCRO0DHFoOR
RRRRRRzRSc:jRRRHV58N8s8IH0>ERR24jRMoCC0sNC-
S-HRVGFRVsNROD4DRd(UU,CR#D0CORRFV0#sH0CN0R0MFRHLCMsoRC#oH0CCs8R
RRRRRRRRRRRRRRkRF0M_C5RH2<'=R4I'RERCM5sN8CNo58I8sHE80-84RF0IMFjR42RR=HC2RDR#C';j'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RWRCIEMNR58C_so85N8HsI8-0E4FR8IFM0R24jRH=R2DRC#'CRj
';RRRRRRRRS8CMRMoCC0sNCcRzjS;
-Q-RVNR58I8sHE80RR<=4Rj2MIFRsCH0RNCMLRDCFFsRkk0b0MRCNCLDRD#CCRO0DHFoOCRMC88C
RRSRSRRzRc4:VRHR85N8HsI8R0E<4=Rjo2RCsMCN
0CSRRRRRRRRRRRR0Fk_5CMH<2R=4R''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=W
 ;RRRRRRRRS8CMRMoCC0sNCcRz4S;
-t-RCsMCNR0C0REC)RqvODCD#MRN8sR0H0-#N#0C
RRRRRRRRcSz.RR:VRFs[MRHRH5I8_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
SSSNs00H0LkCORG_FbsbF#RV)RAq4v_jX.c4:nRRLDNCHDR#1R")peq=&"RRP#sN4D5U+*[48URF0IMFUR4*4[+2RR&"W,R) Qa_7vm R="&sRI_8lFCR;
RRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)RAq4v_jX.c4:nRRLDNCHDR#AR"1Ra"&MRH0CCosl'HN5oCI0H8E&2RR""7RH&RMo0CCHs'lCNo54H*j2.cR"&RW&"RR0HMCsoC'NHlo[C5*24UR"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05R5H+2R4*.4jc8,RCEb02&2RR""XRH&RMo0CCHs'lCNo5+5[442*U
2;SLSSCMoH
RRRRRRRRRRRR)SAq4v_jX.c4:nRRv)qA_4n1
4URRRRRRRRRRRRRRRRRFRbsl0RN5bR7=QR>MRH_osC5*4U[6+4RI8FMR0F4[U*2q,R7R7)=D>RFNI_858sgFR8IFM0R,j2RR h= >Rh1,R1=)R>1R)a
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRW= R>sRI0M_C5,H2RiBpRR=>B,piR57m4R62=F>RkL0_kn#454H,n+*[4,62R57m4Rc2=F>RkL0_kn#454H,n+*[4,c2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7524dRR=>F_k0L4k#n,5H4[n*+24d,mR7524.RR=>F_k0L4k#n,5H4[n*+24.,mR75244RR=>F_k0L4k#n,5H4[n*+244,RR
RRRRRRRRRRRRRRRRRRRRRRRRR7RRmj542>R=R0Fk_#Lk4Hn5,*4n[j+427,Rm25gRR=>F_k0L4k#n,5H4[n*+,g2R57mU=2R>kRF0k_L#54nHn,4*U[+2R,
RRRRRRRRRRRRRRRRRRRRRRRRR7RRm25(RR=>F_k0L4k#n,5H4[n*+,(2R57mn=2R>kRF0k_L#54nHn,4*n[+27,Rm256RR=>F_k0L4k#n,5H4[n*+,62
SSSRRRR7cm52>R=R0Fk_#Lk4Hn5,*4n[2+c,mR75Rd2=F>RkL0_kn#454H,n+*[dR2,7.m52>R=R0Fk_#Lk4Hn5,*4n[2+.,R
RRRRRRRRRRRRRRRRRRRRRRRRRRmR75R42=F>RkL0_kn#454H,n+*[4R2,7jm52>R=R0Fk_#Lk4Hn5,*4n[R2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRu7QRR=>HsM_C4o5U+*[48(RF0IMFUR4*4[+n
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRR75mu4=2R>NRbs$H0_#Lk4Hn5,[.*+,42Ru7m5Rj2=b>RN0sH$k_L#54nH*,.[;22
RRRRRRRRRRRRRRRR0Fk_osC5*4U[<2R=kRF0k_L#54nHn,4*R[2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[2+4RR<=F_k0L4k#n,5H4[n*+R42IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[2+.RR<=F_k0L4k#n,5H4[n*+R.2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[2+dRR<=F_k0L4k#n,5H4[n*+Rd2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[2+cRR<=F_k0L4k#n,5H4[n*+Rc2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[2+6RR<=F_k0L4k#n,5H4[n*+R62IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[2+nRR<=F_k0L4k#n,5H4[n*+Rn2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[2+(RR<=F_k0L4k#n,5H4[n*+R(2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[2+URR<=F_k0L4k#n,5H4[n*+RU2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[2+gRR<=F_k0L4k#n,5H4[n*+Rg2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[j+42=R<R0Fk_#Lk4Hn5,*4n[j+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[4R42<F=RkL0_kn#454H,n+*[4R42IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[.+42=R<R0Fk_#Lk4Hn5,*4n[.+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[4Rd2<F=RkL0_kn#454H,n+*[4Rd2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[c+42=R<R0Fk_#Lk4Hn5,*4n[c+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[4R62<F=RkL0_kn#454H,n+*[4R62IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[n+42=R<RsbNH_0$L4k#n,5H.2*[RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*4[+(<2R=NRbs$H0_#Lk4Hn5,[.*+R42IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRMSC8CRoMNCs0zCRc
.;RRRRRMSC8CRoMNCs0zCRd
g;RRRRCRM8oCCMsCN0RUzd;S

RRRR-t-RCsMCNR0C0REC)RqvODCD#MRN8CR#D0CORoDFHVORF)sRq4vAnd_1nz
Sc:dRRRHV5FOEH_OCI0H8ERR=dRn2oCCMsCN0
-SS-HRVGFRVsNROD4DRd(UU,CR#D0CORRFV0#sH0CN0R0MFRHLCMsoRC#oH0CCs8R
SREzO	RR:H5VRR8N8s8IH0>ERR2gRRMoCC0sNCR
SRzRRO:D	RFbsO#C#Rp5BiS2
SLRRCMoH
RSSRVRHRp5BiP'CCRM0NRM8BRpi=4R''02RE
CMSRSRRRRRNC8so85N8HsI8-0E4FR8IFM0RRg2<N=R8C_so85N8HsI8-0E4FR8IFM0R;g2
RSSRMRC8VRH;S
SCRM8bOsFCR##k	OD;R
SR8CMRMoCC0sNCORzE
	;SRRRRczcRV:RFHsRRRHM5b8C0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CSR--Q5VRNs88I0H8ERR>gM2RCRC80OFRs0CNCsRIHR0CCLMNDNCRMF8Rkk0b0MRCNCLDRD#CCRO0DHFoOS
SS6zcRH:RVNR58I8sHE80Rg>R2CRoMNCs0SC
-V-RHVGRFOsRNRDD4UdU(#,RCODC0VRFRH0s#00NCFRM0CRLHRMosHCo#s0CCS8
SFSSkC0_M25HRR<='R4'IMECR85Ns5CoNs88I0H8ER-48MFI0gFR2RR=HC2RDR#C';j'
SSSS0Is_5CMH<2R= RWRCIEMNR58C_so85N8HsI8-0E4FR8IFM0RRg2=2RHR#CDCjR''S;
SMSC8CRoMNCs0zCRc
6;SR--Q5VRNs88I0H8E=R<RRg2MIFRsCH0RNCMLRDCFFsRkk0b0MRCNCLDRD#CCRO0DHFoOCRMC88C
SSSzRcn:VRHR85N8HsI8R0E<g=R2CRoMNCs0SC
SFSSkC0_M25HRR<=';4'
SSSS0Is_5CMH<2R= RW;S
SS8CMRMoCC0sNCcRznS;
-t-RCsMCNR0C0REC)RqvODCD#MRN8sR0H0-#N#0C
SSSzRc(:FRVsRR[H5MRI0H8Ek_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0SC
S0SN0LsHkR0CGbO_s#FbRRFVAv)q_.64XRd.:NRDLRCDH"#R1q)epR="&sR#P5NDd[n*+Rdn8MFI0dFRn+*[4&2RRR",Wa)Q m_v7" =RI&RsF_l8
C;RRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FAVR)_qv6X4.d:.RRLDNCHDR#AR"1Ra"&MRH0CCosl'HN5oCI0H8E&2RR""7RH&RMo0CCHs'lCNo56H*4R.2&WR""RR&HCM0o'CsHolNC*5[dRn2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50E5+HRR*426,4.Rb8C02E2R"&RX&"RR0HMCsoC'NHlo5C5[2+4*2dn;S
SSoLCHRM
RRRRRRRRRRRRRRRRRRRRRRRRRqA)v4_6..XdR):Rq4vAnd_1nR
RRRRRRRRRRRRRRRRRRRRRRRRRRFRbsl0RN5bR7=QR>MRH_osC5*dn[4+dRI8FMR0Fd[n*2q,R7R7)=F>DI8_N8Us5RI8FMR0FjR2, =hR>hR ,1R1)>R=Ra)1,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRW= R>sRI0M_C5,H2RiBpRR=>B,piR57mdR42=F>RkL0_k.#d5dH,.+*[d,42R57mdRj2=F>RkL0_k.#d5dH,.+*[d,j2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRmg5.2>R=R0Fk_#LkdH.5,*d.[g+.27,RmU5.2>R=R0Fk_#LkdH.5,*d.[U+.27,Rm(5.2>R=R0Fk_#LkdH.5,*d.[(+.2R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR57m.Rn2=F>RkL0_k.#d5dH,.+*[.,n2R57m.R62=F>RkL0_k.#d5dH,.+*[.,62R57m.Rc2=F>RkL0_k.#d5dH,.+*[.,c2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRmd5.2>R=R0Fk_#LkdH.5,*d.[d+.27,Rm.5.2>R=R0Fk_#LkdH.5,*d.[.+.27,Rm45.2>R=R0Fk_#LkdH.5,*d.[4+.2R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR57m.Rj2=F>RkL0_k.#d5dH,.+*[.,j2R57m4Rg2=F>RkL0_k.#d5dH,.+*[4,g2R57m4RU2=F>RkL0_k.#d5dH,.+*[4,U2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRm(542>R=R0Fk_#LkdH.5,*d.[(+427,Rmn542>R=R0Fk_#LkdH.5,*d.[n+427,Rm6542>R=R0Fk_#LkdH.5,*d.[6+42R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR57m4Rc2=F>RkL0_k.#d5dH,.+*[4,c2R57m4Rd2=F>RkL0_k.#d5dH,.+*[4,d2R57m4R.2=F>RkL0_k.#d5dH,.+*[4,.2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR74m54=2R>kRF0k_L#5d.H.,d*4[+4R2,74m5j=2R>kRF0k_L#5d.H.,d*4[+jR2,7gm52>R=R0Fk_#LkdH.5,*d.[2+g,RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR57mU=2R>kRF0k_L#5d.H.,d*U[+27,Rm25(RR=>F_k0Ldk#.,5Hd[.*+,(2R57mn=2R>kRF0k_L#5d.H.,d*n[+2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR75R62=F>RkL0_k.#d5dH,.+*[6R2,7cm52>R=R0Fk_#LkdH.5,*d.[2+c,mR75Rd2=F>RkL0_k.#d5dH,.+*[dR2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRm25.RR=>F_k0Ldk#.,5Hd[.*+,.2R57m4=2R>kRF0k_L#5d.H.,d*4[+27,Rm25jRR=>F_k0Ldk#.,5Hd[.*2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRQR7u>R=R_HMs5Cod[n*+Rd68MFI0dFRn+*[d,.2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRmdu52>R=RsbNH_0$Ldk#.,5Hc+*[dR2,75mu.=2R>NRbs$H0_#LkdH.5,[c*+,.2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRm4u52>R=RsbNH_0$Ldk#.,5Hc+*[4R2,75muj=2R>NRbs$H0_#LkdH.5,[c*2
2;RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*R[2<F=RkL0_k.#d5dH,.2*[RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*+R42<F=RkL0_k.#d5dH,.+*[4I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*.[+2=R<R0Fk_#LkdH.5,*d.[2+.RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*+Rd2<F=RkL0_k.#d5dH,.+*[dI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*c[+2=R<R0Fk_#LkdH.5,*d.[2+cRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*+R62<F=RkL0_k.#d5dH,.+*[6I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*n[+2=R<R0Fk_#LkdH.5,*d.[2+nRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*+R(2<F=RkL0_k.#d5dH,.+*[(I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*U[+2=R<R0Fk_#LkdH.5,*d.[2+URCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*+Rg2<F=RkL0_k.#d5dH,.+*[gI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*4[+j<2R=kRF0k_L#5d.H.,d*4[+jI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*4[+4<2R=kRF0k_L#5d.H.,d*4[+4I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*4[+.<2R=kRF0k_L#5d.H.,d*4[+.I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*4[+d<2R=kRF0k_L#5d.H.,d*4[+dI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*4[+c<2R=kRF0k_L#5d.H.,d*4[+cI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*4[+6<2R=kRF0k_L#5d.H.,d*4[+6I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*4[+n<2R=kRF0k_L#5d.H.,d*4[+nI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*4[+(<2R=kRF0k_L#5d.H.,d*4[+(I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*4[+U<2R=kRF0k_L#5d.H.,d*4[+UI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*4[+g<2R=kRF0k_L#5d.H.,d*4[+gI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*.[+j<2R=kRF0k_L#5d.H.,d*.[+jI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*.[+4<2R=kRF0k_L#5d.H.,d*.[+4I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*.[+.<2R=kRF0k_L#5d.H.,d*.[+.I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*.[+d<2R=kRF0k_L#5d.H.,d*.[+dI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*.[+c<2R=kRF0k_L#5d.H.,d*.[+cI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*.[+6<2R=kRF0k_L#5d.H.,d*.[+6I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*.[+n<2R=kRF0k_L#5d.H.,d*.[+nI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*.[+(<2R=kRF0k_L#5d.H.,d*.[+(I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*.[+U<2R=kRF0k_L#5d.H.,d*.[+UI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*.[+g<2R=kRF0k_L#5d.H.,d*.[+gI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*d[+j<2R=kRF0k_L#5d.H.,d*d[+jI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*d[+4<2R=kRF0k_L#5d.H.,d*d[+4I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*d[+.<2R=NRbs$H0_#LkdH.5,[c*2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[d+d2=R<RsbNH_0$Ldk#.,5Hc+*[4I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*d[+c<2R=NRbs$H0_#LkdH.5,[c*+R.2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[dR62<b=RN0sH$k_L#5d.H*,c[2+dRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;S
SS8CMRMoCC0sNCcRz(S;
S8CMRMoCC0sNCcRzcS;
CRM8oCCMsCN0Rdzc;C

MN8RsHOE00COkRsCLODF	N_sl
;
NEsOHO0C0CksR_MFsOI_E	CORRFV)hqv_R)WHV#
k0MOHRFMVOkM_HHM0R5L:FRLFNDCMs2RCs0kM0R#soHMR
H#LHCoMR
RH5VRL02RE
CMRRRRskC0s"M5hsFRC/N8I0sHCFROMHVDOO0RE	CO3HR1lNkD0MHFR#lHlON0EFRb#L#HD!CR!;"2
CRRD
#CRRRRskC0s"M5'_MFsOI_E	CO'#RHRC0ERl#NC#RNRD'LF_O	s'NlRsVFRM#HoRDCb0FsRv)q#;"2
CRRMH8RVC;
MV8Rk_MOH0MH;0
N0LsHkR0CoCCMsFN0sC_sb0FsR#:R0MsHo-;
-0N0skHL0oCRCsMCNs0F_bsCFRs0FMVRFI_s_COEO:	RRONsECH0Os0kC#RHRMVkOM_HHN058_8ss2Co;k
VMHO0F#MR0MsHoD.#PR5N:0R#soHM2CRs0MksR8#0_oDFHPO_CFO0s#RH
sPNHDNLCDR#PRR:#_08DHFoOC_POs0F5EN'H-oENF'DIFR8IFM0R;j2
sPNHDNLCRRH:MRH0CCosL;
CMoH
VRRFHsRRRHMjFR0RP#D'oEHEFRDFRb
RHRRVNR55EN'H-oEH=2RR''42ER0CSM
RDR#P25HRR:=';4'
DSC#SC
RDR#P25HRR:=';j'
MSC8VRH;R
RCRM8DbFF;R
RskC0s#MRD
P;CRM8#H0sM#o.D
P;VOkM0MHFRP#D.s#0H5MoNRR:#_08DHFoOC_POs0F2CRs0MksRs#0HRMoHP#
NNsHLRDC#RR:#H0sMNo5'oEHE'-ND+FI4FR8IFM0R;42
sPNHDNLCRRH:MRH0CCosL;
CMoH
VRRFHsRRRHMNF'DIFR0REN'HRoEDbFF
RRRRRHV5HN52RR='24'RC0EMR
SRH#5-DN'F4I+2=R:R''4;C
SD
#CS#RR5NH-'IDF+R42:'=Rj
';S8CMR;HV
CRRMD8RF;Fb
sRRCs0kM;R#
8CMRP#D.s#0H;Mo
0N0skHL0GCROs_bFRb#:0R#soHM;-
-O#FM00NMRP#sN:DRR8#0_oDFHPO_CFO0sH5I8-0E4FR8IFM0RRj2:#=R0MsHoD.#P#5s0N_80;N2
R--LHCoMDRLFRO	sRNlHDlbCMlC0HN0F#MRHNoMDV#
k0MOHRFMo_C0OHEFOIC_HE8058IH0:ERR0HMCsoC2CRs0MksR0HMCsoCR
H#PHNsNCLDRDPNRH:RMo0CC:sR=;Rj
sPNHDNLCHR8P,d.RP8H4Rn,8UHP,HR8PRc,8.HP,HR8P:4RR0HMCsoC;C
Lo
HMRHR8PRd.:5=RI0H8E2-4/;dn
8RRHnP4RR:=58IH04E-2U/4;R
R8UHPRR:=58IH04E-2;/g
8RRHRPc:5=RI0H8E2-4/
c;RHR8P:.R=IR5HE80-/42.R;
RP8H4=R:RH5I8-0E4
2;RVRHRH58P>4RRRj20MEC
RRRRDPNRR:=PRND+;R4
CRRMH8RVR;
RRHV5P8H.RR>j02RE
CMRRRRPRND:P=RN+DRR
4;RMRC8VRH;R
RH5VR8cHPRj>R2ER0CRM
RPRRN:DR=NRPDRR+4R;
R8CMR;HV
HRRV8R5HRPU>2RjRC0EMR
RRNRPD=R:RDPNR4+R;R
RCRM8H
V;RVRHRH58PR4n>2RjRC0EMR
RRNRPD=R:RDPNR4+R;R
RCRM8H
V;-R-RH5VR8dHP.RR>j02RE
CM-R-RRNRPD=R:RDPNR4+R;-
-RMRC8VRH;R
RH5VRPRND>2R.RC0EMRR
RsRRCs0kM.R5RR**PRND+RR.*5*RPRND-2Rd2R;
R#CDCR
RRCRs0MksRR5.*P*RN;D2
CRRMH8RVC;
Mo8RCO0_EOFHCH_I8;0E
MVkOF0HMCRo0E_OFCHO_b8C08E5CEb0RH:RMo0CCRs2skC0sHMRMo0CCHsR#N
PsLHND8CR_FOEH_OC80CbERR:HCM0oRCs:j=R;C
Lo
HMRVRHRC58bR0E>4RUgR.20MEC
RRRRO8_EOFHCC_8bR0E:4=RncdU;R
RCHD#V8R5CEb0RR<=U.4gR8NMRb8C0>ERRgcjnRR20MEC
RRRRO8_EOFHCC_8bR0E:U=R4;g.
CRRDV#HRC58bR0E<c=RjRgnNRM880CbERR>.Ujc2ER0CRM
R8RR_FOEH_OC80CbE=R:RgcjnR;
R#CDH5VR80CbE=R<Rc.jUMRN8CR8bR0E>jR4.2cRRC0EMR
RR_R8OHEFO8C_CEb0RR:=.Ujc;R
RCHD#V8R5CEb0RR<=4cj.R8NMRb8C0>ERR.642ER0CRM
R8RR_FOEH_OC80CbE=R:R.4jcR;
R#CDH5VR80CbE=R<R.642ER0CRM
R8RR_FOEH_OC80CbE=R:R.64;R
RCRM8H
V;RCRs0MksRO8_EOFHCC_8b;0E
8CMR0oC_FOEH_OC80CbEV;
k0MOHRFMo_C0I0H8EF_l85_UOHEFOIC_8RR:HCM0o2CsR0sCkRsMHCM0oRCsHP#
NNsHLRDCI0H8EF_l8R_U:MRH0CCosL;
CMoH
HRRVOR5EOFHC8_IRU>R2ER0CRM
RIRRHE80_8lF_:UR=EROFCHO_RI8-OR5EOFHC8_IR8lFR;U2
CRRD
#CRRRRI0H8EF_l8R_U:O=REOFHC8_I;R
RCRM8H
V;RCRs0MksR8IH0lE_FU8_;M
C8CRo0H_I8_0El_F8U
;
O#FM00NMROI_EOFHCH_I8R0E:MRH0CCos=R:R0oC_FOEH_OCI0H8EH5I820E;F
OMN#0MI0R_FOEH_OC80CbERR:HCM0oRCs:4=RncdU/0oC_8IH0lE_FU8_5OI_EOFHCH_I820E;F
OMN#0M80R_FOEH_OC80CbERR:HCM0oRCs:o=RCO0_EOFHCC_8b50E80CbE
2;O#FM00NMRO8_EOFHCH_I8R0E:MRH0CCos=R:Rn54d/Uc8E_OFCHO_b8C0RE2+5R54Undc_/8OHEFO8C_CEb02RR/U
2;
MVkOF0HMCRo0k_MlC_OD5D#I:8RR0HMCsoC;FOEH_OCI:8RR0HMCsoC2CRs0MksR0HMCsoCR
H#PHNsNCLDRlMk_DOCD:#RR0HMCsoC;C
Lo
HMRkRMlC_ODRD#:5=RI48-2E/OFCHO_RI8+;R4
sRRCs0kMkRMlC_OD;D#
8CMR0oC_lMk_DOCD
#;
MVkOF0HMCRo0H_#xIC5M:ORR0HMCsoC;MR8ORR:HCM0o2CsR0sCkRsMHCM0oRCsHL#
CMoH
RRRskC0sIMRM*ORRO8M;M
C8CRo0H_#x
C;
MVkOF0HMCRo0F_LF5D88H_#x:CRR0HMCsoC;_RI#CHxRH:RMo0CCRs;8I_ORH:RMo0CCRs;II_ORH:RMo0CCRs2skC0sHMRMo0CCHsR#C
Lo
HMH5VR8H_#x<CR=_RI#CHx2ER0CRM
R0sCkRsM8I_O;D
C#RC
R0sCkRsMII_O;M
C8VRH;M
C8CRo0F_LF;D8
MVkOF0HMCRo0M_C8C_8b50E#CHxRH:RMo0CC;sRRb8C0:ERR0HMCsoC2CRs0MksR0HMCsoCR
H#PHNsNCLDRMlH_x#HCRR:HCM0oRCs:j=R;C
Lo
HMRHRlMH_#x:CR=CR8b;0E
HRRV#R5HRxC<CR8b20ERC0EMR
RRHRlMH_#x:CR=HR#x
C;RMRC8VRH;R
RskC0slMRH#M_H;xC
8CMR0oC_8CM_b8C0
E;
MOF#M0N0EROFCHO_8IH0:ERR0HMCsoCRR:=o_C0LDFF8C5o0H_#xoC5CM0_kOl_C#DD58IH0RE,8E_OFCHO_8IH0,E2o_C0M_klODCD#C58b,0ERO8_EOFHCC_8b20E2R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRo_C0#CHx50oC_lMk_DOCDI#5HE80,_RIOHEFOIC_HE802C,o0k_MlC_OD5D#80CbEI,R_FOEH_OC80CbE,22
SSSSSSSSSSSRO8_EOFHCH_I8,0EROI_EOFHCH_I820E;F
OMN#0MI0RHE80_lMk_DOCD:#RR0HMCsoCRR:=o_C0LDFF8C5o0H_#xoC5CM0_kOl_C#DD58IH0RE,8E_OFCHO_8IH0,E2o_C0M_klODCD#C58b,0ERO8_EOFHCC_8b20E2R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRoRRC#0_H5xCo_C0M_klODCD#H5I8,0EROI_EOFHCH_I820E,0oC_lMk_DOCD8#5CEb0,_RIOHEFO8C_CEb02
2,SSSSSSSSSRSSR5RRI0H8E2-4/O8_EOFHCH_I8,0ERH5I8-0E4I2/_FOEH_OCI0H8E+2RR
4;O#FM00NMRb8C0ME_kOl_C#DDRH:RMo0CC:sR=CRo0F_LF5D8o_C0#CHx50oC_lMk_DOCDI#5HE80,_R8OHEFOIC_HE802C,o0k_MlC_OD5D#80CbE8,R_FOEH_OC80CbE,22
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRo_C0#CHx50oC_lMk_DOCDI#5HE80,_RIOHEFOIC_HE802C,o0k_MlC_OD5D#80CbEI,R_FOEH_OC80CbE,22
SSSSSSSSRSSR8R5CEb0-/428E_OFCHO_b8C0RE,5b8C04E-2_/IOHEFO8C_CEb02RR+4R;S
MOF#M0N0CRxs:FRR8#0_oDFHPO_CFO0sE5OFCHO_8IH0IE*HE80_lMk_DOCDI#-HE80-84RF0IMF2RjRR:=5EF0CRs#='>Rj;'2
MOF#M0N0sR#P_ND#RDP:0R#8F_Do_HOP0COFOs5EOFHCH_I8*0EI0H8Ek_MlC_OD-D#4FR8IFM0RRj2:x=RCRsF&0R#soHM.P#D50s#_08NN
2;O#FM00NMRP#sN:DRRs#0H5MoOHEFOIC_HE80*8IH0ME_kOl_C#DDRI8FMR0F4:2R=DR#P0.#soHM5P#sN#D_D;P2
#--HNoMDV#RFMsRFDM-#bENCL8RD	FORlsN#$
0bFCRkL0_k_#40C$bRRH#NNss$8R5CEb0_lMk_DOCD4#-RI8FMR0FjI,RHE80_lMk_DOCD4#-RI8FMR0FjF2RV0R#8F_Do;HO
o#HMRNDF_k0L4k#RF:RkL0_k_#40C$b;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFV80FkRM5HbRk000FRs#H-0CN0#02
$RbCF_k0L.k#_b0$C#RHRsNsN5$R80CbEk_MlC_OD-D#4FR8IFM0RRj,.H*I8_0EM_klODCD#R+48MFI0jFR2VRFR8#0_oDFH
O;#MHoNFDRkL0_kR#.:kRF0k_L#0._$;bCRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$F8VRFRk05bHMk00RFsR0H0-#N#0C2$
0bFCRkL0_k_#c0C$bRRH#NNss$8R5CEb0_lMk_DOCD4#-RI8FMR0Fjc,R*8IH0ME_kOl_C#DD+8dRF0IMF2RjRRFV#_08DHFoO#;
HNoMDkRF0k_L#:cRR0Fk_#Lkc$_0bRC;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RVFR8k50RHkMb0FR0RH0s-N#002C#
b0$CkRF0k_L#0U_$RbCHN#Rs$sNRC58b_0EM_klODCD#R-48MFI0jFR,*RUI0H8Ek_MlC_OD+D#(FR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNR0Fk_#LkURR:F_k0LUk#_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFRk8F0HR5M0bkRR0F0-sH#00NC
#20C$bRsbNH_0$LUk#_b0$C#RHRsNsN5$R80CbEk_MlC_OD-D#4FR8IFM0RRj,I0H8Ek_MlC_OD-D#4FR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNRsbNH_0$LUk#Rb:RN0sH$k_L#0U_$;bCRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFRk8F0HR5M0bkRR0F0-sH#00NC
#20C$bR0Fk_#Lk40n_$RbCHN#Rs$sNRC58b_0EM_klODCD#R-48MFI0jFR,nR4*8IH0ME_kOl_C#DD+R468MFI0jFR2VRFR8#0_oDFH
O;#MHoNFDRkL0_kn#4RF:RkL0_kn#4_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFRk8F0HR5M0bkRR0F0-sH#00NC
#20C$bRsbNH_0$L4k#n$_0bHCR#sRNsRN$5b8C0ME_kOl_C#DD-84RF0IMF,RjRI.*HE80_lMk_DOCD4#+RI8FMR0FjF2RV0R#8F_Do;HO
o#HMRNDbHNs0L$_kn#4Rb:RN0sH$k_L#_4n0C$b;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFV80FkRM5HbRk000FRs#H-0CN0#02
$RbCF_k0Ldk#.$_0bHCR#sRNsRN$5b8C0ME_kOl_C#DD-84RF0IMF,RjR*d.I0H8Ek_MlC_OD+D#d84RF0IMF2RjRRFV#_08DHFoO#;
HNoMDkRF0k_L#Rd.:kRF0k_L#_d.0C$b;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFV80FkRM5HbRk000FRs#H-0CN0#02
$RbCbHNs0L$_k.#d_b0$C#RHRsNsN5$R80CbEk_MlC_OD-D#4FR8IFM0RRj,cH*I8_0EM_klODCD#R+d8MFI0jFR2VRFR8#0_oDFH
O;#MHoNbDRN0sH$k_L#Rd.:NRbs$H0_#Lkd0._$;bCRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$F8VRFRk05bHMk00RFsR0H0-#N#0C2H
#oDMNR0Fk_RCM:0R#8F_Do_HOP0COF8s5CEb0_lMk_DOCD4#-RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-C-RMDNLCV#RF0sRs#H-0CN0#H
#oDMNR0Is_RCM:0R#8F_Do_HOP0COF8s5CEb0_lMk_DOCD4#-RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-I-RsCH0RNCML#DCRsVFROCNEFRsIVRFRv)qRDOCD##
HNoMDMRH_osCR#:R0D8_FOoH_OPC05FsI0H8E6+dRI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RCk#8FR0RosCHC#0sQR7h#R
HNoMDkRF0C_soRR:#_08DHFoOC_POs0F58IH0dE+6FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RCk#8FR0RosCHC#0smR7z#a
HNoMD8RN_osCR#:R0D8_FOoH_OPC05FsNs88I0H8ER-48MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--k8#CRR0FsHCo#s0CR7q7)H
#oDMNRIDF_8N8sRR:#_08DHFoOC_POs0F5R4d8MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--Ns88R0LH#MRHbRk00)FRqOvRC#DDRR5cL#H0RJsCkCHs8#2
HNoMD8RNsRCo:0R#8F_Do_HOP0COFNs58I8sHE80-84RF0IMF2Rj;-R-RR0FsHCo#s0CRC0ERD#CCRO0#MHoNFDRVsR0HN#00-C
-MRC8DRLFRO	sRNlHDlbCMlC0HN0F#MRHNoMDN#
0H0sLCk0Rs\3NFl_VCV#0:\RRs#0H;Mo
C
Lo
HMRRR
R-RR-VRQR8N8s8IH0<ERRFOEH_OCI0H8E#RN#MHoR''jRR0Fk#MkCL8RH
0#RRRRzRjR:VRHR85N8HsI8R0E=2R4RMoCC0sNCR
SRDRRFNI_8R8s<"=Rjjjjjjjjjjjjj&"RR_N8s5Coj
2;S8CMRMoCC0sNCjRz;R
RR4RzRRR:H5VRNs88I0H8ERR=.o2RCsMCN
0CSRRRRIDF_8N8s=R<Rj"jjjjjjjjjjRj"&8RN_osC584RF0IMF2Rj;C
SMo8RCsMCNR0Cz
4;RRRRzR.R:VRHR85N8HsI8R0E=2RdRMoCC0sNCR
SRDRRFNI_8R8s<"=Rjjjjjjjjj"jjRN&R8C_soR5.8MFI0jFR2S;
CRM8oCCMsCN0R;z.
RRRRRzdRH:RVNR58I8sHE80Rc=R2CRoMNCs0SC
RRRRD_FINs88RR<="jjjjjjjj"jjRN&R8C_soR5d8MFI0jFR2S;
CRM8oCCMsCN0R;zd
RRRRRzcRH:RVNR58I8sHE80R6=R2CRoMNCs0SC
RRRRD_FINs88RR<="jjjjjjjjRj"&8RN_osC58cRF0IMF2Rj;C
SMo8RCsMCNR0Cz
c;RRRRzR6R:VRHR85N8HsI8R0E=2RnRMoCC0sNCR
SRDRRFNI_8R8s<"=Rjjjjjjjj"RR&Ns8_C6o5RI8FMR0Fj
2;S8CMRMoCC0sNC6Rz;R
RRnRzRRR:H5VRNs88I0H8ERR=(o2RCsMCN
0CSRRRRIDF_8N8s=R<Rj"jjjjjj&"RR_N8s5ConFR8IFM0R;j2
MSC8CRoMNCs0zCRnR;
RzRR(:RRRRHV58N8s8IH0=ERRRU2oCCMsCN0
RSRRFRDI8_N8<sR=jR"jjjjj&"RR_N8s5Co(FR8IFM0R;j2
MSC8CRoMNCs0zCR(R;
RzRRU:RRRRHV58N8s8IH0=ERRRg2oCCMsCN0
RSRRFRDI8_N8<sR=jR"jjjj"RR&Ns8_CUo5RI8FMR0Fj
2;S8CMRMoCC0sNCURz;R
RRgRzRRR:H5VRNs88I0H8ERR=4Rj2oCCMsCN0
RSRRFRDI8_N8<sR=jR"j"jjRN&R8C_soR5g8MFI0jFR2S;
CRM8oCCMsCN0R;zg
RRRRjz4RRR:H5VRNs88I0H8ERR=4R42oCCMsCN0
RSRRFRDI8_N8<sR=jR"jRj"&8RN_osC5R4j8MFI0jFR2S;
CRM8oCCMsCN0Rjz4;R
RR4Rz4:RRRRHV58N8s8IH0=ERR24.RMoCC0sNCR
SRDRRFNI_8R8s<"=RjRj"&8RN_osC5R448MFI0jFR2S;
CRM8oCCMsCN0R4z4;R
RR4Rz.:RRRRHV58N8s8IH0=ERR24dRMoCC0sNCR
SRDRRFNI_8R8s<'=Rj&'RR_N8s5Co48.RF0IMF2Rj;C
SMo8RCsMCNR0Cz;4.
RRRRdz4RRR:H5VRNs88I0H8ERR>4Rd2oCCMsCN0
RSRRFRDI8_N8<sR=8RN_osC5R4d8MFI0jFR2S;
CRM8oCCMsCN0Rdz4;R

R-RR-VRQRH58MC_sos2RC#oH0RCs7RQhkM#HopRBiR
RR4Rzc:RRRRHV5M8H_osC2CRoMNCs0RC
RRRRRbRRsCFO#5#RB,piRh7Q2CRLo
HMRRRRRRRRRRRRH5VRBRpi=4R''MRN8pRBiP'CC2M0RC0EMR
RRRRRRRRRRRRRRMRH_osCRR<=5j"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjRj"&QR7h
2;RRRRRRRRRRRRCRM8H
V;RRRRRRRRCRM8bOsFC;##
MSC8CRoMNCs0zCR4
c;RRRRzR46RH:RVMR5F80RHsM_CRo2oCCMsCN0
RRRRRRRRRRRR_HMsRCo<5=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj&"RRh7Q2S;
CRM8oCCMsCN0R6z4;R

R7RRmRza<F=Rks0_CIo5HE80-84RF0IMF2Rj;R

RNRR8C_so=R<R7q7)R;
R-RR-CRtMNCs00CRE)CRqOvRC#DDR8NMRD#CCRO0DHFoOFRVsqR)vnA4__141R4
RzRR4:URRRHV5FOEH_OCI0H8ERR=4o2RCsMCN
0CSzRRORE	:VRHRN5R8I8sHE80R4>RcRR2oCCMsCN0
RRRRRRRRDzO	b:RsCFO#5#RB2pi
RSRRRRRLHCoMR
SRRRRRVRHRp5BiP'CCRM0NRM8BRpi=4R''02RE
CMSRRRRRRRRNRR8osC58N8s8IH04E-RI8FMR0F4Rc2<N=R8C_so85N8HsI8-0E4FR8IFM0R24c;S
SRCRRMH8RVS;
S8CMRFbsO#C#RDkO	S;
RMRC8CRoMNCs0zCRO;E	
RRRRRRRRgz4RV:RFHsRRRHM5b8C0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CRRRR-Q-RVNR58I8sHE80R4>RcM2RCRC80OFRs0CNCsRIHR0CCLMNDNCRMF8Rkk0b0MRCNCLDRD#CCRO0DHFoOR
RRRRRRzRS.:jRRRHV58N8s8IH0>ERR24cRMoCC0sNC-
S-HRVGFRVsNROD4DRd(UU,CR#D0CORRFV0#sH0CN0R0MFRHLCMsoRC#oH0CCs8R
RRRRRRRRRRRRRRkRF0M_C5RH2<'=R4I'RERCM5sN8CNo58I8sHE80-84RF0IMFcR42RR=HC2RDR#C';j'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RWRCIEMNR58C_so85N8HsI8-0E4FR8IFM0R24cRH=R2DRC#'CRj
';RRRRRRRRS8CMRMoCC0sNC.RzjR;
R-RR-VRQR85N8HsI8R0E<4=R.M2RFsRIHR0CCLMNDFCRskRF00bkRNCMLRDC#CCDOD0RFOoHRCMC8
C8RRRRRRRRRRRRzR.4:VRHR85N8HsI8R0E<4=Rco2RCsMCN
0CRRRRRRRRRRRRRRRRF_k0CHM52=R<R''4;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R R;
RRRRRRRRRCRRMo8RCsMCNR0Cz;.4
RRRRR--tCCMsCN0RC0ERv)qRDOCDN#RM08Rs#H-0CN0#R
RRRRRRzRS.:.RRsVFRH[RMIR5HE80_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNCS
SS0N0skHL0GCROs_bFRb#FAVR)_qv4UndcRX4:NRDLRCDH"#R1q)epR="&sR#P5ND[2+4R"&R,)RWQ_a v m7=&"RR_IslCF8;R
RRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqA)vn_4dXUc4RR:DCNLD#RHR1"Aa&"RR0HMCsoC'NHloIC5HE802RR&"R7"&MRH0CCosl'HN5oCHn*4d2UcR"&RW&"RR0HMCsoC'NHlo[C52RR&"R "&MRH0CCosl'HN5oCo_C0C_M880CbEH55R4+R2n*4d,UcRb8C02E2R"&RX&"RR0HMCsoC'NHlo[C5+;42
SSSLHCoMR
RRRRRRRRRRARS)_qv4UndcRX4:qR)vnA4_
14SRRRRRRRRRRRRsbF0NRlb7R5Q25jRR=>HsM_C[o52q,R7R7)=D>RFNI_858s48dRF0IMF2Rj,hR RR=> Rh,1R1)=)>R1
a,SSSSW= R>sRI0M_C5,H2RiBpRR=>B,piR57mj=2R>kRF0k_L#H45,2[2;R
RRRRRRRRRRRRRRkRF0C_so25[RR<=F_k0L4k#5[H,2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRSRRCRM8oCCMsCN0R.z.;R
RRRRRRMRC8CRoMNCs0zCR4
g;RRRRCRM8oCCMsCN0RUz4;RRRRR
RRRRR
RRRRR--tCCMsCN0RC0ERv)qRDOCDN#RM#8RCODC0FRDoRHOVRFs)Aqv41n_.z
S.:dRRRHV5FOEH_OCI0H8ERR=.o2RCsMCN
0CS-S-RGVHRsVFRDONDdR4U,U(RD#CCRO0F0VRs0H#NR0CMRF0LMCHoCRso0H#C8sC
RSRz	OERH:RVRR5Ns88I0H8ERR>4Rd2oCCMsCN0
RRRRRRRRDzO	b:RsCFO#5#RB2pi
RSRRRRRLHCoMR
SRRRRRVRHRp5BiP'CCRM0NRM8BRpi=4R''02RE
CMSRRRRRRRRNRR8osC58N8s8IH04E-RI8FMR0F4Rd2<N=R8C_so85N8HsI8-0E4FR8IFM0R24d;S
SRCRRMH8RVS;
S8CMRFbsO#C#RDkO	S;
RMRC8CRoMNCs0zCRO;E	
RRRR.SzcRR:VRFsHMRHRC58b_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
-S-RRQV58N8s8IH0>ERR24dRCMC8FR0RCOsNR0CI0sHCMRCNCLDR8NMR0FkbRk0CLMND#CRCODC0FRDo
HORRRRRRRRS6z.RH:RVNR58I8sHE80R4>Rdo2RCsMCN
0CSR--VRHGVRFsODNDRU4dUR(,#CCDOF0RVsR0HN#00MCRFL0RCoHMRosCHC#0s
C8RRRRRRRRRRRRRRRRF_k0CHM52=R<R''4RCIEMNR58osC58N8s8IH04E-RI8FMR0F4Rd2=2RHR#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=WI RERCM5_N8s5CoNs88I0H8ER-48MFI04FRd=2RRRH2CCD#R''j;R
RRRRRRCRSMo8RCsMCNR0Cz;.6
-S-RRQV58N8s8IH0<ER=dR42FRMRHIs0CCRMDNLCsRFR0FkbRk0CLMND#CRCODC0FRDoRHOM8CCCR8
SRRRR.SznRR:H5VRNs88I0H8E=R<R24dRMoCC0sNCR
SRRRRRRRRRFRRkC0_M25HRR<=';4'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RW;R
RRRRRRCRSMo8RCsMCNR0Cz;.n
-S-RMtCC0sNCER0CqR)vCRODRD#NRM80-sH#00NCR#
RRRRRSRRzR.(:FRVsRR[H5MRI0H8Ek_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0SC
S0SN0LsHkR0CGbO_s#FbRRFVAv)q_gU4.RX.:NRDLRCDH"#R1q)epR="&sR#P5ND.+*[.FR8IFM0R[.*+R42&,R"RQW)av _m=7 "RR&Ils_F;8C
RRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVAv)q_gU4.RX.:NRDLRCDH"#RA"1aRH&RMo0CCHs'lCNo58IH0RE2&7R""RR&HCM0o'CsHolNC*5HU.4g2RR&"RW"&MRH0CCosl'HN5oC[2*.R"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05R5H+2R4*gU4.8,RCEb02&2RR""XRH&RMo0CCHs'lCNo5+5[4.2*2S;
SCSLo
HMRRRRRRRRRRRRSqA)v4_Ug..XR):Rq4vAn._1
RSRRRRRRRRRRFRbsl0RN5bR7=QR>MRH_osC5[.*+84RF0IMF*R.[R2,q)77RR=>D_FINs885R4.8MFI0jFR2 ,Rh>R=R, hR)11RR=>),1a
SSSSRW =I>RsC0_M25H,pRBi>R=RiBp,mR75R42=F>RkL0_k5#.H*,.[2+4,mR75Rj2=F>RkL0_k5#.H.,R*2[2;R
RRRRRRRRRRRRRRkRF0C_so*5.[<2R=kRF0k_L#H.5,[.*2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C.o5*4[+2=R<R0Fk_#Lk.,5H.+*[4I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRS8CMRMoCC0sNC.Rz(R;
RRRRS8CMRMoCC0sNC.RzcR;
RCRRMo8RCsMCNR0Cz;.dR
R
SRRRRR--tCCMsCN0RC0ERv)qRDOCDN#RM#8RCODC0FRDoRHOVRFs)Aqv41n_cz
S.:URRRHV5FOEH_OCI0H8ERR=co2RCsMCN
0CS-S-RGVHRsVFRDONDdR4U,U(RD#CCRO0F0VRs0H#NR0CMRF0LMCHoCRso0H#C8sC
RSRz	OERH:RVNR58I8sHE80R4>R.o2RCsMCN
0CRRRRRRRRz	OD:sRbF#OC#BR5p
i2SRRRRLRRCMoH
RSRRRRRRRHV5iBp'CCPMN0RMB8Rp=iRR''42ER0CSM
RRRRRRRRR8RNs5CoNs88I0H8ER-48MFI04FR.<2R=8RN_osC58N8s8IH04E-RI8FMR0F4;.2
RSSRMRC8VRH;S
SCRM8bOsFCR##k	OD;R
SR8CMRMoCC0sNCORzE
	;RRRRSgz.RV:RFHsRRRHM5b8C0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CSR--Q5VRNs88I0H8ERR>4R.2M8CCRR0FONsC0ICRsCH0RNCMLRDCNRM8Fbk0kC0RMDNLCCR#D0CORoDFHRO
RRRRRSRRzRdj:VRHR85N8HsI8R0E>.R42CRoMNCs0SC
-V-RHVGRFOsRNRDD4UdU(#,RCODC0VRFRH0s#00NCFRM0CRLHRMosHCo#s0CCR8
RRRRRRRRRRRRRFRRkC0_M25HRR<='R4'IMECR85Ns5CoNs88I0H8ER-48MFI04FR.=2RRRH2CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R ERIC5MRNs8_CNo58I8sHE80-84RF0IMF.R42RR=HC2RDR#C';j'
RRRRRRRRMSC8CRoMNCs0zCRd
j;SR--Q5VRNs88I0H8E=R<R24.RRMFI0sHCMRCNCLDRRFsFbk0kC0RMDNLCCR#D0CORoDFHMORCCC88S
RRRRRS4zdRH:RVNR58I8sHE80RR<=4R.2oCCMsCN0
RSRRRRRRRRRRkRF0M_C5RH2<'=R4
';RRRRRRRRRRRRRRRRI_s0CHM52=R<R;W 
RRRRRRRRMSC8CRoMNCs0zCRd
4;SR--tCCMsCN0RC0ERv)qRDOCDN#RM08Rs#H-0CN0#R
RRRRRRzRSd:.RRsVFRH[RMIR5HE80_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNCS
SS0N0skHL0GCROs_bFRb#FAVR)_qvcnjgX:cRRLDNCHDR#1R")peq=&"RRP#sNcD5*c[+RI8FMR0Fc+*[4&2RRR",Wa)Q m_v7" =RI&RsF_l8
C;RRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FAVR)_qvcnjgX:cRRLDNCHDR#AR"1Ra"&MRH0CCosl'HN5oCI0H8E&2RR""7RH&RMo0CCHs'lCNo5cH*j2gnR"&RW&"RR0HMCsoC'NHlo[C5*Rc2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50E5+HRR*42cnjg,CR8b20E2RR&"RX"&MRH0CCosl'HN5oC54[+22*c;S
SSoLCHRM
RRRRRRRRRSRRAv)q_gcjnRXc:qR)vnA4_
1cSRRRRRRRRRRRRsbF0NRlb7R5Q>R=R_HMs5Coc+*[dFR8IFM0R[c*2q,R7R7)=D>RFNI_858s484RF0IMF2Rj,hR RR=> Rh,1R1)=)>R1Ra,
SSSSRW =I>RsC0_M25H,pRBi>R=RiBp,mR75Rd2=F>RkL0_k5#cHc,R*d[+27,Rm25.RR=>F_k0Lck#5cH,*.[+2
,RSSSS74m52>R=R0Fk_#Lkc,5Hc+*[4R2,7jm52>R=R0Fk_#Lkc,5HR[c*2
2;RRRRRRRRRRRRRRRRF_k0s5Coc2*[RR<=F_k0Lck#5cH,*R[2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5[c*+R42<F=RkL0_k5#cH*,c[2+4RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so*5c[2+.RR<=F_k0Lck#5cH,*.[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cco5*d[+2=R<R0Fk_#Lkc,5Hc+*[dI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRS8CMRMoCC0sNCdRz.R;
RRRRS8CMRMoCC0sNC.RzgR;
RCRRMo8RCsMCNR0Cz;.U
R
SR-RR-CRtMNCs00CRE)CRqOvRC#DDR8NMRD#CCRO0DHFoOFRVsqR)vnA4_
1gSdzdRH:RVOR5EOFHCH_I8R0E=2RgRMoCC0sNCS
S-V-RHVGRFOsRNRDD4UdU(#,RCODC0VRFRH0s#00NCFRM0CRLHRMosHCo#s0CCS8
RORzE:	RRRHV58RN8HsI8R0E>4R42CRoMNCs0RC
RRRRRzRRO:D	RFbsO#C#Rp5BiS2
RRRRRCRLo
HMSRRRRRRRH5VRB'piCMPC0MRN8pRBiRR='24'RC0EMR
SRRRRRRRRRsN8CNo58I8sHE80-84RF0IMF4R42=R<R_N8s5CoNs88I0H8ER-48MFI04FR4
2;SRSRR8CMR;HV
CSSMb8RsCFO#k#RO;D	
RSRCRM8oCCMsCN0REzO	R;
RSRRzRdc:FRVsRRHH5MR80CbEk_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0SC
-Q-RVNR58I8sHE80R4>R4M2RCRC80OFRs0CNCsRIHR0CCLMNDNCRMF8Rkk0b0MRCNCLDRD#CCRO0DHFoOR
RRRRRRzRSd:6RRRHV58N8s8IH0>ERR244RMoCC0sNC-
S-HRVGFRVsNROD4DRd(UU,CR#D0CORRFV0#sH0CN0R0MFRHLCMsoRC#oH0CCs8R
RRRRRRRRRRRRRRkRF0M_C5RH2<'=R4I'RERCM5sN8CNo58I8sHE80-84RF0IMF4R42RR=HC2RDR#C';j'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RWRCIEMNR58C_so85N8HsI8-0E4FR8IFM0R244RH=R2DRC#'CRj
';RRRRRRRRS8CMRMoCC0sNCdRz6S;
-Q-RVNR58I8sHE80RR<=4R42MIFRsCH0RNCMLRDCFFsRkk0b0MRCNCLDRD#CCRO0DHFoOCRMC88C
RRSRSRRzRdn:VRHR85N8HsI8R0E<4=R4o2RCsMCN
0CSRRRRRRRRRRRR0Fk_5CMH<2R=4R''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=W
 ;RRRRRRRRS8CMRMoCC0sNCdRznS;
-t-RCsMCNR0C0REC)RqvODCD#MRN8sR0H0-#N#0C
RRRRRRRRdSz(RR:VRFs[MRHRH5I8_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
SSSNs00H0LkCORG_FbsbF#RV)RAq.v_jXcUURR:DCNLD#RHR)"1e=qp"RR&#NsPD*5g[R+g8MFI0gFR*4[+2RR&"W,R) Qa_7vm R="&sRI_8lFCR;
RRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)RAq.v_jXcUURR:DCNLD#RHR1"Aa&"RR0HMCsoC'NHloIC5HE802RR&"R7"&MRH0CCosl'HN5oCHj*.cRU2&WR""RR&HCM0o'CsHolNC*5[g&2RR"" RH&RMo0CCHs'lCNo50oC_8CM_b8C05E5HRR+4.2*j,cURb8C02E2R"&RX&"RR0HMCsoC'NHlo5C5[2+4*;g2
SSSLHCoMR
RRRRRRRRRRARS)_qv.UjcX:URRv)qA_4n1Sg
RRRRRRRRRRRRb0FsRblNRQ57RR=>HsM_Cgo5*([+RI8FMR0Fg2*[,7Rq7=)R>FRDI8_N84s5jFR8IFM0R,j2RR h= >Rh1,R1=)R>1R)a
,RSSSSW= R>sRI0M_C5,H2RiBpRR=>B,piR57m(=2R>kRF0k_L#HU5,[U*+,(2R57mn=2R>kRF0k_L#HU5,[U*+,n2RS
SSmS75R62=F>RkL0_k5#UH*,U[2+6,mR75Rc2=F>RkL0_k5#UH*,U[2+c,mR75Rd2=F>RkL0_k5#UH*,U[2+d,SR
S7SSm25.RR=>F_k0LUk#5UH,*.[+27,Rm254RR=>F_k0LUk#5UH,*4[+27,Rm25jRR=>F_k0LUk#5UH,*,[2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75Quj=2R>MRH_osC5[g*+,U2Ru7m5Rj2=b>RN0sH$k_L#HU5,2[2;R
RRRRRRRRRRRRRRkRF0C_so*5g[<2R=kRF0k_L#HU5,[U*2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cgo5*4[+2=R<R0Fk_#LkU,5HU+*[4I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cog+*[.<2R=kRF0k_L#HU5,[U*+R.2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5[g*+Rd2<F=RkL0_k5#UH*,U[2+dRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so*5g[2+cRR<=F_k0LUk#5UH,*c[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cgo5*6[+2=R<R0Fk_#LkU,5HU+*[6I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cog+*[n<2R=kRF0k_L#HU5,[U*+Rn2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5[g*+R(2<F=RkL0_k5#UH*,U[2+(RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so*5g[2+URR<=bHNs0L$_k5#UH2,[RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRCRSMo8RCsMCNR0Cz;d(
RRRRCRSMo8RCsMCNR0Cz;dc
RRRR8CMRMoCC0sNCdRzd
;
SRRRRR--tCCMsCN0RC0ERv)qRDOCDN#RM#8RCODC0FRDoRHOVRFs)Aqv41n_4SU
zRdU:VRHRE5OFCHO_8IH0=ERR24URMoCC0sNCS
S-V-RHVGRFOsRNRDD4UdU(#,RCODC0VRFRH0s#00NCFRM0CRLHRMosHCo#s0CCS8
RORzE:	RRRHV58RN8HsI8R0E>jR4Ro2RCsMCN
0CRRRRRRRRz	OD:sRbF#OC#BR5p
i2SRRRRLRRCMoH
RSRRRRRRRHV5iBp'CCPMN0RMB8Rp=iRR''42ER0CSM
RRRRRRRRR8RNs5CoNs88I0H8ER-48MFI04FRj<2R=8RN_osC58N8s8IH04E-RI8FMR0F4;j2
RSSRMRC8VRH;S
SCRM8bOsFCR##k	OD;R
SR8CMRMoCC0sNCORzE
	;RRRRSgzdRV:RFHsRRRHM5b8C0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CSR--Q5VRNs88I0H8ERR>4Rj2M8CCRR0FONsC0ICRsCH0RNCMLRDCNRM8Fbk0kC0RMDNLCCR#D0CORoDFHRO
RRRRRSRRzRcj:VRHR85N8HsI8R0E>jR42CRoMNCs0SC
-V-RHVGRFOsRNRDD4UdU(#,RCODC0VRFRH0s#00NCFRM0CRLHRMosHCo#s0CCR8
RRRRRRRRRRRRRFRRkC0_M25HRR<='R4'IMECR85Ns5CoNs88I0H8ER-48MFI04FRj=2RRRH2CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R ERIC5MRNs8_CNo58I8sHE80-84RF0IMFjR42RR=HC2RDR#C';j'
RRRRRRRRMSC8CRoMNCs0zCRc
j;SR--Q5VRNs88I0H8E=R<R24jRRMFI0sHCMRCNCLDRRFsFbk0kC0RMDNLCCR#D0CORoDFHMORCCC88S
RRRRRS4zcRH:RVNR58I8sHE80RR<=4Rj2oCCMsCN0
RSRRRRRRRRRRkRF0M_C5RH2<'=R4
';RRRRRRRRRRRRRRRRI_s0CHM52=R<R;W 
RRRRRRRRMSC8CRoMNCs0zCRc
4;SR--tCCMsCN0RC0ERv)qRDOCDN#RM08Rs#H-0CN0#R
RRRRRRzRSc:.RRsVFRH[RMIR5HE80_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNCS
SS0N0skHL0GCROs_bFRb#FAVR)_qv4cj.XR4n:NRDLRCDH"#R1q)epR="&sR#P5ND4[U*+R4U8MFI04FRU+*[4&2RRR",Wa)Q m_v7" =RI&RsF_l8
C;RRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FAVR)_qv4cj.XR4n:NRDLRCDH"#RA"1aRH&RMo0CCHs'lCNo58IH0RE2&7R""RR&HCM0o'CsHolNC*5H4cj.2RR&"RW"&MRH0CCosl'HN5oC[U*42RR&"R "&MRH0CCosl'HN5oCo_C0C_M880CbEH55R4+R2j*4.Rc,80CbER22&XR""RR&HCM0o'CsHolNC[55+*424;U2
SSSLHCoMR
RRRRRRRRRRARS)_qv4cj.XR4n:qR)vnA4_U14
RRRRRRRRRRRRRRRRbRRFRs0lRNb5R7Q=H>RMC_soU54*4[+6FR8IFM0R*4U[R2,q)77RR=>D_FINs8858gRF0IMF2Rj,hR RR=> Rh,1R1)=)>R1Ra,
SSSSRW =I>RsC0_M25H,pRBi>R=RiBp,mR75246RR=>F_k0L4k#n,5H4[n*+246,mR7524cRR=>F_k0L4k#n,5H4[n*+24c,SR
S7SSmd542>R=R0Fk_#Lk4Hn5,*4n[d+427,Rm.542>R=R0Fk_#Lk4Hn5,*4n[.+427,Rm4542>R=R0Fk_#Lk4Hn5,*4n[4+42
,RSSSS74m5j=2R>kRF0k_L#54nHn,4*4[+jR2,7gm52>R=R0Fk_#Lk4Hn5,*4n[2+g,mR75RU2=F>RkL0_kn#454H,n+*[U
2,SSSS7(m52>R=R0Fk_#Lk4Hn5,*4n[2+(,mR75Rn2=F>RkL0_kn#454H,n+*[nR2,76m52>R=R0Fk_#Lk4Hn5,*4n[2+6,S
SSRRRR57mc=2R>kRF0k_L#54nHn,4*c[+27,Rm25dRR=>F_k0L4k#n,5H4[n*+,d2R57m.=2R>kRF0k_L#54nHn,4*.[+2S,
SRRRRRRRR57m4=2R>kRF0k_L#54nHn,4*4[+27,Rm25jRR=>F_k0L4k#n,5H4[n*2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRR7RQu=H>RMC_soU54*4[+(FR8IFM0R*4U[n+42R,
RRRRRRRRRRRRRRRRRRRRRRRRR7RRm4u52>R=RsbNH_0$L4k#n,5H.+*[4R2,75muj=2R>NRbs$H0_#Lk4Hn5,[.*2
2;RRRRRRRRRRRRRRRRF_k0s5Co4[U*2=R<R0Fk_#Lk4Hn5,*4n[I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+R42<F=RkL0_kn#454H,n+*[4I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+R.2<F=RkL0_kn#454H,n+*[.I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+Rd2<F=RkL0_kn#454H,n+*[dI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+Rc2<F=RkL0_kn#454H,n+*[cI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+R62<F=RkL0_kn#454H,n+*[6I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+Rn2<F=RkL0_kn#454H,n+*[nI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+R(2<F=RkL0_kn#454H,n+*[(I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+RU2<F=RkL0_kn#454H,n+*[UI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+Rg2<F=RkL0_kn#454H,n+*[gI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+24jRR<=F_k0L4k#n,5H4[n*+24jRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*4[+4<2R=kRF0k_L#54nHn,4*4[+4I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+24.RR<=F_k0L4k#n,5H4[n*+24.RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*4[+d<2R=kRF0k_L#54nHn,4*4[+dI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+24cRR<=F_k0L4k#n,5H4[n*+24cRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*4[+6<2R=kRF0k_L#54nHn,4*4[+6I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+24nRR<=bHNs0L$_kn#45.H,*R[2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[(+42=R<RsbNH_0$L4k#n,5H.+*[4I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRS8CMRMoCC0sNCcRz.R;
RRRRS8CMRMoCC0sNCdRzgR;
RCRRMo8RCsMCNR0Cz;dU
R
SR-RR-CRtMNCs00CRE)CRqOvRC#DDR8NMRD#CCRO0DHFoOFRVsqR)vnA4_n1d
cSzdRR:H5VROHEFOIC_HE80Rd=Rno2RCsMCN
0CS-S-RGVHRsVFRDONDdR4U,U(RD#CCRO0F0VRs0H#NR0CMRF0LMCHoCRso0H#C8sC
RSRz	OERH:RVRR5Ns88I0H8ERR>gRR2oCCMsCN0
RSRRORzDR	:bOsFCR##5iBp2S
SRCRLo
HMSRSRRRHV5iBp'CCPMN0RMB8Rp=iRR''42ER0CSM
SRRRRNRR8osC58N8s8IH04E-RI8FMR0Fg<2R=8RN_osC58N8s8IH04E-RI8FMR0Fg
2;SRSRR8CMR;HV
CSSMb8RsCFO#k#RO;D	
RSRCRM8oCCMsCN0REzO	S;
RRRRzRcc:FRVsRRHH5MR80CbEk_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0SC
-Q-RVNR58I8sHE80Rg>R2CRMC08RFsROCCN0RHIs0CCRMDNLCMRN8kRF00bkRNCMLRDC#CCDOD0RFOoH
SSSzRc6:VRHR85N8HsI8R0E>2RgRMoCC0sNC-
S-HRVGFRVsNROD4DRd(UU,CR#D0CORRFV0#sH0CN0R0MFRHLCMsoRC#oH0CCs8S
SSkSF0M_C5RH2<'=R4I'RERCM5sN8CNo58I8sHE80-84RF0IMF2RgRH=R2DRC#'CRj
';SSSSI_s0CHM52=R<RRW IMECR85N_osC58N8s8IH04E-RI8FMR0Fg=2RRRH2CCD#R''j;S
SS8CMRMoCC0sNCcRz6S;
-Q-RVNR58I8sHE80RR<=gM2RFsRIHR0CCLMNDFCRskRF00bkRNCMLRDC#CCDOD0RFOoHRCMC8
C8SzSSc:nRRRHV58N8s8IH0<ER=2RgRMoCC0sNCS
SSkSF0M_C5RH2<'=R4
';SSSSI_s0CHM52=R<R;W 
SSSCRM8oCCMsCN0Rnzc;-
S-CRtMNCs00CRE)CRqOvRC#DDR8NMRH0s-N#00
C#SzSSc:(RRsVFRH[RMIR5HE80_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNCS
SS0N0skHL0GCROs_bFRb#FAVR)_qv6X4.d:.RRLDNCHDR#1R")peq=&"RRP#sNdD5n+*[d8nRF0IMFnRd*4[+2RR&"W,R) Qa_7vm R="&sRI_8lFCR;
RRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)RAq6v_4d.X.RR:DCNLD#RHR1"Aa&"RR0HMCsoC'NHloIC5HE802RR&"R7"&MRH0CCosl'HN5oCH4*6.&2RR""WRH&RMo0CCHs'lCNo5d[*n&2RR"" RH&RMo0CCHs'lCNo50oC_8CM_b8C05E5HRR+462*4R.,80CbER22&XR""RR&HCM0o'CsHolNC[55+*42d;n2
SSSLHCoMS
SS)SAq6v_4d.X.RR:)Aqv41n_dRn
RRRRRRRRRRRRRRRRRRRRRRRRRbRRFRs0lRNb5R7Q=H>RMC_son5d*d[+4FR8IFM0R*dn[R2,q)77RD=>FNI_858sUFR8IFM0R,j2RR h= >Rh1,R1=)R>1R)aS,
SWSS >R=R0Is_5CMHR2,BRpi=B>RpRi,7dm54=2R>kRF0k_L#5d.H.,d*d[+4R2,7dm5j=2R>kRF0k_L#5d.H.,d*d[+j
2,SSSS7.m5g=2R>kRF0k_L#5d.H.,d*.[+gR2,7.m5U=2R>kRF0k_L#5d.H.,d*.[+UR2,7.m5(=2R>kRF0k_L#5d.H.,d*.[+(
2,SSSS7.m5n=2R>kRF0k_L#5d.H.,d*.[+nR2,7.m56=2R>kRF0k_L#5d.H.,d*.[+6R2,7.m5c=2R>kRF0k_L#5d.H.,d*.[+c
2,SSSS7.m5d=2R>kRF0k_L#5d.H.,d*.[+dR2,7.m5.=2R>kRF0k_L#5d.H.,d*.[+.R2,7.m54=2R>kRF0k_L#5d.H.,d*.[+4
2,SSSS7.m5j=2R>kRF0k_L#5d.H.,d*.[+jR2,74m5g=2R>kRF0k_L#5d.H.,d*4[+gR2,74m5U=2R>kRF0k_L#5d.H.,d*4[+U
2,SSSS74m5(=2R>kRF0k_L#5d.H.,d*4[+(R2,74m5n=2R>kRF0k_L#5d.H.,d*4[+nR2,74m56=2R>kRF0k_L#5d.H.,d*4[+6
2,SSSS74m5c=2R>kRF0k_L#5d.H.,d*4[+cR2,74m5d=2R>kRF0k_L#5d.H.,d*4[+dR2,74m5.=2R>kRF0k_L#5d.H.,d*4[+.R2,
SSSS57m4R42=F>RkL0_k.#d5dH,.+*[4,42R57m4Rj2=F>RkL0_k.#d5dH,.+*[4,j2R57mg=2R>kRF0k_L#5d.H.,d*g[+2
,RSSSS7Um52>R=R0Fk_#LkdH.5,*d.[2+U,mR75R(2=F>RkL0_k.#d5dH,.+*[(R2,7nm52>R=R0Fk_#LkdH.5,*d.[2+n,SR
S7SSm256RR=>F_k0Ldk#.,5Hd[.*+,62R57mc=2R>kRF0k_L#5d.H.,d*c[+27,Rm25dRR=>F_k0Ldk#.,5Hd[.*+,d2RS
SSmS75R.2=F>RkL0_k.#d5dH,.+*[.R2,74m52>R=R0Fk_#LkdH.5,*d.[2+4,mR75Rj2=F>RkL0_k.#d5dH,.2*[,RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRu7QRR=>HsM_Cdo5n+*[d86RF0IMFnRd*d[+.
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7u25dRR=>bHNs0L$_k.#d5cH,*d[+27,Rm.u52>R=RsbNH_0$Ldk#.,5Hc+*[.
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7u254RR=>bHNs0L$_k.#d5cH,*4[+27,Rmju52>R=RsbNH_0$Ldk#.,5Hc2*[2R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[<2R=kRF0k_L#5d.H.,d*R[2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[4<2R=kRF0k_L#5d.H.,d*4[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[2+.RR<=F_k0Ldk#.,5Hd[.*+R.2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[d<2R=kRF0k_L#5d.H.,d*d[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[2+cRR<=F_k0Ldk#.,5Hd[.*+Rc2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[6<2R=kRF0k_L#5d.H.,d*6[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[2+nRR<=F_k0Ldk#.,5Hd[.*+Rn2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[(<2R=kRF0k_L#5d.H.,d*([+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[2+URR<=F_k0Ldk#.,5Hd[.*+RU2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[g<2R=kRF0k_L#5d.H.,d*g[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[j+42=R<R0Fk_#LkdH.5,*d.[j+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[4+42=R<R0Fk_#LkdH.5,*d.[4+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[.+42=R<R0Fk_#LkdH.5,*d.[.+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[d+42=R<R0Fk_#LkdH.5,*d.[d+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[c+42=R<R0Fk_#LkdH.5,*d.[c+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[6+42=R<R0Fk_#LkdH.5,*d.[6+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[n+42=R<R0Fk_#LkdH.5,*d.[n+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[(+42=R<R0Fk_#LkdH.5,*d.[(+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[U+42=R<R0Fk_#LkdH.5,*d.[U+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[g+42=R<R0Fk_#LkdH.5,*d.[g+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[j+.2=R<R0Fk_#LkdH.5,*d.[j+.2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[4+.2=R<R0Fk_#LkdH.5,*d.[4+.2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[.+.2=R<R0Fk_#LkdH.5,*d.[.+.2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[d+.2=R<R0Fk_#LkdH.5,*d.[d+.2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[c+.2=R<R0Fk_#LkdH.5,*d.[c+.2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[6+.2=R<R0Fk_#LkdH.5,*d.[6+.2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[n+.2=R<R0Fk_#LkdH.5,*d.[n+.2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[(+.2=R<R0Fk_#LkdH.5,*d.[(+.2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[U+.2=R<R0Fk_#LkdH.5,*d.[U+.2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[g+.2=R<R0Fk_#LkdH.5,*d.[g+.2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[j+d2=R<R0Fk_#LkdH.5,*d.[j+d2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[4+d2=R<R0Fk_#LkdH.5,*d.[4+d2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[.+d2=R<RsbNH_0$Ldk#.,5Hc2*[RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*+2ddRR<=bHNs0L$_k.#d5cH,*4[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[c+d2=R<RsbNH_0$Ldk#.,5Hc+*[.I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*d[+6<2R=NRbs$H0_#LkdH.5,[c*+Rd2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
SSSCRM8oCCMsCN0R(zc;S
SCRM8oCCMsCN0Rczc;C
SMo8RCsMCNR0Cz;cd
M
C8sRNO0EHCkO0sMCRFI_s_COEO
	;
R--p0N#RbHlDCClM00NHRFMH8#RCkVNDN0
sHOE00COkRsC#CCDOs0_NFlRVqR)v)h_W#RH
MVkOF0HMCRo0M_C8C_8b50E#CHxRH:RMo0CC;sRRb8C0:ERR0HMCsoC2CRs0MksR0HMCsoCR
H#PHNsNCLDRMlH_x#HCRR:HCM0oRCs:j=R;C
Lo
HMRHRlMH_#x:CR=CR8b;0E
HRRV#R5HRxC<CR8b20ERC0EMR
RRHRlMH_#x:CR=HR#x
C;RMRC8VRH;R
RskC0slMRH#M_H;xC
8CMR0oC_8CM_b8C0
E;O#FM00NMRlMk_DOCD:#RR0HMCsoCRR:=5855CEb0R4-R2RR/dR.2+5R55b8C0-ERRR42lRF8dR.2/nR42R2;R-R-RFyRVqR)vXd.4O1RC#DDRCMC8RC8
MOF#M0N0CRDVF0_PRCs:MRH0CCos=R:R55580CbERR+4R62lRF8dR.2/nR42R;RRRRRRRRRRRRRRRRRRRRRR-RR-RRyF)VRqnv4XR41M8CCCV8RFDsRCRV0FsPCRsIF80#
$RbCF_k0L_k#0C$bRRH#NNss$MR5kOl_C#DDRI8FMR0FjI,RHE80-84RF0IMF2RjRRFV#_08DHFoO#;
HNoMDkRF0k_L#RR:F_k0L_k#0C$b;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFV80FkRM5HbRk000FRs#H-0CN0##2
HNoMDkRF0M_CR#:R0D8_FOoH_OPC05FsM_klODCD#FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--CLMNDRC#VRFs0-sH#00NC##
HNoMDkRF0M_C_R4n:0R#8F_Do;HO
o#HMRNDI_s0C:MRR8#0_oDFHPO_CFO0sk5MlC_ODRD#8MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-sRIHR0CCLMNDRC#VRFsCENORIsFRRFV)RqvODCD#H
#oDMNR0Is__CM4:nRR8#0_oDFH
O;#MHoNHDRMC_soRR:#_08DHFoOC_POs0F58IH04E-RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RCk#8FR0RosCHC#0sQR7h#R
HNoMDkRF0C_soRR:#_08DHFoOC_POs0F58IH04E-RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--k8#CRR0FsHCo#s0CRz7maH
#oDMNR_N8sRCo:0R#8F_Do_HOP0COFNs58I8sHE80-84RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-k-R#RC80sFRC#oH0RCsq)77
o#HMRNDD_FINs88R#:R0D8_FOoH_OPC05FscFR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-8RN8LsRHR0#HkMb0FR0Rv)qRDOCD5#RcHRL0s#RCHJks2C8
0N0skHL0\CR3lsN_VFV#\C0R#:R0MsHo
;
LHCoMR

R-RR-VRQR8N8s8IH0<ERRN6R#o#HMjR''FR0RkkM#RC8L#H0
RRRRRzjRH:RVNR58I8sHE80R4=R2CRoMNCs0RC
RRRRRDRRFNI_8R8s<"=Rjjjj"RR&Ns8_Cjo52R;
RCRRMo8RCsMCNR0Cz
j;RRRRzR4R:VRHR85N8HsI8R0E=2R.RMoCC0sNCR
RRRRRRFRDI8_N8<sR=jR"jRj"&8RN_osC584RF0IMF2Rj;R
RRMRC8CRoMNCs0zCR4R;
RzRR.:RRRRHV58N8s8IH0=ERRRd2oCCMsCN0
RRRRRRRRIDF_8N8s=R<Rj"j"RR&Ns8_C.o5RI8FMR0Fj
2;RRRRCRM8oCCMsCN0R;z.
RRRRRzdRH:RVNR58I8sHE80Rc=R2CRoMNCs0RC
RRRRRDRRFNI_8R8s<'=Rj&'RR_N8s5CodFR8IFM0R;j2
RRRR8CMRMoCC0sNCdRz;R
RRcRzRRR:H5VRNs88I0H8ERR>co2RCsMCN
0CRRRRRRRRD_FINs88RR<=Ns8_Cco5RI8FMR0Fj
2;RRRRCRM8oCCMsCN0R;zc
R
RR-R-RRQV5M8H_osC2CRso0H#C7sRQkhR#oHMRiBp
RRRRRz6RH:RV8R5HsM_CRo2oCCMsCN0
RRRRRRRRFbsO#C#Rp5Bi7,RQRh2LHCoMR
RRRRRRRRRRVRHRp5BiRR='R4'NRM8B'piCMPC002RE
CMRRRRRRRRRRRRRRRRHsM_C<oR=QR7hR;
RRRRRRRRRCRRMH8RVR;
RRRRRCRRMb8RsCFO#
#;RRRRCRM8oCCMsCN0R;z6
RRRRRznRH:RVMR5F80RHsM_CRo2oCCMsCN0
RRRRRRRRRRRR_HMsRCo<7=RQ
h;RRRRCRM8oCCMsCN0R;zn
R
RR-R-RRQV5k8F0C_sos2RC#oH0RCs7amzRHk#MmoRB
piRRRRzR(R:VRHRF58ks0_CRo2oCCMsCN0
RRRRRRRRFbsO#C#RB5mpRi,F_k0s2CoRoLCHRM
RRRRRRRRRHRRVmR5BRpi=4R''MRN8BRmpCi'P0CM2ER0CRM
RRRRRRRRRRRRR7RRmRza<F=Rks0_C
o;RRRRRRRRRRRRCRM8H
V;RRRRRRRRCRM8bOsFC;##
RRRRRRRR8CMRMoCC0sNC(Rz;R
RRURzRRR:H5VRMRF080Fk_osC2CRoMNCs0RC
RRRRRRRRR7RRmRza<F=Rks0_C
o;RRRRCRM8oCCMsCN0R;zU
R
RR-R-RRQV58N8sC_sos2RC#oH0RCsq)77RHk#MBoRpRi
RzRRg:RRRRHV58N8sC_soo2RCsMCN
0CRRRRRRRRbOsFCR##5iBp,7Rq7R)2LHCoMR
RRRRRRRRRRVRHRp5BiRR='R4'NRM8B'piCMPC002RE
CMRRRRRRRRRRRRRRRRNs8_C<oR=7Rq7N)58I8sHE80-84RF0IMF2Rj;R
RRRRRRRRRRMRC8VRH;R
RRRRRRMRC8sRbF#OC#R;
RCRRMo8RCsMCNR0Cz
g;RRRRzR4j:VRHRF5M08RN8ss_CRo2oCCMsCN0
RRRRRRRRRRRR_N8sRCo<q=R7;7)
RRRR8CMRMoCC0sNC4RzjR;
RRRRR
RRRRRR-t-RCsMCNR0C0REC)RqvODCD#MRN8CR#D0CORoDFHRO
RzRR4:4RRsVFRHHRMMR5kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CRRRR-Q-RVNR58I8sHE80R6>R2CRMC08RFsROCCN0RHIs0CCRMDNLCMRN8kRF00bkRNCMLRDC#CCDOD0RFOoH
RRRRRRRR.z4RH:RVNR58I8sHE80R6>R2CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_M25HRR<='R4'IMECR85N_osC58N8s8IH04E-RI8FMR0F6=2RRRH2CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R ERIC5MRNs8_CNo58I8sHE80-84RF0IMF2R6RH=R2DRC#'CRj
';RRRRRRRRRRRRCRM8oCCMsCN0R.z4;R
RR-R-RRQV58N8s8IH0<ER=2R6RRMFI0sHCMRCNCLDRRFsFbk0kC0RMDNLCCR#D0CORoDFHMORCCC88R
RRRRRR4RzdRR:H5VRNs88I0H8E=R<RR62oCCMsCN0
RRRRRRRRRRRRRRRR0Fk_5CMH<2R=4R''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=W
 ;RRRRRRRRRRRRCRM8oCCMsCN0Rdz4;R
RR-R-RMtCC0sNCER0CqR)vCRODRD#NRM80-sH#00NCR#
RRRRRzRR4:cRRsVFRH[RMIR5HE80R4-R2FR8IFM0RojRCsMCN
0CRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FzVR)dqv.RR:DCNLD#RHR1"1a&"RR0HMCsoC'NHloIC5HE802RR&"R7"&MRH0CCosl'HN5oCH.*d2RR&"RW"&MRH0CCosl'HN5oC[&2RR"" RH&RMo0CCHs'lCNo50oC_8CM_b8C05E5HRR+4d2*.8,RCEb02&2RR""XRH&RMo0CCHs'lCNo54[+2R;
RRRRRRRRRLRRCMoH
RRRRRRRRRRRRqz)vRd.:qR)vXd.4
1RRRRRRRRRRRRRRRRRb0FsRblNRR57=H>RMC_so25[,jRqRR=>D_FINs885,j2RRq4=D>RFNI_858s4R2,q=.R>FRDI8_N8.s52R,
RRRRRRRRRRRRRRRRRRRRRRRRRRqd=D>RFNI_858sdR2,q=cR>FRDI8_N8cs52W,R >R=R0Is_5CMHR2,WiBpRR=>B,piR=mR>kRF0k_L#,5H[;22
RRRRRRRRRRRRRRRR0Fk_osC5R[2<F=RkL0_kH#5,R[2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRR8CMRMoCC0sNC4RzcR;
RRRRRCRRMo8RCsMCNR0Cz;44RRRRRRRRRRRR
RRRR
RRRRRR-t-RCsMCNR0CNnR4RsIF8CR8C)bRqOvRCRDDHNVRbFbsbNsH0RCRRRRRRRRRRRRRRR
RR4Rz6RR:H5VRD0CV_CFPsRR=4o2RCsMCN
0CRRRR-Q-RVNR58I8sHE80R6>R2CRMC08RFsROCCN0RHIs0CCRMDNLCMRN8kRF00bkRNCMLRDC#CCDOD0RFOoH
RRRRRRRRnz4RH:RVNR58I8sHE80R6>R2CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_Mn_4RR<='R4'IMECRN558C_so85N8HsI8-0E4FR8IFM0RR62=kRMlC_OD2D#R8NMR85N_osC5Rc2=jR''R22CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C_R4n<W=R ERIC5MR5_N8s5CoNs88I0H8ER-48MFI06FR2RR=M_klODCD#N2RM58RNs8_Cco52RR='2j'2DRC#'CRj
';RRRRRRRRRRRRCRM8oCCMsCN0Rnz4;R
RR-R-RRQV58N8s8IH0<ER=2R6RRMFI0sHCMRCNCLDRRFsFbk0kC0RMDNLCCR#D0CORoDFHMORCCC88R
RRRRRR4Rz(RR:H5VRNs88I0H8E=R<RR62oCCMsCN0
RRRRRRRRRRRRRRRR0Fk__CM4<nR=4R''R;
RRRRRRRRRRRRRIRRsC0_Mn_4RR<=W
 ;RRRRRRRRRRRRCRM8oCCMsCN0R(z4;R
RR-R-RMtCC0sNCER0CqR)vCRODNDRM08Rs#H-0CN0
RRRRRRRRUz4RV:RF[sRRRHM58IH0-ERRR428MFI0jFRRMoCC0sNCR
RRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqz)vR4n:NRDLRCDH"#R1"1aRH&RMo0CCHs'lCNo58IH0RE2&7R""RR&HCM0o'CsHolNCk5MlC_OD*D#dR.2&WR""RR&HCM0o'CsHolNC25[R"&R &"RR0HMCsoC'NHlo8C5CEb02RR&"RX"&MRH0CCosl'HN5oC[2+4;R
RRRRRRRRRRCRLo
HMRRRRRRRRRRRRzv)q4:nRRv)q44nX1RR
RRRRRRRRRRRRRbRRFRs0lRNb5=7R>MRH_osC5,[2RRqj=D>RFNI_858sjR2,q=4R>FRDI8_N84s52q,R.>R=RIDF_8N8s25.,R
RRRRRRRRRRRRRRRRRRRRRRRRRq=dR>FRDI8_N8ds52W,R >R=R0Is__CM4Rn,WiBpRR=>B,piR=mR>kRF0k_L#k5MlC_OD,D#[;22
RRRRRRRRRRRRRRRR0Fk_osC5R[2<F=RkL0_kM#5kOl_C#DD,R[2IMECRk5F0M_C_R4n=4R''C2RDR#C';Z'
RRRRRRRRRRRR8CMRMoCC0sNC4RzUR;
RRRRRCRRMo8RCsMCNR0Cz;46RRRRRRRRR
R
CRM8NEsOHO0C0CksRD#CC_O0s;Nl
