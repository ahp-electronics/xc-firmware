--
@ER--B$FbsEHo0OR52gR4g-cRRj.jd$R1MHbDO$H0ROQM
R--fN]C8:CsR#//$DMbH0OH$N/lb0DN.Uj4J4.b/blNb#Cs/0N0/LDH/MoC_OFsN/dOs_NlsPI3E48yR-f
-


---
-HR1lCbDRv)qR0IHEHR#MCoDR7q7)1 1RsVFRNsC8MRN8sRIH
0C-a-RNCso0RR:pCkOM-0RRBm)qBRd

--DsHLNRs$HCCC;#
kCCRHC#C30D8_FOoH_n44cD3NDk;
#HCRC3CC#_08DHFoOH_#o8MC3DND;#
kCCRHC#C30D8_FOoH_HNs0NE3D
D;DsHLNRs$FNsOdk;
#FCRsdON3OFsNlOFbD3NDC;
M00H$qR)vW_)R
H#RRRRoCCMsRHO5R
RRRRRRNRVl$HD:0R#soHMRR:="MMFC
";RRRRRRRRI0H8ERR:HCM0oRCs:(=R;RR
RRRRRNRR8I8sHE80RH:RMo0CC:sR=;R(RRRRRRRR-L-RHCoRMoFkEFRVsCR8b
0ERRRRRRRR80CbERR:HCM0oRCs:R=R4;.U
RRRRRRRRk8F0C_soRR:LDFFCRNM:V=RNCD#;RRRR-R-R#ENR0FkbRk0s
CoRRRRRRRR8_HMsRCo:FRLFNDCM=R:RDVN#RC;RRRRRR--ERN#8NN0RbHMks0RCRo
RRRRRNRR8_8ssRCo:FRLFNDCM=R:RDVN#RCRRRRR-E-RNs8RCRN8Ns88CR##s
CoRRRRRRRR2R;
RbRRFRs05R
RRRRRRmR7zRaR:kRF00R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj;R
RRRRRRQR7hRRR:MRHR0R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj;R
RRRRRR7Rq7R)R:MRHR0R#8F_Do_HOP0COFNs58I8sHE80-84RF0IMF2Rj;R
RRRRRR RWRRRR:MRHR0R#8F_Do;HORRRRR-RR-sRIHR0CCLMNDVCRFssRNRl
RRRRRBRRpRiRRH:RM#RR0D8_FOoH;RRRRRRR-O-RD	FORsVFRlsN,8RN8Rs,8
HMRRRRRRRRmiBpRRR:HRMR#_08DHFoORRRRRRRRR--FRb0OODF	FRVsFR8kR0
RRRRR2RR;M
C8MRC0$H0Rv)q_;)W
-
-
R--w#Hs0lRHblDCCNM00MHFR#lk0CRLRDONDRC8NEsOj-
-
ONsECH0Os0kCsRNOREjF)VRq)v_W#RH
MOF#M0N0kRMlC_OD_D#8bCCRH:RMo0CC:sR=5R580CbERR-4d2/.R2;RRRRRRRR-y-RRRFVs#FIRRFV)dB .RXcODCD#CRMC88C
MOF#M0N0kRMlC_OD_D#ICH8RH:RMo0CC:sR=5R5I0H8ERR-4c2/2R;RRRRRRRRR-y-RRRFVOkFDlRM#F)VRB. dXOcRC#DDRCMC8
C80C$bR0Fk_#Lk_b0$C#RHRsNsN5$RM_klODCD#C_8C8bRF0IMF,RjRk5MlC_OD_D#ICH8*+c2dFR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNR0Fk_#LkR:RRR0Fk_#Lk_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFV80FkRM5HbRk000FRs#H-0CN0##2
HNoMDkRF0M_CRRRR:0R#8F_Do_HOP0COFMs5kOl_C#DD_C8CbFR8IFM0R;j2R-R-RNCML#DCRsVFRH0s-N#00
C##MHoNIDRb_CjCRMRR#:R0D8_FOoH_OPC05FsM_klODCD#C_8C8bRF0IMF2Rj;-RR-sRIHR0CCLMNDRC#VRFsCENORIsFRRFV)RqvODCD#H
#oDMNRCIb4M_CR:RRR8#0_oDFHPO_CFO0sk5MlC_OD_D#8bCCRI8FMR0FjR2;RR--I0sHCMRCNCLD#FRVsNRCOsERFFIRVqR)vCROD
D##MHoNHDRMC_soRRRR#:R0D8_FOoH_OPC05FsI0H8ER+d8MFI0jFR2R;RRRRRR-RR-#RkC08RFCRso0H#C7sRQ
hR#MHoNFDRks0_CRoRR#:R0D8_FOoH_OPC05FsI0H8ER+d8MFI0jFR2R;RRRRRR-RR-#RkC08RFCRso0H#C7sRm
za#MHoNWDR  _)tR4RR#:R0D8_FOoH;H
#oDMNR_HMs4CoR:RRR8#0_oDFHPO_CFO0sH5I8+0EdFR8IFM0R;j2RRRR
o#HMRNDNs8_CRoRRRR:#_08DHFoOC_POs0F58N8s8IH04E-RI8FMR0FjR2;RRRR-k-R#RC80sFRC#oH0RCsq)77
o#HMRNDD_FINs88RRR:#_08DHFoOC_POs0F58cRF0IMF2Rj;RRRRRRRRRRRRRRR-N-R8R8sL#H0RbHMk00RFqR)vCRODRD#5L6RHR0#skCJH8sC2$
0b0CRlNb_8_8s0C$bRRH#NNss$MR5kOl_C#DD_C8CbFR8IFM0RRj2F#VR0D8_FOoH_OPC0RFs58gRF0IMF2Rj;H
#oDMNRb0l_8N8s:RRRb0l_8N8s$_0b
C;
oLCH
M
RRRR-Q-RV8RN8HsI8R0E<RR6NH##o'MRj0'RFMRkk8#CR0LH#R
RR4RzRRR:H5VRNs88I0H8ERR=4o2RCsMCN
0CRRRRRRRRD_FINs88RR<="jjjj&"RR_N8s5Coj
2;RRRRCRM8oCCMsCN0R;z4
RRRRRz.RH:RVNR58I8sHE80R.=R2CRoMNCs0RC
RRRRRDRRFNI_8R8s<"=Rj"jjRN&R8C_soR548MFI0jFR2R;
RCRRMo8RCsMCNR0Cz
.;RRRRzRdR:VRHR85N8HsI8R0E=2RdRMoCC0sNCR
RRRRRRFRDI8_N8<sR=jR"j&"RR_N8s5Co.FR8IFM0R;j2
RRRR8CMRMoCC0sNCdRz;R
RRcRzRRR:H5VRNs88I0H8ERR=co2RCsMCN
0CRRRRRRRRD_FINs88RR<='Rj'&8RN_osC58dRF0IMF2Rj;R
RRMRC8CRoMNCs0zCRcR;
RzRR6:RRRRHV58N8s8IH0>ERRRc2oCCMsCN0
RRRRRRRRIDF_8N8s=R<R_N8s5CocFR8IFM0R;j2
RRRR8CMRMoCC0sNC6Rz;R

R-RR-VRQRH58MC_sos2RC#oH0RCs7RQhkM#HopRBiR
RRnRzRRR:H5VR8_HMs2CoRMoCC0sNCR
RRRRRRsRbF#OC#BR5pRi,72QhRoLCHRM
RRRRRRRRRHRRVBR5p=iRR''4R8NMRiBp'CCPMR020MEC
RRRRRRRRRRRRRRRR_HMsRCo<5=R"jjjj&"RRh7Q2R;
RRRRRRRRRCRRMH8RVR;
RRRRRCRRMb8RsCFO#
#;RRRRCRM8oCCMsCN0R;zn
RRRRRz(RH:RVMR5F80RHsM_CRo2oCCMsCN0
RRRRRRRRRRRR_HMsRCo<5=R"jjjj&"RRh7Q2R;
RCRRMo8RCsMCNR0Cz
(;
RRRRFbsO#C#Rp5BiW,R H,RMC_soL2RCMoH
RRRRRRRRRHV5iBpR'=R4N'RMB8RpCi'P0CM2ER0CRM
RRRRRRRRRWRR  _)t<4R= RW;R
RRRRRRRRRRMRH_osC4=R<R_HMs;Co
RRRRRRRR8CMR;HV
RRRR8CMRFbsO#C#;R

R-RR-VRQR85N8ss_CRo2sHCo#s0CR7q7)#RkHRMoB
piRRRRzR4.RH:RVNR58_8ss2CoRMoCC0sNCR
RRRRRRsRbF#OC#BR5pRi,q)772CRLo
HMRRRRRRRRRRRRH5VRBRpi=4R''MRN8pRBiP'CC2M0RC0EMR
RRRRRRRRRRRRRR8RN_osCRR<=q)7758N8s8IH04E-RI8FMR0Fj
2;RRRRRRRRRRRRCRM8H
V;RRRRRRRRCRM8bOsFC;##
RRRR8CMRMoCC0sNC4Rz.
;
RRRRzR4d:VRHRF5M08RN8ss_CRo2oCCMsCN0
RRRRRRRRRRRR_N8sRCo<q=R757)Ns88I0H8ER-48MFI0jFR2R;
RCRRMo8RCsMCNR0Cz;4d
R
RR.Rzn:RRRRHV5k8F0C_soo2RCsMCN
0CRRRRRRRRbOsFCR##5pmBiF,Rks0_CRo2LHCoMR
RRRRRRRRRRVRHRB5mp=iRR''4R8NMRpmBiP'CC2M0RC0EMR
RRRRRRRRRRRRRRmR7z<aR=kRF0C_soH5I8-0E4FR8IFM0R;j2
RRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMRFbsO#C#;R
RRMRC8CRoMNCs0zCR.
n;
RRRRR--tCCMsCN0RC0ERD#CCRO0DHFoOR
RR4RzcRR:VRFsHMRHRlMk_DOCD8#_CRCb8MFI0jFRRMoCC0sNCR
RR-R-RHAkDF8Rkk0b0MRCNCLDRD#CCRO0DHFoOR
RRRRRR-R-RRQV58N8s8IH0>ERR246RM8F'k0R#1CRpRQBODCD#R
RRRRRR Rm4:nRRRHV58N8s8IH0>ERR246RMoCC0sNCR
RRRRRRRRRRRRRRkRF0M_C5RH2<'=R4I'RERCM5_N8s5CoNs88I0H8ER-48MFI06FR2RR=HC2RDR#C';j'
RRRRRRRR8CMRMoCC0sNC Rm4
n;RRRRRRRR-Q-RVNR58I8sHE80R6>R2hRq7NR58I8sHE80RR<=4R62kR#C1BpQRDOCDR#
RRRRRmRR R46:VRHR85N8HsI8R0E=6R42CRoMNCs0RC
RRRRRRRRRRRRR0RRlNb_858sHg25RI8FMR0Fj<2R=mRhaF5OM#P_0D8_FOoH_OPC05FsH4,RjR22XRm)Ns8_CNo58I8sHE80-84RF0IMF2R6;R
RRRRRRRRRRRRRRqR1h47_6RR:17qh4bjRFRs0lRNb5=qR>lR0b8_N8Hs5225j,RRA=0>RlNb_858sH4252B,RRR=>0_lbNs8855H2.R2,7>R=Rb0l_8N8s25H5,d2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR >R=Rb0l_8N8s25H5,c2R=wR>lR0b8_N8Hs52256,RRt=0>RlNb_858sHn252],RRR=>0_lbNs8855H2(R2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRQ>R=Rb0l_8N8s25H5,U2R=KR>lR0b8_N8Hs5225g,RRZ=F>RkC0_M25H2R;
RRRRRCRRMo8RCsMCNR0Cm6 4;R
RRRRRR Rm4:cRRRHV58N8s8IH0=ERR24cRMoCC0sNCR
RRRRRRRRRRRRRRlR0b8_N8Hs52R5U8MFI0jFR2=R<Rahm5MOFP0_#8F_Do_HOP0COFHs5,2Rg2mRX)8RN_osC58N8s8IH04E-RI8FMR0F6
2;RRRRRRRRRRRRRRRR17qh_R4c:qR1hj74RsbF0NRlbqR5RR=>0_lbNs8855H2jR2,A>R=Rb0l_8N8s25H5,42R=BR>lR0b8_N8Hs5225.,RR7=0>RlNb_858sHd252R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR =0>RlNb_858sHc252w,RRR=>0_lbNs8855H26R2,t>R=Rb0l_8N8s25H5,n2R=]R>lR0b8_N8Hs5225(,RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRQ=0>RlNb_858sHU252K,RRR=>',4'R=ZR>kRF0M_C52H2;R
RRRRRRMRC8CRoMNCs0mCR ;4c
RRRRRRRR4m dRR:H5VRNs88I0H8ERR=4Rd2oCCMsCN0
RRRRRRRRRRRRRRRRb0l_8N8s25H58(RF0IMF2RjRR<=h5maOPFM_8#0_oDFHPO_CFO0s,5HR2U2R)XmR_N8s5CoNs88I0H8ER-48MFI06FR2R;
RRRRRRRRRRRRR1RRq_h74:dRRh1q7RURb0FsRblNRR5q=0>RlNb_858sHj252A,RRR=>0_lbNs8855H24R2,B>R=Rb0l_8N8s25H5,.2R=7R>lR0b8_N8Hs5225d,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR= R>lR0b8_N8Hs5225c,RRw=0>RlNb_858sH6252t,RRR=>0_lbNs8855H2nR2,]>R=Rb0l_8N8s25H5,(2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR=ZR>kRF0M_C52H2;R
RRRRRRMRC8CRoMNCs0mCR ;4d
RRRRRRRR4m .RR:H5VRNs88I0H8ERR=4R.2oCCMsCN0
RRRRRRRRRRRRRRRRb0l_8N8s25H58nRF0IMF2RjRR<=h5maOPFM_8#0_oDFHPO_CFO0s,5HR2(2R)XmR_N8s5CoNs88I0H8ER-48MFI06FR2R;
RRRRRRRRRRRRR1RRq_h74:.RRh1q7RURb0FsRblNRR5q=0>RlNb_858sHj252A,RRR=>0_lbNs8855H24R2,B>R=Rb0l_8N8s25H5,.2R=7R>lR0b8_N8Hs5225d,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR= R>lR0b8_N8Hs5225c,RRw=0>RlNb_858sH6252t,RRR=>0_lbNs8855H2nR2,]>R=R''4,RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRZ=F>RkC0_M25H2R;
RRRRRCRRMo8RCsMCNR0Cm. 4;R
RRRRRR Rm4:4RRRHV58N8s8IH0=ERR244RMoCC0sNCR
RRRRRRRRRRRRRRlR0b8_N8Hs52R568MFI0jFR2=R<Rahm5MOFP0_#8F_Do_HOP0COFHs5,2Rn2mRX)8RN_osC58N8s8IH04E-RI8FMR0F6
2;RRRRRRRRRRRRRRRR17qh_R44:qR1hR7nRsbF0NRlbqR5RR=>0_lbNs8855H2jR2,A>R=Rb0l_8N8s25H5,42R=BR>lR0b8_N8Hs5225.,RR7=0>RlNb_858sHd252R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR =0>RlNb_858sHc252w,RRR=>0_lbNs8855H26R2,Z>R=R0Fk_5CMH;22
RRRRRRRR8CMRMoCC0sNC Rm4
4;RRRRRRRRmj 4RH:RVNR58I8sHE80R4=Rjo2RCsMCN
0CRRRRRRRRRRRRRRRR0_lbNs8855H2cFR8IFM0RRj2<h=RmOa5F_MP#_08DHFoOC_POs0F5RH,6R22XRm)Ns8_CNo58I8sHE80-84RF0IMF2R6;R
RRRRRRRRRRRRRRqR1h47_jRR:17qhnbRRFRs0lRNb5=qR>lR0b8_N8Hs5225j,RRA=0>RlNb_858sH4252B,RRR=>0_lbNs8855H2.R2,7>R=Rb0l_8N8s25H5,d2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR >R=Rb0l_8N8s25H5,c2R=wR>4R''Z,RRR=>F_k0CHM52
2;RRRRRRRRCRM8oCCMsCN0R4m jR;
RRRRRmRR RgR:VRHR85N8HsI8R0E=2RgRMoCC0sNCR
RRRRRRRRRRRRRRlR0b8_N8Hs52R5d8MFI0jFR2=R<Rahm5MOFP0_#8F_Do_HOP0COFHs5,2Rc2mRX)8RN_osC58N8s8IH04E-RI8FMR0F6
2;RRRRRRRRRRRRRRRR17qh_:gRRh1q7RcRRsbF0NRlbqR5RR=>0_lbNs8855H2jR2,A>R=Rb0l_8N8s25H5,42R=BR>lR0b8_N8Hs5225.,RR7=0>RlNb_858sHd252R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRZ=F>RkC0_M25H2R;
RRRRRCRRMo8RCsMCNR0Cm; g
RRRRRRRRUm RRR:H5VRNs88I0H8ERR=Uo2RCsMCN
0CRRRRRRRRRRRRRRRR0_lbNs8855H2.FR8IFM0RRj2<h=RmOa5F_MP#_08DHFoOC_POs0F5RH,dR22XRm)Ns8_CNo58I8sHE80-84RF0IMF2R6;R
RRRRRRRRRRRRRRqR1hU7_R1:Rqch7RbRRFRs0lRNb5=qR>lR0b8_N8Hs5225j,RRA=0>RlNb_858sH4252B,RRR=>0_lbNs8855H2.R2,7>R=R''4,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR=ZR>kRF0M_C52H2;R
RRRRRRMRC8CRoMNCs0mCR 
U;RRRRRRRRmR (RH:RVNR58I8sHE80R(=R2CRoMNCs0RC
RRRRRRRRRRRRR0RRlNb_858sH425RI8FMR0Fj<2R=mRhaF5OM#P_0D8_FOoH_OPC05FsH.,R2X2RmN)R8C_so85N8HsI8-0E4FR8IFM0R;62
RRRRRRRRRRRRRRRRh1q7R_(:qR1hR7.RFRbsl0RN5bRq>R=Rb0l_8N8s25H5,j2R=AR>lR0b8_N8Hs52254,RRZ=F>RkC0_M25H2R;
RRRRRCRRMo8RCsMCNR0Cm; (
RRRRRRRRnm RRR:H5VRNs88I0H8ERR=no2RCsMCN
0CRRRRRRRRRRRRRRRRF_k0CHM52=R<R''4RCIEMNR58C_so256RO=RF_MP#_08DHFoOC_POs0F54H,225j2DRC#'CRj
';RRRRRRRRCRM8oCCMsCN0Rnm ;R
RR-R-RRQV58N8s8IH0<ER=2R6RRMFFbk0kC0RMDNLCCR#D0CORoDFHMORCCC88RR/lRNb8CHsO$0DRR0F)'qv#8RN8#sC#HRDM
C#RRRRRRRRmR 6:VRHR85N8HsI8R0E<6=R2CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_M25HRR<=';4'
RRRRRRRR8CMRMoCC0sNC Rm6
;
RRRR-Q-RVNR58I8sHE80Rg>R2#RkCuRW 0jRFCR8OCF8R8N8s#C#R0LH#RRn0FEskRoEgMRN8uRW 04RFCR8OCF8R0LH#jR4RR+
RRRRRWRR R4j:VRHR85N8HsI8R0E>2RgRMoCC0sNCR
RRRRRRRRRRRRRRbRICCj_M25HRR<='R4'IMECR85N_osC58URF0IMF2R6RO=RF_MP#_08DHFoOC_POs0F5.H,jd25RI8FMR0FjR22CCD#R''j;R
RRRRRRRRRRRRRRbRICC4_M25HRR<='R4'IMECR85N_osC58N8s8IH04E-RI8FMR0Fg=2RRMOFP0_#8F_Do_HOP0COFHs5,2.j58N8s8IH0nE-RI8FMR0FcR22CCD#R''j;R
RRRRRRRRRRMRC8CRoMNCs0WCR ;4j
RRRRR--Q5VRNs88I0H8ERR=UsRFRRg2kR#CWju RR0F8FCO8NCR8C8s#L#RHR0#nER0soFkE
RgRRRRRRRRWR gRH:RV5R5Ns88I0H8ERR=Um2R)NR58I8sHE80Rg=R2o2RCsMCN
0CRRRRRRRRRRRRRRRRIjbC_5CMH<2R=4R''ERIC5MRNs8_CNo58I8sHE80-84RF0IMF2R6RH=R2DRC#'CRj
';RRRRRRRRRRRRRRRRI4bC_5CMH<2R=4R''R;
RRRRRRRRRCRRMo8RCsMCNR0CW; g
RRRRR--Q5VRNs88I0H8ERR=(k2R#WCRuR j08FRC8OFCER0C0RnE8RN8#sC#HRL0RR&W4u RR0F8FCO80CRE(CR0NER8C8s#L#RHR0
RRRRRWRR R(R:VRHR85N8HsI8R0E=2R(RMoCC0sNCR
RRRRRRRRRRRRRRbRICCj_M25HRR<='R4'IMECR85N_osC5R62=FROM#P_0D8_FOoH_OPC05FsH2,.52j2R#CDCjR''R;
RRRRRRRRRRRRRIRRb_C4CHM52=R<R''4RCIEMNR58C_so25nRO=RF_MP#_08DHFoOC_POs0F5.H,22542DRC#'CRj
';RRRRRRRRCRM8oCCMsCN0R(W ;R
RR-R-RRQV58N8s8IH0=ERRRn2kR#CWju RR0F8FCO80CREnCR0NER8C8s#L#RHR0
RRRRRWRR RnR:VRHR85N8HsI8R0E=2RnRMoCC0sNCR
RRRRRRRRRRRRRRbRICCj_M25HRR<='R4'IMECR85N_osC5R62=FROM#P_0D8_FOoH_OPC05FsH2,452j2R#CDCjR''R;
RRRRRRRRRRRRRIRRb_C4CHM52=R<R''4;R
RRRRRRMRC8CRoMNCs0WCR 
n;RRRR-Q-RVNR58I8sHE80RR<=6M2RFsRIHR0CCLMND#CRCODC0FRDoRHOM8CCCR8
RRRRRWRR R6R:VRHR85N8HsI8R0E<6=R2CRoMNCs0RC
RRRRRRRRRRRRRIRRb_CjCHM52=R<R''4;R
RRRRRRRRRRRRRRbRICC4_M25HRR<=';4'
RRRRRRRR8CMRMoCC0sNC RW6
;
RRRRCRM8oCCMsCN0Rcz4;R

RzRR.:6RRRHV50MFRk8F0C_soo2RCsMCN
0CRRRRRRRRz44(:sRbF#OC#WR5  _)tR4,HsM_C,o4R0Fk_osC2R
RRRRRRCRLo
HMRRRRRRRRRRRRH5VRW) _ Rt4=4R''02RE
CMRRRRRRRRRRRRRRRR7amzRR<=HsM_C5o4I0H8ER-48MFI0jFR2R;
RRRRRRRRRCRRD
#CRRRRRRRRRRRRRRRR7amzRR<=F_k0s5CoI0H8ER-48MFI0jFR2R;
RRRRRRRRRCRRMH8RVR;
RRRRRCRRMb8RsCFO#z#R4;(4
RRRR8CMRMoCC0sNC.Rz6
;
RRRR-t-RCsMCNR0C0REC)RqvODCD#HRI00ERs#H-0CN0#R
RR4Rz6RR:VRFsHMRHRlMk_DOCD8#_CRCb8MFI0jFRRMoCC0sNCR
RRRRRR4Rz(RR:VRFs[MRHRlMk_DOCDI#_HR8C8MFI0jFRRMoCC0sNCR
RRRRRRRRRR)RzqRv:)dB .RXc
RRRRRRRRRRRRRRRRsbF0NRlb7R5Q=jR>MRH_osC5*5[c,22R47QRR=>HsM_C5o5[2*c+,42R.7QRR=>HsM_C5o5[2*c+,.2Rd7QRR=>HsM_C5o5[2*c+,d2
RRRRRRRRRRRRRRRRRRRRRRRRqRR7=jR>FRDI8_N8js52q,R7=4R>FRDI8_N84s52q,R7=.R>FRDI8_N8.s52q,R7=dR>FRDI8_N8ds52q,R7=cR>FRDI8_N8cs52-,
-RRRRRRRRRRRRRRRRRRRRRRRRWRR)R h=W>R W,RuR j=I>Rb_CjCHM52W,RuR 4=I>Rb_C4CHM52B,Ri>R=RahmRiBp,RR
RRRRRRRRRRRRRRRRRRRRRRRRR W)h>R=R,W R Wuj>R=RCIbjM_C5,H2R Wu4>R=RCIb4M_C5,H2RRBi=B>RpRi,tR1)='>R4R',
RRRRRRRRRRRRRRRRRRRRRRRR7RRm=jR>kRF0k_L#,5H5c[*2R2,7Rm4=F>RkL0_kH#5,*5[c42+27,Rm=.R>kRF0k_L#,5H5c[*22+.,mR7d>R=R0Fk_#Lk55H,[2*c+2d2;R
RRRRRRRRRRRRRRkRF0C_so[55*2c2RR<=F_k0L5k#H[,5*2c2RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so[55*+c24<2R=kRF0k_L#,5H5c[*22+4RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so[55*+c2.<2R=kRF0k_L#,5H5c[*22+.RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so[55*+c2d<2R=kRF0k_L#,5H5c[*22+dRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRMRC8CRoMNCs0zCR4
(;RRRRRRRRCRM8oCCMsCN0R6z4;-

-zRR.:URRRHV5k8F0C_soo2RCsMCN
0C-R-RRRRRR4RznRR:VRFsHMRHRlMk_DOCD8#_CRCb8MFI0jFRRMoCC0sNC-
-RRRRRRRRzR4U:FRVsRR[HMMRkOl_C#DD_8IHCFR8IFM0RojRCsMCN
0C-R-RRRRRRRRRR)RzqRv:)dB .RXc
R--RRRRRRRRRRRRRbRRFRs0lRNb5j7QRR=>HsM_C5o5[2*c27,RQ=4R>MRH_osC5*5[c42+27,RQ=.R>MRH_osC5*5[c.2+27,RQ=dR>MRH_osC5*5[cd2+2-,
-RRRRRRRRRRRRRRRRRRRRRRRRqRR7=jR>FRDI8_N8js52q,R7=4R>FRDI8_N84s52q,R7=.R>FRDI8_N8.s52q,R7=dR>FRDI8_N8ds52q,R7=cR>FRDI8_N8cs52-,
-RRRRRRRRRRRRRRRRRRRRRRRRWRR)R h=W>R W,RuR j=I>Rb_CjCHM52W,RuR 4=I>Rb_C4CHM52B,Ri>R=RahmRiBp,-R
-RRRRRRRRRRRRRRRRRRRRRRRRTRR7Rmj=F>RkL0_kH#5,*5[c,22RmT74>R=R0Fk_#Lk55H,[2*c+,42RmT7.>R=R0Fk_#Lk55H,[2*c+,.2RmT7d>R=R0Fk_#Lk55H,[2*c+2d2;-
-RRRRRRRRRRRRRRRRF_k0s5Co5c[*2<2R=kRF0k_L#,5H5c[*2I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';-R-RRRRRRRRRRRRRRkRF0C_so[55*+c24<2R=kRF0k_L#,5H5c[*22+4RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;-
-RRRRRRRRRRRRRRRRF_k0s5Co5c[*22+.RR<=F_k0L5k#H[,5*+c2.I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';-R-RRRRRRRRRRRRRRkRF0C_so[55*+c2d<2R=kRF0k_L#,5H5c[*22+dRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;-
-RRRRRRRRRRRRCRM8oCCMsCN0RUz4;-
-RRRRRCRRMo8RCsMCNR0Cz;4n
R--RCRRMo8RCsMCNR0Cz;.U
-
-RRRRRURkRH:RV8R5F_k0s2CoRMoCC0sNC-
-RRRRRRRRRmR7z<aR=kRF0C_soH5I8-0E4FR8IFM0R;j2
R--R8CMRMoCC0sNCURk;R
RRRRRRRRRRRRRR
RRCRM8NEsOHO0C0CksRONsE
j;
