--$Header: //synplicity/maplat2018q2p1/designware/dw03.vhd#1 $
@E---------------------------------------------------------------------------------------------------

---w-RHRDCRRRRR:RRRj8IdE3P8-
-R#7CHRoMRRRRRB:RFNM0HRM#4LURNO#HR#7CHWoMNRsCObFlFMMC0
#R-B-RFNlbMR$RR:RRRM1$bODHHR0$Q3MO
R--7CN0RRRRRRRR:kRqo6R.,jR.j-U
-kRq0sEFRRRRRRR:1PCDN)lR
R--e#CsHRFMRRRR:3Rd4-
-
---------------------------------------------------------------------------------------------------
H
DLssN$CRHC
C;kR#CHCCC38#0_oDFH4O_43ncN;DD
Ck#RCHCC03#8F_Do_HOkHM#o8MC3DND;


CHM007$RW_jdbCHb_osCR
H#RRRRoCCMs5HORRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR
RRRRRRRRRIRRHE80RQ:Rhta  :)R=R6;RRRRRRRRRRRRRRRRRRRRRRRRRRRR
RRRRRRRRRRRRb8C0:ERRaQh )t R(:=RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR
RRRRRRRRR2RR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR
RRRRRRRRsbF0R5RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR
RRRRRRRRRRRRRRqRRR:MRHR8#0_oDFHPO_CFO0sH5I8-0E4FR8IFM0R;j2RRR
RRRRRRRRRORRD:	RRRHM#_08DHFoOR;RRRRRRRRRRRRRRRRRRRRRRRRRRR
RRRRRRRRRRRRARRR:FRk0#_08DHFoOC_POs0F58IH04E-RI8FMR0FjR2R
RRRRRRRRRRRRR2;RRRR
R--Ns00H0LkCCR8OsDNNF0HMFRVsHR#MCoDRk#FsROC8HC#oNMIsRC
RRRRRNRR0H0sLCk0RM#$_HLkDM0H_R8k:0R#soHM;R
RRRRRR0RN0LsHkR0C#_$MLDkH0_HM8FkRVWR7jbd_H_bCsRCo:MRC0$H0RRH#"NIC	R";RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR
RRR8CMRj7WdH_bbsC_C
o;
ONsECH0Os0kC0RsDVRFRj7WdH_bbsC_CHoR#-

-0RN0LsHkR0C8DCON0sNHRFMVRFs#oHMD#CRFOksCCR8#MHoICNsR0
N0LsHkR0C#_$MLDkH0_HM8:kRRs#0H;Mo
0N0skHL0#CR$LM_k0HDH8M_kVRFRDs0RN:RsHOE00COkRsCH"#RI	CN"
;
-w-RF#sRHDMoCFR#kCsOR,7WRONsECH0Os0kCER#F8kDRRLC8lkl$0
N0LsHkR0C#_$MLODN	F_LGRR:LDFFC;NM
0N0skHL0#CR$LM_D	NO_GLFRRFVsR0D:sRNO0EHCkO0sHCR#sR0k
C;
oLCH
M
CRM8s;0D
-
--------------------------------------------------------------------------
---S-S HM00N$RMN8RsHOE00COkRsCVRFs7qW_1wYvQBwma1p_4w_7R-R----------------
----------------------------------------------------------------------------
D

HNLssQ$R ,  Rj7Wdk;
#QCR 3  #_08DHFoO4_4nNc3D
D;kR#CHCCC38#0_oDFHkO_Mo#HM3C8N;DD
Ck#RCHCC03#8F_Do_HON0sHED3ND
;RkR#C8dIj3j8IdF_OlMbFC#M03DND;


S0CMHR0$7NW_#V$lHOVF0#D_4V_8R
H#SCSoMHCsO
R5S8SSN_0NHIM_HE80RRS:Q hatR ):U=R;S
SS08NNk_F0H_I8R0ESQ:Rhta  :)R=nR4;S
SSb8C0SERSQ:Rhta  :)R=;RU
SSSC_sslCF8R:SSRaQh )t RR:=4S;
S#Ss0F_l8SCRSQ:Rhta  :)R=;R4
SSSLC$0_8FsCSsRSQ:Rhta  :)R=
RjS2SS;S
Sb0FsRS5
SDSO	SRSSH:RM0R#8F_Do;HO
SSSs_#0MSRSSH:RM0R#8F_Do;HO
SSSbEk#_JsC_SMRSH:RM0R#8F_Do;HO
SSSV#DkER_MSRS:H#MR0D8_FOoH;S
SSbbF_JsC_SMRSH:RM0R#8F_Do;HO
SSS8oHN_SMRSRS:H#MR0D8_FOoH;S
SS_NCDCCPDRRRRRS:HRMR#_08DHFoOC_POs0F50LH_8IH08E5CEb02R-48MFI0jFR2
;RSNSSVE_0sEC#RSRR:MRHR0R#8F_Do_HOP0COFLs5HI0_HE805b8C0-E24FR8IFM0R;j2RS
SS08NNM_HR:SSRRHM#_08DHFoOC_POs0F508NNM_H_8IH04E-RI8FMR0Fj
2;SsSS8N_80SNRSH:RM0R#8F_Do_HOP0COFls5NlGHk8l5N_0NHIM_HE80,NR80FN_kI0_HE802R-48MFI0jFR2S;
SCSI_SMRSRS:FRk0#_08DHFoOS;
SlSCbR0$S:SSR0FkR8#0_oDFH
O;SNSSD#lF0l_CbR0$SF:Rk#0R0D8_FOoH;S
SSDENVk_VDSDRSF:Rk#0R0D8_FOoH;S
SSlNDF_#0VDkDRRS:FRk0#_08DHFoOS;
SkSVDSDRSRS:FRk0#_08DHFoOS;
SNSslk_VDSDRSF:Rk#0R0D8_FOoH;S
SSsCsFSsRSRS:FRk0#_08DHFoOS;
SNSbsI0_8SRS:kRF00R#8F_Do;HO
SSSI8s_NR0NSRS:FRk0#_08DHFoOC_POs0F5GlNHllk508NNM_H_8IH0RE,8NN0_0Fk_8IH0-E24FR8IFM0R;j2
SSSINs_8R8sSRS:FRk0#_08DHFoOC_POs0F50LH_8IH08E5CEb02R-48MFI0jFR2S;
S8Ss_8N8sSRS:kRF00R#8F_Do_HOP0COFLs5HI0_HE805b8C0-E24FR8IFM0R;j2
SSS8NN0_0FkR:SSR0FkR8#0_oDFHPO_CFO0sN580FN_kI0_HE80-84RF0IMF2Rj
SSS2
;
-N-R0H0sLCk0RO8CDNNs0MHFRsVFRM#HoRDC#sFkO8CRCo#HMsINCR
RRRRRR0RN0LsHkR0C#_$MLDkH0_HM8:kRRs#0H;Mo
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kVRFR_7WNl#$VFHVO_0D#84_VRR:CHM00H$R#IR"C"N	;
RR
MSC8WR7_$N#lVVHFDO0__#48
V;Rs
NO0EHCkO0ssCR0FDRVWR7_$N#lVVHFDO0__#48HVR#-

-0RN0LsHkR0C8DCON0sNHRFMVRFs#oHMD#CRFOksCCR8#MHoICNsR0
N0LsHkR0C#_$MLDkH0_HM8:kRRs#0H;Mo
0N0skHL0#CR$LM_k0HDH8M_kVRFRDs0RN:RsHOE00COkRsCH"#RI	CN"
;
-w-RF#sRHDMoCFR#kCsOR,7WRONsECH0Os0kCER#F8kDRRLC8lkl$0
N0LsHkR0C#_$MLODN	F_LGRR:LDFFC;NM
0N0skHL0#CR$LM_D	NO_GLFRRFVsR0D:sRNO0EHCkO0sHCR#sR0k
C;S
R
LHCoM

SCRM8s;0D
-

----------------------------------------------------------------------------
H
DLssN$ RQ R ,7dWj;#
kC RQ # 30D8_FOoH_n44cD3NDk;
#HCRC3CC#_08DHFoOM_k#MHoCN83D
D;kR#CHCCC38#0_oDFHNO_sEH03DND;kR
#8CRI3jd8dIj_lOFbCFMM30#N;DD
C

M00H$WR7_$N#lVVHFDO0__#4#HVR#o
SCsMCH
O5S8SSN_0NHIM_HE80RRRR:hSQa  t)=R:R
U;S8SSN_0NF_k0I0H8ERRR:hSQa  t)=R:R;4n
SSS80CbESSSRQ:Shta  :)R=;RU
RRRRRRRRRRRR_NCDCCPDRSRR:RRRhRQa  t)=R:R
c;SNSSVC_DPSCDRRRRRQ:Shta  :)R=;Rc
SSSC_sslCF8RRSS:hSQa  t)=R:R
4;SsSS#l0_FS8CSSR:Q hatR ):4=R;S
SS0L$Cs_F8SCsRRRRRQ:Shta  :)R=
RjSSSS
SSS2R;S
R
RRRRRRsbF0RR5
RRRRRRRRRRRR	ODRRSRR:RRRRHM#_08DHFoO
R;SsSS#M0_RRSRR:RRRRHM#_08DHFoO
R;RRRRRRRRS#bkEC_sJS_MRH:RM0R#8F_DoRHO;S
SSkVD#ME_RRS:H#MR0D8_FOoH;S
SSbbF_JsC_RMS:MRHR8#0_oDFH;OR
SSS8oHN_SMS:MRHR8#0_oDFH
O;S8SSN_0NHRMSR:RRRRHM#_08DHFoOC_POs0FR55RR08NNM_H_8IH0-ERR24RRI8FMR0Fj;R2
RSSRsRR8N_80SNS:MRHR8#0_oDFHPO_CFO0sRR5lHNGl5kl8NN0__HMI0H8E8,RN_0NF_k0I0H8E42-RI8FMR0FjS2;
SSSIMC_S:SRR0FkR8#0_oDFH
O;SCSSl$b0SF:Rk#0R0D8_FOoH;S
SSlNDF_#0C0lb$RS:FRk0#_08DHFoOS;
SNSEDVV_kSDD:kRF00R#8F_Do;HOS
SSSNSSD#lF0k_VD:DRR0FkR8#0_oDFHSO;SSS
SkSVDSDS:kRF00R#8F_Do;HOS
SSSsSSNVl_kSDD:kRF00R#8F_Do;HO
SSSCFsssRS:FRk0#_08DHFoOS;
SNSbsI0_8:SSR0FkR8#0_oDFHSO;S
S
SISSsN_80SNS:kRF00R#8F_Do_HOP0COF5sRRGlNHllk508NNM_H_8IH0RE,8NN0_0Fk_8IH0-E24FR8IFM0R;j2SSR
S8Ss_8N8s:SSR0FkR8#0_oDFHPO_CFO0sRR55HRL0H_I850E80CbER2R-2R4RI8FMR0Fj
2;
SSSINs_8S8sSF:Rk#0R0D8_FOoH_OPC0RFs5RR5L_H0I0H8EC58b20ERRR-482RF0IMF2Rj;S
SS08NNk_F0RRRRF:Rk#0R0D8_FOoH_OPC0RFs5RR58NN0_0Fk_8IH0-ERR24RRI8FMR0Fj
R2
SSS
2SS;-

-0RN0LsHkR0C8DCON0sNHRFMVRFs#oHMD#CRFOksCCR8#MHoICNs
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kRR:#H0sM
o;RRRRRRRRNs00H0LkC$R#Mk_LHHD0Mk_8RRFV7NW_#V$lHOVF0#D_4V_#RC:RM00H$#RHRC"IN;	"R
R
R
RR
8CMR_7WNl#$VFHVO_0D##4_V
;
NEsOHO0C0CksRDs0RRFV7NW_#V$lHOVF0#D_4V_#R
H#
R--Ns00H0LkCCR8OsDNNF0HMFRVsHR#MCoDRk#FsROC8HC#oNMIs
CRNs00H0LkC$R#Mk_LHHD0Mk_8R#:R0MsHoN;
0H0sLCk0RM#$_HLkDM0H_R8kFsVR0:DRRONsECH0Os0kC#RHRC"IN;	"
-
-RswFRM#HoRDC#sFkO7CRWN,RsHOE00COkRsC#kEFDL8RCkR8l
l$Ns00H0LkC$R#MD_LN_O	LRFG:FRLFNDCMN;
0H0sLCk0RM#$_NLDOL	_FFGRV0RsDRR:NEsOHO0C0CksRRH#0Csk;L

CMoH
M
C80RsD
;

----------------------------------------------------------------------------D-
HNLssQ$R ,  Rj7Wdk;
#QCR 3  #_08DHFoO4_4nNc3D
D;kR#CHCCC38#0_oDFHkO_Mo#HM3C8N;DD
Ck#RCHCC03#8F_Do_HON0sHED3ND
;RkR#C8dIj3j8IdF_OlMbFC#M03DND;


S0CMHR0$7VW_HOVF0#D_4V_#R
H#SCSoMHCsO
R5S8SSCEb0RRRR:hRQa  t)=R:R
c;SNSSCC_DPRCD:hRQa  t)=R:R
4;SNSSVC_DPRCD:hRQa  t)=R:R
4;SCSSsls_FR8C:hRQa  t)=R:R
j;SsSS#l0_FR8C:hRQa  t)=R:RSj
S;S2
bSSFRs05S
SS	ODRSSS:MRHR8#0_oDFH
O;SsSS#M0_RSSS:MRHR8#0_oDFH
O;SbSSk_#Es_CJMSRS:MRHR8#0_oDFH
O;SbSSFsb_CMJ_R:SSRRHM#_08DHFoOS;
SHS8NMo_RSSS:MRHR8#0_oDFH
O;SISSCR_MS:SSR0FkR8#0_oDFH
O;SCSSl$b0RSSS:kRF00R#8F_Do;HO
SSSNFDl#C0_l$b0RRS:FRk0#_08DHFoOS;
SNSEDVV_kRDDSRS:FRk0#_08DHFoOS;
SDSNl0F#_DVkD:RSR0FkR8#0_oDFH
O;SVSSkRDDS:SSR0FkR8#0_oDFH
O;SCSSsssFRSSS:kRF00R#8F_Do;HO
SSSINs_8R8sSRS:FRk0#_08DHFoOC_POs0F50LH_8IH08E5CEb02R-48MFI0jFR2S;
S8Ss_8N8sSRS:kRF00R#8F_Do_HOP0COFLs5HI0_HE805b8C0-E24FR8IFM0R
j2S2SS;-

-0RN0LsHkR0C8DCON0sNHRFMVRFs#oHMD#CRFOksCCR8#MHoICNs
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kRR:#H0sM
o;RRRRRRRRNs00H0LkC$R#Mk_LHHD0Mk_8RRFV7VW_HOVF0#D_4V_#RC:RM00H$#RHRC"IN;	"R
R
S8CMR_7WVFHVO_0D##4_V
;
NEsOHO0C0CksRDs0RRFV7VW_HOVF0#D_4V_#R
H#
R--Ns00H0LkCCR8OsDNNF0HMFRVsHR#MCoDRk#FsROC8HC#oNMIs
CRNs00H0LkC$R#Mk_LHHD0Mk_8R#:R0MsHoN;
0H0sLCk0RM#$_HLkDM0H_R8kFsVR0:DRRONsECH0Os0kC#RHRC"IN;	"
-
-RswFRM#HoRDC#sFkO7CRWN,RsHOE00COkRsC#kEFDL8RCkR8l
l$Ns00H0LkC$R#MD_LN_O	LRFG:FRLFNDCMN;
0H0sLCk0RM#$_NLDOL	_FFGRV0RsDRR:NEsOHO0C0CksRRH#0Csk;L

CMoH
M
C80RsD
;
-----------------------------------------------------------------------------S

DsHLNRs$HCCC,IR8j
d;SCk#RCHCC03#8F_Do_HO4c4n3DND;k
S#HCRC3CC#_08DHFoOM_k#MHoCN83D
D;SCk#RCHCC03#8F_Do_HON0sHED3NDS;
kR#C8dIj3j8IdF_OlMbFC#M03DND;

SS0CMHR0$7#W_0	NOOR0DHS#
SMoCCOsHRS5
SCS8bR0ER:RRRaQh )t RR:=US;
SsSCsF_l8:CRRaQh )t RR:=4S;
S#Ss0F_l8:CRRaQh )t RR:=4S
SS
2;SFSbs50R
SSSORD	SRS:H#MR0D8_FOoH;S
SS0s#_SMRSH:RM0R#8F_Do;HO
SSSbEk#_JsC_RMR:MRHR8#0_oDFH
O;SbSSFsb_CMJ_R:RRRRHM#_08DHFoOS;
SCSI_SMRSF:Rk#0R0D8_FOoH;S
SSbCl0S$RSF:Rk#0R0D8_FOoH;S
SSDVkDSRS:kRF00R#8F_Do;HO
SSSCFsssSRS:kRF00R#8F_Do;HO
SSSINs_8S8sRRRR:kRF00R#8F_Do_HOP0COFLs5HI0_HE805b8C0-E24FR8IFM0R;j2
SSSsN8_8R8sSF:Rk#0R0D8_FOoH_OPC05FsL_H0I0H8EC58b20E-84RF0IMF2Rj
SSS2
;
-N-R0H0sLCk0RO8CDNNs0MHFRsVFRM#HoRDC#sFkO8CRCo#HMsINCR
RRRRRR0RN0LsHkR0C#_$MLDkH0_HM8:kRRs#0H;Mo
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kVRFR_7W#O0N	DO0RC:RM00H$#RHRC"IN;	"R
R
S8CMR_7W#O0N	DO0R
;

sSNO0EHCkO0ssCR0FDRVWR7_N#0O0	OD#RH
-
-R0N0skHL08CRCNODsHN0FVMRF#sRHDMoCFR#kCsOR#8CHIoMNRsC
0N0skHL0#CR$LM_k0HDH8M_kRR:#H0sM
o;Ns00H0LkC$R#Mk_LHHD0Mk_8RRFVsR0D:sRNO0EHCkO0sHCR#IR"C"N	;-

-FRwsHR#MCoDRk#FsROC7RW,NEsOHO0C0CksRF#EkRD8L8CRk$ll
0N0skHL0#CR$LM_D	NO_GLFRL:RFCFDN
M;Ns00H0LkC$R#MD_LN_O	LRFGFsVR0:DRRONsECH0Os0kC#RHRk0sC
;
S
S
LHCoMC

Ms8R0
D;
-
--------------------------------------------------------------------------
--DsHLNRs$Q   ,WR7j
d;kR#CQ   38#0_oDFH4O_43ncN;DD
Ck#RCHCC03#8F_Do_HOkHM#o8MC3DND;#
kCCRHC#C30D8_FOoH_HNs0NE3D
D;kR#C8dIj3j8IdF_OlMbFC#M03DND;S

CHM007$RWH_VV0FOD4_#_R8VHS#
SMoCCOsHRS5
SCS8bR0ESRR:Q hatR ):c=R;S
SSsCs_8lFCRR:Q hatR ):j=R;S
SS0s#_8lFCRR:Q hatR ):j=R
SSS2S;
SsbF0
R5SOSSDS	RSRS:H#MR0D8_FOoH;S
SS0s#_SMRSRS:H#MR0D8_FOoH;S
SS#bkEC_sJR_MSRS:H#MR0D8_FOoH;S
SSbbF_JsC_SMRSH:RM0R#8F_Do;HO
SSS8oHN_SMRSRS:H#MR0D8_FOoH;S
SS_NCDCCPDSRS:MRHR8#0_oDFHPO_CFO0sH5L0H_I850E80CbE42-RI8FMR0Fj
2;SNSSVE_0sEC#R:SSRRHM#_08DHFoOC_POs0F50LH_8IH08E5CEb02R-48MFI0jFR2S;
SCSI_SMRSRS:FRk0#_08DHFoOS;
SlSCbR0$S:SSR0FkR8#0_oDFH
O;SNSSD#lF0l_CbR0$SF:Rk#0R0D8_FOoH;S
SSDENVk_VDSDRSF:Rk#0R0D8_FOoH;S
SSlNDF_#0VDkDRRS:FRk0#_08DHFoOS;
SkSVDSDRSRS:FRk0#_08DHFoOS;
SsSCsRFsS:SSR0FkR8#0_oDFH
O;SISSs8_N8SsRSF:Rk#0R0D8_FOoH_OPC05FsL_H0I0H8EC58b20E-84RF0IMF2Rj;S
SS_s8Ns88R:SSR0FkR8#0_oDFHPO_CFO0sH5L0H_I850E80CbE42-RI8FMR0FjS2
S;S2
R--Ns00H0LkCCR8OsDNNF0HMFRVsHR#MCoDRk#FsROC8HC#oNMIsRC
RRRRRNRR0H0sLCk0RM#$_HLkDM0H_R8k:0R#soHM;R
RRRRRR0RN0LsHkR0C#_$MLDkH0_HM8FkRVWR7_VVHFDO0__#48:VRR0CMHR0$H"#RI	CN"R;R
M
C8WR7_VVHFDO0__#48
V;
ONsECH0Os0kC0RsDVRFR_7WVFHVO_0D#84_V#RH
-
-R0N0skHL08CRCNODsHN0FVMRF#sRHDMoCFR#kCsOR#8CHIoMNRsC
0N0skHL0#CR$LM_k0HDH8M_kRR:#H0sM
o;Ns00H0LkC$R#Mk_LHHD0Mk_8RRFVsR0D:sRNO0EHCkO0sHCR#IR"C"N	;-

-FRwsHR#MCoDRk#FsROC7RW,NEsOHO0C0CksRF#EkRD8L8CRk$ll
0N0skHL0#CR$LM_D	NO_GLFRL:RFCFDN
M;Ns00H0LkC$R#MD_LN_O	LRFGFsVR0:DRRONsECH0Os0kC#RHRk0sC
;
LHCoMC

Ms8R0
D;
----------------------------------------------------------------------------D-
HNLssH$RC;CC
Ck#RCHCC03#8F_Do_HO4c4n3DND;#
kCCRHC#C30D8_FOoH_#kMHCoM8D3ND
;
S0CMHR0$7dWj_V#E0osCR
H#SCSoMHCsO
R5SDSSC0MoERR:hzqa)Rqp:c=R
SSS2S;
SsbF0
R5SOSSDS	R:MRHR8#0_oDFH
O;S#SS_RHMSH:RM0R#8F_Do;HO
SSSbM_HRRS:H#MR0D8_FOoH_OPC05FsDoCM04E-RI8FMR0Fj
2;S#SSE0HV_:MRRRHM#_08DHFoOS;
SFSDNM8_RRS:H#MR0D8_FOoH;S
SSFb_kS0R:kRF00R#8F_Do_HOP0COFDs5C0MoER-48MFI0jFR2S
SS
2;
R--Ns00H0LkCCR8OsDNNF0HMFRVsHR#MCoDRk#FsROC8HC#oNMIsRC
RRRRRNRR0H0sLCk0RM#$_HLkDM0H_R8k:0R#soHM;R
RRRRRR0RN0LsHkR0C#_$MLDkH0_HM8FkRVWR7j#d_EsV0C:oRR0CMHR0$H"#RI	CN"R;R
C
SM78RW_jd#0EVs;Co
N

sHOE00COkRsCsR0DF7VRW_jd#0EVsRCoH
#
-N-R0H0sLCk0RO8CDNNs0MHFRsVFRM#HoRDC#sFkO8CRCo#HMsINCNR
0H0sLCk0RM#$_HLkDM0H_R8k:0R#soHM;0
N0LsHkR0C#_$MLDkH0_HM8FkRV0RsDRR:NEsOHO0C0CksRRH#"NIC	
";
R--wRFs#oHMD#CRFOksCWR7,sRNO0EHCkO0s#CREDFk8CRLRl8klN$
0H0sLCk0RM#$_NLDOL	_F:GRRFLFDMCN;0
N0LsHkR0C#_$MLODN	F_LGVRFRDs0RN:RsHOE00COkRsCH0#Rs;kC
C
Lo
HM
8CMRDs0;SSSRRR

------------------------------------------------------------------------------
--S-- -SM00H$MRN8sRNO0EHCkO0sVCRF7sRW_jdp)w1_h7BaRmRR-R-----------------
----------------------------------------------------------------------------D-
HNLssH$RC;CC
Ck#RCHCC03#8F_Do_HO4c4n3DND;#
kCCRHC#C30D8_FOoH_#kMHCoM8D3ND
;
S0CMHR0$7dWj_#DVsO_8MR0FHS#
SMoCCOsHRS5
SHSI8R0E:hRQa  t)=R:RSd
S;S2
bSSFRs05S
SS08NNSRS:MRHR8#0_oDFHPO_CFO0sH5I8-0E4FR8IFM0R;j2
SSSOMFk0F_0RRS:H#MR0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2S;
SFSDNS8RSH:RM0R#8F_Do;HO
SSSORCMSRS:H#MR0D8_FOoH;S
SS	ODR:SSRRHM#_08DHFoOS;
SCSs#RC0SRS:H#MR0D8_FOoH;S
SSkOFMS0RSF:Rk#0R0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2S;
SCS0s0OMR:SSR0FkR8#0_oDFHSO
S;S2
R--Ns00H0LkCCR8OsDNNF0HMFRVsHR#MCoDRk#FsROC8HC#oNMIsRC
RRRRRNRR0H0sLCk0RM#$_HLkDM0H_R8k:0R#soHM;R
RRRRRR0RN0LsHkR0C#_$MLDkH0_HM8FkRVWR7jDd_V_#s80OMFRR:CHM00H$R#IR"C"N	;
RR
MSC8WR7jDd_V_#s80OMF
;

ONsECH0Os0kC0RsDVRFRj7WdV_D#8s_OFM0R
H#
R--Ns00H0LkCCR8OsDNNF0HMFRVsHR#MCoDRk#FsROC8HC#oNMIs
CRNs00H0LkC$R#Mk_LHHD0Mk_8R#:R0MsHoN;
0H0sLCk0RM#$_HLkDM0H_R8kFsVR0:DRRONsECH0Os0kC#RHRC"IN;	"
-
-RswFRM#HoRDC#sFkO7CRWN,RsHOE00COkRsC#kEFDL8RCkR8l
l$Ns00H0LkC$R#MD_LN_O	LRFG:FRLFNDCMN;
0H0sLCk0RM#$_NLDOL	_FFGRV0RsDRR:NEsOHO0C0CksRRH#0Csk;


LHCoMC

Ms8R0
D;
-
--------------------------------------------------------------------------
--DsHLNRs$HCCC;#
kCCRHC#C30D8_FOoH_n44cD3NDk;
#HCRC3CC#_08DHFoOM_k#MHoCN83D
D;
0CMHR0$7dWj_#DVsO_#MR0FHo#
CsMCH
O5SHSI8S0ESQ:Rhta  :)R=;Rd
OSSF0kM_R0FSQ:Rhta  :)R=
RdS;S2
bSSF5s0RS
SS08NNSRS:MRHR8#0_oDFHPO_CFO0sH5I8-0E4FR8IFM0R;j2
SSSD8FNR:SSRRHM#_08DHFoOS;
SCSOMSRS:MRHR8#0_oDFH
O;SOSSDS	RSH:RM0R#8F_Do;HO
SSSsCC#0SRS:MRHR8#0_oDFH
O;SOSSF0kMR:SSR0FkR8#0_oDFHPO_CFO0sH5I8-0E4FR8IFM0R;j2
SSS0OCsMS0RSF:Rk#0R0D8_FOoH
RRRR2SS;-

-0RN0LsHkR0C8DCON0sNHRFMVRFs#oHMD#CRFOksCCR8#MHoICNs
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kRR:#H0sM
o;RRRRRRRRNs00H0LkC$R#Mk_LHHD0Mk_8RRFV7dWj_#DVsO_#MR0F:MRC0$H0RRH#"NIC	R";RC

M78RW_jdDsV#_M#O0
F;
s
NO0EHCkO0ssCR0FDRVWR7jDd_V_#s#0OMF#RH
-
-R0N0skHL08CRCNODsHN0FVMRF#sRHDMoCFR#kCsOR#8CHIoMNRsC
0N0skHL0#CR$LM_k0HDH8M_kRR:#H0sM
o;Ns00H0LkC$R#Mk_LHHD0Mk_8RRFVsR0D:sRNO0EHCkO0sHCR#IR"C"N	;-

-FRwsHR#MCoDRk#FsROC7RW,NEsOHO0C0CksRF#EkRD8L8CRk$ll
0N0skHL0#CR$LM_D	NO_GLFRL:RFCFDN
M;Ns00H0LkC$R#MD_LN_O	LRFGFsVR0:DRRONsECH0Os0kC#RHRk0sC
;
LHCoMC

Ms8R0
D;
-
--------------------------------------------------------------------------
--
LDHs$NsR Q  k;
#QCR 3  #_08DHFoO4_4nNc3D
D;kR#CQ   38#0_oDFHkO_Mo#HM3C8N;DD
Ck#R Q  03#8F_Do_HON0sHED3ND
;
S0CMHR0$7dWj_osC_b#_D#RH
oSSCsMCH5ORRS
SS8IH0RERRRRRRQ:Rhta  :)R=;Rd
RRRRSRSsCC#0N_PDRkC:hRQa  t):RR=RR(
SSS2S;
SsbF0
R5S8SSRRRRR:RRRRHM#_08DHFoOC_POs0F58IH04E-RI8FMR0Fj
2;SOSSDR	RR:RRRRHM#_08DHFoOS;
SCSs#_C0MRR:H#MR0D8_FOoH;S
SSNCMLRDCRH:RM0R#8F_Do;HO
SSSJRRRRRRR:kRF00R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj
SSS2
;
-N-R0H0sLCk0RO8CDNNs0MHFRsVFRM#HoRDC#sFkO8CRCo#HMsINCR
RRRRRR0RN0LsHkR0C#_$MLDkH0_HM8:kRRs#0H;Mo
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kVRFRj7WdC_so__#b:DRR0CMHR0$H"#RI	CN"R;R
C
SM88RI_jds_Co#D_b;N

sHOE00COkRsCsR0DF8VRI_jds_Co#D_bRRH#
R--Ns00H0LkCCR8OsDNNF0HMFRVsHR#MCoDRk#FsROC8HC#oNMIs
CRNs00H0LkC$R#Mk_LHHD0Mk_8R#:R0MsHoN;
0H0sLCk0RM#$_HLkDM0H_R8kFsVR0:DRRONsECH0Os0kC#RHRC"IN;	"
-
-RswFRM#HoRDC#sFkO7CRWN,RsHOE00COkRsC#kEFDL8RCkR8l
l$Ns00H0LkC$R#MD_LN_O	LRFG:FRLFNDCMN;
0H0sLCk0RM#$_NLDOL	_FFGRV0RsDRR:NEsOHO0C0CksRRH#0Csk;L

CMoH
M
C80RsD
;
-----------------------------------------------------------------------------D

HNLssH$RC;CC
Ck#RCHCC03#8F_Do_HO4c4n3DND;#
kCCRHC#C30D8_FOoH_#kMHCoM8D3ND
;
S0CMHR0$7dWj_#DVsb_k8HMR#S
SoCCMsRHO5S
SS8IH0:ERRaQh )t RR:=US
SS
2;SFSbs50R
SSSkMb8RRS:H#MR0D8_FOoH;S
SSMOCRRS:H#MR0D8_FOoH;S
SS	ODRRS:H#MR0D8_FOoH;S
SS#sCCS0R:MRHR8#0_oDFH
O;SOSSF0kMRRS:FRk0#_08DHFoOC_POs0F58IH04E-RI8FMR0Fj
2;S0SSCMsO0:RRR0FkR8#0_oDFHSO
S;S2
R--Ns00H0LkCCR8OsDNNF0HMFRVsHR#MCoDRk#FsROC8HC#oNMIsRC
RRRRRNRR0H0sLCk0RM#$_HLkDM0H_R8k:0R#soHM;R
RRRRRR0RN0LsHkR0C#_$MLDkH0_HM8FkRVWR7jDd_V_#skMb8RC:RM00H$#RHRC"IN;	"R
R
S8CMRj8IdV_D#ks_b;8M
N

sHOE00COkRsCsR0DF8VRI_jdDsV#_8kbM#RH
-
-R0N0skHL08CRCNODsHN0FVMRF#sRHDMoCFR#kCsOR#8CHIoMNRsC
0N0skHL0#CR$LM_k0HDH8M_kRR:#H0sM
o;Ns00H0LkC$R#Mk_LHHD0Mk_8RRFVsR0D:sRNO0EHCkO0sHCR#IR"C"N	;-

-FRwsHR#MCoDRk#FsROC7RW,NEsOHO0C0CksRF#EkRD8L8CRk$ll
0N0skHL0#CR$LM_D	NO_GLFRL:RFCFDN
M;Ns00H0LkC$R#MD_LN_O	LRFGFsVR0:DRRONsECH0Os0kC#RHRk0sCS;
RR
R
oLCH
M
CRM8s;0D
-

----------------------------------------------------------------------------
DS
HNLssH$RC;CC
Ck#RCHCC03#8F_Do_HO4c4n3DND;#
kCCRHC#C30D8_FOoH_#kMHCoM8D3ND
;
S0CMHR0$7dWj_#DVsF_DNH8R#S
SoCCMsRHO5S
SS8IH0:ERRaQh )t RR:=d
2;SFSbs50R
SSS8NN0RRS:H#MR0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2S;
SFSDNS8R:MRHR8#0_oDFH
O;SOSSCSMR:MRHR8#0_oDFH
O;SOSSDS	R:MRHR8#0_oDFH
O;SsSSC0#CRRS:H#MR0D8_FOoH;S
SSkOFMS0R:kRF00R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj
SSS2-;
-0RN0LsHkR0C8DCON0sNHRFMVRFs#oHMD#CRFOksCCR8#MHoICNs
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kRR:#H0sM
o;RRRRRRRRNs00H0LkC$R#Mk_LHHD0Mk_8RRFV7dWj_#DVsF_DN:8RR0CMHR0$H"#RI	CN"R;R
C
SM88RI_jdDsV#_NDF8
;

ONsECH0Os0kC0RsDVRFRj8IdV_D#Ds_FRN8H
#
-N-R0H0sLCk0RO8CDNNs0MHFRsVFRM#HoRDC#sFkO8CRCo#HMsINCNR
0H0sLCk0RM#$_HLkDM0H_R8k:0R#soHM;0
N0LsHkR0C#_$MLDkH0_HM8FkRV0RsDRR:NEsOHO0C0CksRRH#"NIC	
";
R--wRFs#oHMD#CRFOksCWR7,sRNO0EHCkO0s#CREDFk8CRLRl8klN$
0H0sLCk0RM#$_NLDOL	_F:GRRFLFDMCN;0
N0LsHkR0C#_$MLODN	F_LGVRFRDs0RN:RsHOE00COkRsCH0#Rs;kC
C
Lo
HM
8CMRDs0;-

----------------------------------------------------------------------------
S------S0 MHR0$NRM8NEsOHO0C0CksRsVFRj7WdQ_AB_a)1aBhmRRRR------------------
----------------------------------------------------------------------------
LDHs$NsRCHCCk;
#RCRHCCC38#0_oDFH4O_43ncN;DD
Ck#RCHCC03#8F_Do_HOkHM#o8MC3DND;S

CHM007$RW_jdL0HOsO_#MR0FHS#
SMoCCOsHRS5
SHSI8R0ESRR:Q hatR ):.=R;S
SSkOFM00_FRR:Q hatR ):.=R
SSS2S;
SsbF0
R5S8SSNR0NSH:RM0R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj;S
SS_kb8SMR:MRHR8#0_oDFH
O;SDSSFRN8SH:RM0R#8F_Do;HO
SSSORCMSH:RM0R#8F_Do;HO
SSSORD	SH:RM0R#8F_Do;HO
SSSsCC#0:RSRRHM#_08DHFoOS;
SFSOkRM0SF:Rk#0R0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2S;
SCS0s0OMRRS:FRk0#_08DHFoOS
SS
2;-N-R0H0sLCk0RO8CDNNs0MHFRsVFRM#HoRDC#sFkO8CRCo#HMsINCR
RRRRRR0RN0LsHkR0C#_$MLDkH0_HM8:kRRs#0H;Mo
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kVRFRj7WdH_LO_0s#0OMFRR:CHM00H$R#IR"C"N	;
RR
MSC8WR7jLd_HsO0_M#O0
F;
ONsECH0Os0kC0RsDVRFRj7WdH_LO_0s#0OMF#RH
-
-R0N0skHL08CRCNODsHN0FVMRF#sRHDMoCFR#kCsOR#8CHIoMNRsC
0N0skHL0#CR$LM_k0HDH8M_kRR:#H0sM
o;Ns00H0LkC$R#Mk_LHHD0Mk_8RRFVsR0D:sRNO0EHCkO0sHCR#IR"C"N	;-

-FRwsHR#MCoDRk#FsROC7RW,NEsOHO0C0CksRF#EkRD8L8CRk$ll
0N0skHL0#CR$LM_D	NO_GLFRL:RFCFDN
M;Ns00H0LkC$R#MD_LN_O	LRFGFsVR0:DRRONsECH0Os0kC#RHRk0sC
;
LHCoM

SCRM8s;0D
-
--------------------------------------------------------------------------
--
LDHs$NsRCHCCk;
#RCRHCCC38#0_oDFH4O_43ncN;DD
Ck#RCHCC03#8F_Do_HOkHM#o8MC3DND;S

CHM007$RW_jdL0HOsO_8MR0FH
#RSCSoMHCsO
R5SISSHE80RH:SMo0CC:sS=
R.S2SS;S
Sb0FsRS5
SNS80:NSRRHMS8#0_oDFHPO_CFO0sH5I8-0E4FR8IFM0R;j2
SSSOMFk0F_0:MRHR0S#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj;S
SS_kb8:MSRRHMS8#0_oDFH
O;SDSSFSN8:MRHR0S#8F_Do;HO
SSSOSCMSH:RM#RS0D8_FOoH;S
SS	ODSRS:HSMR#_08DHFoOS;
SCSs#SC0:MRHR0S#8F_Do;HOS
SSSOSSF0kMSF:RkS0R#_08DHFoOC_POs0F58IH04E-RI8FMR0Fj
2;S0SSCMsO0RS:FRk0S8#0_oDFHSO
S;S2
R--Ns00H0LkCCR8OsDNNF0HMFRVsHR#MCoDRk#FsROC8HC#oNMIsRC
RRRRRNRR0H0sLCk0RM#$_HLkDM0H_R8k:0R#soHM;R
RRRRRR0RN0LsHkR0C#_$MLDkH0_HM8FkRVWR7jLd_HsO0_M8O0:FRR0CMHR0$H"#RI	CN"R;R
C
SM78RW_jdL0HOsO_8M;0FRN

sHOE00COkRsCsR0DF7VRW_jdL0HOsO_8MR0FH
#
-N-R0H0sLCk0RO8CDNNs0MHFRsVFRM#HoRDC#sFkO8CRCo#HMsINCNR
0H0sLCk0RM#$_HLkDM0H_R8k:0R#soHM;0
N0LsHkR0C#_$MLDkH0_HM8FkRV0RsDRR:NEsOHO0C0CksRRH#"NIC	
";
R--wRFs#oHMD#CRFOksCWR7,sRNO0EHCkO0s#CREDFk8CRLRl8klN$
0H0sLCk0RM#$_NLDOL	_F:GRRFLFDMCN;0
N0LsHkR0C#_$MLODN	F_LGVRFRDs0RN:RsHOE00COkRsCH0#Rs;kC


SLHCoM

SCRM8s;0D
-
--------------------------------------------------------------------------
-----S-S-- HM00N$RMN8RsHOE00COkRsCVRFs7dWj_BAQa7)_ 7Bm RRRR-R---------------
--------------------------------------------------------------------------
--DsHLNRs$HCCC;#
kCCRHC#C30D8_FOoH_n44cD3NDk;
#HCRC3CC#_08DHFoOM_k#MHoCN83D
D;kR#CHCCC38#0_oDFHNO_sEH03DND;#
kCCRHCMC3kslCH#O_0N83D
D;
MSC0$H0Rj7WdH_LO_0s8FCO8HCR#S
SoCCMs5HO
SSSI0H8EQ:Rhta  :)R=
RdS2SS;S
Sb0FsRS5
SNS80SNS:MRHR0S#8F_Do_HOP0COF5s5I0H8E2-4RI8FMR0Fj
2;SkSSbM_8SRS:HSMR#_08DHFoOS;
SFSDNS8S:MRHR0S#8F_Do;HO
SSSOSCMSRS:HSMR#_08DHFoOS;SSS
SS	ODS:SSRRHMS8#0_oDFH
O;SsSSC0#CSRS:HSMR#_08DHFoOS;
SFSOk_M08SCO:0FkS8#0_oDFHPO_CFO0s.55*H*I8-0E482RF0IMF2Rj;S
SSs0COSM0SF:RkS0R#_08DHFoOSSS
SSS2
;
-N-R0H0sLCk0RO8CDNNs0MHFRsVFRM#HoRDC#sFkO8CRCo#HMsINCR
RRRRRR0RN0LsHkR0C#_$MLDkH0_HM8:kRRs#0H;Mo
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kVRFRj7WdH_LO_0s8FCO8:CRR0CMHR0$H"#RI	CN"R;R
C
SM78RW_jdL0HOsC_8OCF8;N

sHOE00COkRsCsR0DF7VRW_jdL0HOsC_8OCF8R
H#-N-R0H0sLCk0RO8CDNNs0MHFRsVFRM#HoRDC#sFkO8CRCo#HMsINCNR
0H0sLCk0RM#$_HLkDM0H_R8k:0R#soHM;0
N0LsHkR0C#_$MLDkH0_HM8FkRV0RsDRR:NEsOHO0C0CksRRH#"NIC	
";
R--wRFs#oHMD#CRFOksCWR7,sRNO0EHCkO0s#CREDFk8CRLRl8klN$
0H0sLCk0RM#$_NLDOL	_F:GRRFLFDMCN;0
N0LsHkR0C#_$MLODN	F_LGVRFRDs0RN:RsHOE00COkRsCH0#Rs;kC
C
Lo
HMSM
C80RsD
;
------------------------------------------------------------------------------
-S----MS 0$H0R8NMRONsECH0Os0kCFRVsWR7jBd_h_a)tY)qRRRR-----------------
-------------------------------------------------------------------------------H
DLssN$ RQ ; R
Ck#RRRRR Q  0318F_po_HO4c4n3pqpRk;
#RCRRQRR 3  1_08pHFoOs_qH30EqRpp;#
kCRRRR RQ 1 30p8_FOoH_#zMHCoM8p3qp
R;
0CMHR0$7dWj_0OMss_oNH$R#S
SoCCMsRHO5S
SS8IH0:ERRaQh )t RR:=dS
SS
2;SFSbs50R
SSSORD	SRRRRH:RM0R#8F_Do;HO
SSSsCC#0SRS:MRHR8#0_oDFH
O;SOSSCSMRSH:RM0R#8F_Do;HO
SSSOMFk0SRS:kRF00R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj;S
SSO8CF_8CFRk0SF:Rk#0R0D8_FOoH_OPC05Fs.I**HE80-84RF0IMF2Rj
SSS2-;
-0RN0LsHkR0C8DCON0sNHRFMVRFs#oHMD#CRFOksCCR8#MHoICNs
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kRR:#H0sM
o;RRRRRRRRNs00H0LkC$R#Mk_LHHD0Mk_8RRFV7dWj_0OMss_oN:$RR0CMHR0$H"#RI	CN"R;R
C
SM78RW_jdOsM0_Nos$
R;
ONsECH0Os0kC0RsDVRFRj7WdM_O0os_sRN$H-#
-0RN0LsHkR0C8DCON0sNHRFMVRFs#oHMD#CRFOksCCR8#MHoICNsR0
N0LsHkR0C#_$MLDkH0_HM8:kRRs#0H;Mo
0N0skHL0#CR$LM_k0HDH8M_kVRFRDs0RN:RsHOE00COkRsCH"#RI	CN"
;
-w-RF#sRHDMoCFR#kCsOR,7WRONsECH0Os0kCER#F8kDRRLC8lkl$0
N0LsHkR0C#_$MLODN	F_LGRR:LDFFC;NM
0N0skHL0#CR$LM_D	NO_GLFRRFVsR0D:sRNO0EHCkO0sHCR#sR0k
C;
C
Lo
HMSM
C80RsDRR;
-
--------------------------------------------------------------------------
-----S-S-- HM00N$RMN8RsHOE00COkRsCVRFs7dWj_7zuha_B)RRRR---------------------
--------------------------------------------------------------------------
--DsHLNRs$Q   ;#
kC RQ # 30D8_FOoH_n44cD3NDk;
#QCR 3  #_08DHFoOM_k#MHoCN83D
D;
MSC0$H0Rj7Wdb_k8OM_0HsR#S
SoCCMs5HO
SSSI0H8ERR:Q hatR ):U=R
SSS2
;RSFSbs
05S8SSNS0N:MRHR#RS0D8_FOoH_OPC05FsRH5I8-0E482RF0IMF2Rj;S
SS_kb8:MSRRHMR0S#8F_Do;HO
SSSD8FNSH:RMSRR#_08DHFoOS;
SCSOM:SSRRHMR0S#8F_Do;HO
SSSOSD	SH:RMSRR#_08DHFoOS;
SCSs#SC0:MRHR#RS0D8_FOoH;S
SSkOFM:0SR0FkR0S#8F_Do_HOP0COF5s5R8IH04E-2FR8IFM0R;j2
SSS0OCsM:0SR0FkR0S#8F_Do
HOS2SS;-
-R0N0skHL08CRCNODsHN0FVMRF#sRHDMoCFR#kCsOR#8CHIoMN
sCRRRRRRRRNs00H0LkC$R#Mk_LHHD0Mk_8R#:R0MsHoR;
RRRRRNRR0H0sLCk0RM#$_HLkDM0H_R8kF7VRW_jdkMb8_sO0RC:RM00H$#RHRC"IN;	"R
R
S8CMRj7Wdb_k8OM_0
s;
ONsECH0Os0kC0RsDVRFRj7Wdb_k8OM_0HsR#-R
-0RN0LsHkR0C8DCON0sNHRFMVRFs#oHMD#CRFOksCCR8#MHoICNsR0
N0LsHkR0C#_$MLDkH0_HM8:kRRs#0H;Mo
0N0skHL0#CR$LM_k0HDH8M_kVRFRDs0RN:RsHOE00COkRsCH"#RI	CN"
;
-w-RF#sRHDMoCFR#kCsOR,7WRONsECH0Os0kCER#F8kDRRLC8lkl$0
N0LsHkR0C#_$MLODN	F_LGRR:LDFFC;NM
0N0skHL0#CR$LM_D	NO_GLFRRFVsR0D:sRNO0EHCkO0sHCR#sR0k
C;
oLCH
M
CRM8s;0D
----------------------------------------------------------------------------
-
DsHLNRs$Q   ,j8Idk;
#QCR 3  #_08DHFoO4_4nNc3D
D;kR#CQ   38#0_oDFHNO_sEH03DND;#
kC RQ # 30D8_FOoH_#kMHCoM8D3NDk;
#8CRI3jd8dIj_lOFbCFMM30#N;DD
M
C0$H0R_7WVFHVO_0D##._V#RH
CSoMHCsOS5
SCS8bR0ESRS:Q hatR ):U=R;S
SS#bkEC_N_DDPRQ:Rhta  :)R=;R.
SSSbEk#__NVDRPD:hRQa  t)=R:R
.;SbSSFNb_CP_DD:RRRaQh )t RR:=.S;
SFSbbV_N_DDPRRR:Q hatR ):.=R;S
SSsCs_8lFCRRRRQ:Rhta  :)R=;Rj
SSSbEk#_M#$ORRR:hRQa  t)=R:R
4;SbSSF#b_$RMOR:RRRaQh )t RR:=4S;
S#Ss0F_l8RCRRRR:Q hatR ):j=R;S
SS00#_8lFCRRRRRRRRQ:Rhta  :)R=RRj
SSS
SSS2R;S
SSS

S
RRRRRbRRFRs05RR
RRRRRRRRRORRDb	_kR#ESRR:H#MR0D8_FOoHRS;
SDSO	F_bb:SRRRHM#_08DHFoOR;
RRRRRSRRs_#0MRRS:MRHR8#0_oDFH;OR
RRRRRRRRkSb#sE_CMJ_SRR:H#MR0D8_FOoHRS;
SFSbbC_sJS_MRH:RM0R#8F_DoRHO;S
SS_ICMRSS:kRF00R#8F_Do;HO
SSSbEk#_bCl0R$S:kRF00R#8F_Do;HO
SSSbEk#_SNCRF:Rk#0R0D8_FOoH;S
SS#bkEV_ESRR:FRk0#_08DHFoOS;
SkSb#NE_V:SRR0FkR8#0_oDFH
O;SbSSk_#EVDkDSRR:FRk0#_08DHFoOS;
SkSb#CE_sssFSRR:FRk0#_08DHFoOS;
SFSbbl_CbS0$RF:Rk#0R0D8_FOoH;S
SSbbF_SNCRF:Rk#0R0D8_FOoH;S
SSbbF_SEVRF:Rk#0R0D8_FOoH;S
SSbbF_SNVRF:Rk#0R0D8_FOoH;S
SSbbF_DVkD:SRR0FkR8#0_oDFH
O;SSRSb_FbCFsss:SRR0FkR8#0_oDFH
O;SISSs8_N8RsS:kRF00R#8F_Do_HOP0COFRs55HRL0H_I850E80CbER2R-2R4RI8FMR0Fj
2;SsSS88_N8RsS:kRF00R#8F_Do_HOP0COFRs55HRL0H_I850E80CbE-2RRR428MFI0jFR2S;
SkSb#IE_F_s8OMFk0RR:FRk0#_08DHFoOC_POs0F50LH_8IH08E5CEb0+-424FR8IFM0R;j2
RRRRRRRRRRRRRRRRRRRRRRRRbbF_sIF8F_OkRM0:kRF00R#8F_Do_HOP0COFLs5HI0_HE805b8C04E+2R-48MFI0jFR2R;
RRRRRRRRRRRRRRRRRRRRR0RRCR#0:MRHR8#0_oDFH
O
S;S2
-
-R0N0skHL08CRCNODsHN0FVMRF#sRHDMoCFR#kCsOR#8CHIoMN
sCRRRRRRRRNs00H0LkC$R#Mk_LHHD0Mk_8R#:R0MsHoR;
RRRRRNRR0H0sLCk0RM#$_HLkDM0H_R8kF7VRWH_VV0FOD._#_R#V:MRC0$H0RRH#"NIC	R";RR
SR
R
CRM87VW_HOVF0#D_.V_#R
;R
ONsECH0Os0kC0R#s0kORRFV7VW_HOVF0#D_.V_#RRH#
-
-R0N0skHL08CRCNODsHN0FVMRF#sRHDMoCFR#kCsOR#8CHIoMNRsC
0N0skHL0#CR$LM_k0HDH8M_kRR:#H0sM
o;Ns00H0LkC$R#Mk_LHHD0Mk_8RRFV#k0sO:0RRONsECH0Os0kC#RHRC"IN;	"
-
-RswFRM#HoRDC#sFkO7CRWN,RsHOE00COkRsC#kEFDL8RCkR8l
l$Ns00H0LkC$R#MD_LN_O	LRFG:FRLFNDCMN;
0H0sLCk0RM#$_NLDOL	_FFGRV0R#s0kORN:RsHOE00COkRsCH0#Rs;kC
L

CMoH
C

M#8R0Osk0
;





