--------------------------------------------------
@ES--a1m_am7ptRQBVOkM0MHFRObN	CNo
------------------------------------------------
--
LDHs$NsSCHCCk;
#HCRC3CC#_08DHFoO4_4nNc3D
D;
ObN	CNoS8#0_oDFH1O_AHaR#R

RwRRzahBQRmha1F_0F8poRHORRRRRRR5LRR:ARQaRRRRRRRRRRRRRRR2)z a)#hR0D8_FOoH;R
RRCR
M#8R0D8_FOoH_a1A;b

NNO	oLCRFR8$#_08DHFoOA_1a#RH
-
------------------------------------------------------------------R-
RwRRzahBQRmha1F_0F8poRHORRRRRRR5LRR:ARQaRRRRRRRRRRRRRRR2)z a)#hR0D8_FOoHR
Q1RRRRAQ thR
RRRRRRqRB1L RR
Q1RRRRRRRRRRRRWh] R''jRR=>)z a)'hRj
';RRRRRRRRRRRRWh] R''4RR=>)z a)'hR4
';RRRRRRRR Rh7B q1;R
RRhR 7
;
CRM8#_08DHFoOA_1a
;

=--=========================================================================
==-1-RAq_B)R)Y
=--=========================================================================
==
R
RRHRDLssN$CRHC
C;RRRRkR#CHCCC38#0_oDFH4O_43ncN;DD
RRRRCk#RCHCC03#8F_Do_HOkHM#o8MC3DND;R
RRRR
R
RRCHM001$RAq_B)R)YHu#
FRs05QRRjRR:HRMR#_08DHFoOR;
RRRRRQRR4RR:HRMR#_08DHFoOR;
RRRRRBRRQRR:HRMR#_08DHFoOR;
RRRRRBRRmRR:FRk0R8#0_oDFHROR2C;
M18RAq_B);)Y
0N0skHL0#CR$LM_D	NO_GLFRRFV1BA_qY))RO:RFFlbM0CMRRH#0Csk;N

sHOE00COkRsCVOkMRRFV1BA_qY))R
H##MHoNBDRQM_H0#R:0D8_FOoH:j=''L;
CMoH
FbsO#C#52BQ
CSLoRHM
RSRRRHV5RBQ=4R'')RmRRBQ=jR''02RERCMBHQ_M=0<B
Q;SRRRCCD#R_BQH<M0=jR''S;
RCRRMH8RVR;
R8CMRFbsO#C#;B

m=R<RQ5B_0HMR8NMR2QjRRFs5_BQHRM0NRM8QR42F5sRQNjRMQ8R4
2;RM
C8kRVMRO;
-

-============================================================================-
-R_1AB)q)Yh_Q_XvzR-
-============================================================================
R
RRHRDLssN$CRHC
C;RRRRkR#CHCCC38#0_oDFH4O_43ncN;DD
RRRRCk#RCHCC03#8F_Do_HOkHM#o8MC3DND;C

M00H$AR1_)Bq)QY_hz_vX#RH
MoCCOsH5QB_h:QaL_H0P0COF4s5RI8FMR0Fj:2R=jR"j;"2
RRRRsbF0RR5
RSROsNs$M_HHF0_kR0R:kRF0#RR0D8_FOoH;R
SRsONsH$_M_H0HRMR:MRHR0R#8F_DoRHOR;R2
M
C8AR1_)Bq)QY_hz_vX
;RNs00H0LkC$R#MD_LN_O	LRFGF1VRAq_B)_)YQvh_z:XRRlOFbCFMMH0R#sR0k
C;Rs
NO0EHCkO0sVCRkRMOF1VRAq_B)_)YQvh_zHXR#H
#oDMNRD#CC_O0L#H0R0:#8F_Do_HOP0COF4s5RI8FMR0Fj
2;
oLCHbM
sCFO###5CODC0H_L0O#,N$ss_HHM0M_H2L
SCMoHRR
SR#ONCCR#D0CO_0LH##RH
RSRRIRRERCM""jj=N>Os_s$H0MH_0Fk<j=''S;
RRRRRCIEMjR"4>"=OsNs$M_HHF0_k=0<';4'
RSRRIRRERCM""4j=N>Os_s$H0MH_0Fk<N=Os_s$H0MH_;HM
RSRRIRRERCM""44=N>Os_s$H0MH_0Fk<N=Os_s$H0MH_;HM
RSRRIRRERCMFC0Es=#R>sONsH$_M_H0F<k0=''j;R
SR8CMR#ONCS;
RRRR
RRRCRM8bOsFC;##
RRR#CCDOL0_HR0#<a=Rma_17tpmQ BeB)am5QB_h2Qa;

RCRM8VOkM;
R
-=-==========================================================================-=
-AR1_apzc-R
-============================================================================R

RDRRHNLssH$RC;CC
RRRRCk#RCHCC03#8F_Do_HO4c4n3DND;R
RR#RkCCRHC#C30D8_FOoH_#kMHCoM8D3NDR;
R
RRCHM001$RAz_paHcR#R
RRMoCCOsH5apz_QQhaH:L0C_POs0F5R468MFI0jFR2=R:Rj"jjjjjjjjjjjjjj2j";R
RRsbF0RR5
RSRm:RRR0FkR0R#8F_Do;HO
RSRQRjR:MRHR0R#8F_Do;HO
RSRQR4R:MRHR0R#8F_Do;HO
RSRQR.R:MRHR0R#8F_Do;HO
RSRQRdR:MRHR0R#8F_DoRHOR;R2
M
C8AR1_apzc
;RNs00H0LkC$R#MD_LN_O	LRFGF1VRAz_pa:cRRlOFbCFMMH0R#sR0k
C;Rs
NO0EHCkO0sVCRkRMOF1VRAz_paHcR#H
#oDMNR#lN	#R:0D8_FOoH_OPC05Fs486RF0IMF2Rj;H
#oDMNR0Dk#0:#8F_Do:HO=''j;H
#oDMNR_QdH#M:0D8_FOoH:j=''#;
HNoMD.RQ_:HM#_08DHFoO':=j
';#MHoNQDR4M_H:8#0_oDFH=O:';j'
o#HMRNDQHj_M0:#8F_Do:HO=''j;H
#oDMNRuQhz:a1#_08DHFoOC_POs0F58dRF0IMF2Rj;C
Lo
HM
s
bF#OC#d5Q_,HMQH._M4,Q_,HMQHj_MS2
LHCoMRR
RRRRRRRRR_QdH<MR=dRQ;R
RRRRRRRRRQH._M=R<R;Q.
RRRRRRRRQRR4M_HRR<=Q
4;RRRRRRRRRjRQ_RHM<Q=RjS;
RRRRRNRl#<	R=mRa_71apQmtBBe a5m)p_zaQahQ2R;
RRRRRRRRmD<=k;0#
RSRRRRRRuQhz<a1=_QdH&MRR_Q.H&MRR_Q4H&MRR_QjH
M;SR
SRNRO#QCRhauz1#RH
RSRRIRRERCM"jjjj>"=D#k0<l=RN5#	jV2N0RCsj43jR;M#
RSRRIRRERCM"jjj4>"=D#k0<l=RN5#	4V2N0RCsj43jR;M#
RSRRIRRERCM"4jjj>"=D#k0<l=RN5#	.V2N0RCsj43jR;M#
RSRRIRRERCM"4jj4>"=D#k0<l=RN5#	dV2N0RCsj43jR;M#
RSRRIRRERCM"jj4j>"=D#k0<l=RN5#	cV2N0RCsj43jR;M#
RSRRIRRERCM"jj44>"=D#k0<l=RN5#	6V2N0RCsj43jR;M#
RSRRIRRERCM"4j4j>"=D#k0<l=RN5#	nV2N0RCsj43jR;M#
RSRRIRRERCM"4j44>"=D#k0<l=RN5#	(V2N0RCsj43jR;M#
RSSRERIC"MR4jjj"D=>k<0#=NRl#U	520NVCjsR3Rj4M
#;SRRRRERIC"MR44jj"D=>k<0#=NRl#g	520NVCjsR3Rj4M
#;SRRRRERIC"MR4jj4"D=>k<0#=NRl#4	5jV2N0RCsj43jR;M#
RSRRIRRERCM"44j4>"=D#k0<l=RN5#	4N42Vs0CRjj34#RM;R
SRRRRIMECR4"4j=j">0Dk#R<=l	N#524.NCV0s3RjjM4R#S;
RRRRRCIEM4R"4"j4=k>D0=#<R#lN	d5420NVCjsR3Rj4M
#;SRRRRERIC"MR4j44"D=>k<0#=NRl#4	5cV2N0RCsj43jR;M#
RSRRIRRERCM"4444>"=D#k0<l=RN5#	4N62Vs0CRjj34#RM;R
SRRRRIMECREF0C=s#>0Dk#R<=l	N#5Nj2Vs0CRjj34#RM;R
SRMRC8NRO#
C;RMRC8sRbF#OC#
;RCRM8VOkM;


-=-==========================================================================-=
-AR1_w7wR-
-============================================================================
R
RRHRDLssN$CRHC
C;RRRRkR#CHCCC38#0_oDFH4O_43ncN;DD
RRRRCk#RCHCC03#8F_Do_HOkHM#o8MC3DND;C

M00H$AR1_w7wR
H#RbRRFRs05SR
RRRTRF:RkR0R#_08DHFoOS;
RRR7RH:RM#RR0D8_FOoH;R
SRRBR:MRHR0R#8F_DoRHOR
2;S
RRCRM817A_wRw;
0N0skHL0#CR$LM_D	NO_GLFRRFV17A_w:wRRlOFbCFMMH0R#sR0k
C;Rs
NO0EHCkO0sVCRkRMOF1VRAw_7w#RH
oLCHRM
bOsFC5##BR2
RCRLo
HMSHRRV'RBCMPC0MRN8RRB=4R''ER0CSM
SRRT<7=R;R
RRRRRCRM8H
V;RCRRMb8RsCFO#
#;CRM8RMVkO
;

=--=========================================================================
==-1-RAw_7wR1)
=--=========================================================================
==
RRRRLDHs$NsRCHCCR;
RkRR#HCRC3CC#_08DHFoO4_4nNc3D
D;RRRRkR#CHCCC38#0_oDFHkO_Mo#HM3C8N;DD
M
C0$H0R_1A71ww)#RH
RRRb0FsR
5RRRRR):RRRRHMR8#0_oDFH
O;STRRRRR:FRk0R8#0_oDFH
O;S7RRRRR:HRMR#_08DHFoOS;
RRRBRH:RM#RR0D8_FOoHR;R2
RSR
8CMR_1A71ww)
;RNs00H0LkC$R#MD_LN_O	LRFGF1VRAw_7wR1):FROlMbFCRM0H0#Rs;kC
NR
sHOE00COkRsCVOkMRRFV17A_w)w1R
H#LHCoMb
RsCFO#B#52R
RRoLCHSM
RVRHRCB'P0CMR8NMR=BRR''4RC0EMR
SRRRRH)VRR'=R4E'0CSM
SRRRRRRRR<TR=jR''S;
SRRRCCD#
RSSRRRRRTRRRR<=7R;
RRRRRMRC8VRH;R
RRMRC8VRH;R
RR8CMRFbsO#C#;M
C8VRRk;MO
-

-============================================================================-
-R_1A71ww1-R
-============================================================================R

RDRRHNLssH$RC;CC
RRRRCk#RCHCC03#8F_Do_HO4c4n3DND;R
RR#RkCCRHC#C30D8_FOoH_#kMHCoM8D3ND
;
CHM001$RAw_7wR11HR#
RFRbs50RRR
RRRR1RH:RM#RR0D8_FOoH;R
SRRTR:kRF0#RR0D8_FOoH;R
SRR7R:MRHR0R#8F_Do;HO
RSRB:RRRRHMR8#0_oDFHROR2S;
RCR
M18RAw_7w;11R0
N0LsHkR0C#_$MLODN	F_LGVRFR_1A71ww1RR:ObFlFMMC0#RHRk0sCR;

ONsECH0Os0kCkRVMFORVAR1_w7w1H1R#C
Lo
HMRFbsO#C#5
B2RLRRCMoH
RSRHBVR'CCPMN0RMB8RR'=R40'RE
CMSRRRRVRHR=1RR''40MEC
RSSRRRRRTRRRR<=';4'
RSSRDRC#SC
SRRRRRRRR<TR=;R7
RRRRRRRCRM8H
V;RRRRCRM8H
V;RCRRMb8RsCFO#
#;CRM8RMVkO
;

-
-============================================================================
R--17A_wRw)
=--=========================================================================
==
RRRRLDHs$NsRCHCCR;
RkRR#HCRC3CC#_08DHFoO4_4nNc3D
D;RRRRkR#CHCCC38#0_oDFHkO_Mo#HM3C8N;DD
C

M00H$AR1_w7w)#RH
RRRb0FsR
5RRRRR):RRRRHMR8#0_oDFH
O;STRRRRR:FRk0R8#0_oDFH
O;S7RRRRR:HRMR#_08DHFoOS;
RRRBRH:RM#RR0D8_FOoHR;R2
RSR
8CMR_1A7)ww;NR
0H0sLCk0RM#$_NLDOL	_FFGRVAR1_w7w)RR:ObFlFMMC0#RHRk0sCR;

ONsECH0Os0kCkRVMFORVAR1_w7w)#RH
oLCHRM
bOsFC5##BRR,)
R2RLRRCMoH
RSRH5VRBP'CCRM0NRM8BRR='24'RRm)5C)'P0CMR8NMR=)RR''420RRE
CMSRRRRVRHR=)RR''40MEC
RSSRRRRRTRRRR<=';j'
RSSRDRC#SC
SRRRRRRRR<TR=;R7
RRRRRRRCRM8H
V;RRRRCRM8H
V;RCRRMb8RsCFO#
#;CRM8RMVkO
;

=--=========================================================================
==-1-RAw_7w
1R-=-==========================================================================
=
RRRRDsHLNRs$HCCC;R
RR#RkCCRHC#C30D8_FOoH_n44cD3NDR;
RkRR#HCRC3CC#_08DHFoOM_k#MHoCN83D
D;
0CMHR0$17A_wRw1HR#
RFRbs50RRR
RRRR1RH:RM#RR0D8_FOoH;R
SRRTR:kRF0#RR0D8_FOoH;R
SRR7R:MRHR0R#8F_Do;HO
RSRB:RRRRHMR8#0_oDFHROR2S;
RCR
M18RAw_7wR1;
0N0skHL0#CR$LM_D	NO_GLFRRFV17A_wRw1:FROlMbFCRM0H0#Rs;kC
NR
sHOE00COkRsCVOkMRRFV17A_wRw1HL#
CMoH
sRbF#OC#R5B,RR12R
RRoLCHSM
RVRHR'5BCMPC0MRN8RRB=4R''m2R)1R5'CCPMN0RM18RR'=R4R'2RC0EMR
SRRRRH1VRR'=R4E'0CSM
SRRRRRRRR<TR=4R''S;
SRRRCCD#
RSSRRRRRTRRRR<=7R;
RRRRRMRC8VRH;R
RRMRC8VRH;R
RR8CMRFbsO#C#;M
C8VRRk;MO
-

-============================================================================-
-R_1A7 wwR-
-============================================================================
R
RRHRDLssN$CRHC
C;RRRRkR#CHCCC38#0_oDFH4O_43ncN;DD
RRRRCk#RCHCC03#8F_Do_HOkHM#o8MC3DND;


CHM001$RAw_7wH R#R
RRsbF0RR5
RRRRR R:MRHR0R#8F_DoRHO:'=R]
';STRRRRR:FRk0R8#0_oDFH
O;S7RRRRR:HRMR#_08DHFoOS;
RRRBRH:RM#RR0D8_FOoHR;R2
RSR
8CMR_1A7 ww;NR
0H0sLCk0RM#$_NLDOL	_FFGRVAR1_w7w RR:ObFlFMMC0#RHRk0sCR;

ONsECH0Os0kCkRVMFORVAR1_w7w #RH
oLCHRM
bOsFC5##BR2
RCRLo
HMSHRRV'RBCMPC0MRN8RRB=4R''0RRE
CMSRRRRVRHR= RR''40MEC
RSSRRRRRTRRRR<=7S;
SRRRCRM8H
V;RRRRCRM8H
V;RCRRMb8RsCFO#
#;CRM8RMVkO
;

=--=========================================================================
==-1-RAw_7w) 1R-
-============================================================================
R
RRHRDLssN$CRHC
C;RRRRkR#CHCCC38#0_oDFH4O_43ncN;DD
RRRRCk#RCHCC03#8F_Do_HOkHM#o8MC3DND;


CHM001$RAw_7w) 1R
H#RbRRFRs05RR
R RRRRR:HRMR#_08DHFoO=R:R''];R
RRRR)RH:RM#RR0D8_FOoH;R
SRRTR:kRF0#RR0D8_FOoH;R
SRR7R:MRHR0R#8F_Do;HO
RSRB:RRRRHMR8#0_oDFHROR2S;
RCR
M18RAw_7w) 1;NR
0H0sLCk0RM#$_NLDOL	_FFGRVAR1_w7w R1):FROlMbFCRM0H0#Rs;kC
NR
sHOE00COkRsCVOkMRRFV17A_w1w )#RH
oLCHRM
bOsFC5##BR2
RCRLo
HMSHRRV'RBCMPC0MRN8RRB=4R''ER0CSM
RRRRH VRR'=R40'RERCMRR
SRRRRRVRHR=)RR''40MEC
RSSRRRRRRRRR<TR=jR''S;
SRRRRDRC#SC
SRRRRRRRRTRRRR<=7R;
RRRRRMRC8VRH;R
RRRRRCRM8H
V;RRRRCRM8H
V;RCRRMb8RsCFO#
#;CRM8RMVkO
;

=--=========================================================================
==-1-RAw_7w1 1R-
-============================================================================
R
RRHRDLssN$CRHC
C;RRRRkR#CHCCC38#0_oDFH4O_43ncN;DD
RRRRCk#RCHCC03#8F_Do_HOkHM#o8MC3DND;


CHM001$RAw_7w1 1R
H#RbRRFRs05RR
R RRRRR:HRMR#_08DHFoO=R:R''];R
RRRR1RH:RM#RR0D8_FOoH;R
SRRTR:kRF0#RR0D8_FOoH;R
SRR7R:MRHR0R#8F_Do;HO
RSRB:RRRRHMR8#0_oDFHROR2S;
RCR
M18RAw_7w1 1;NR
0H0sLCk0RM#$_NLDOL	_FFGRVAR1_w7w R11:FROlMbFCRM0H0#Rs;kC
NR
sHOE00COkRsCVOkMRRFV17A_w1w 1#RH
oLCHRM
bOsFC5##BR2
RCRLo
HMSHRRV'RBCMPC0MRN8RRB=4R''ER0CSM
RRRRH VRR'=R40'RERCMRR
SRRRRRVRHR=1RR''40MEC
RSSRRRRRRRRR<TR=4R''S;
SRRRRDRC#SC
SRRRRRRRRTRRRR<=7R;
RRRRRMRC8VRH;R
RRRRRCRM8H
V;RRRRCRM8H
V;RCRRMb8RsCFO#
#;CRM8RMVkO
;

=--=========================================================================
==-1-RAw_7wR )
=--=========================================================================
==
RRRRLDHs$NsRCHCCR;
RkRR#HCRC3CC#_08DHFoO4_4nNc3D
D;RRRRkR#CHCCC38#0_oDFHkO_Mo#HM3C8N;DD
C

M00H$AR1_w7w H)R#R
RRsbF0RR5
RRRRR R:MRHR0R#8F_DoRHO:'=R]
';RRRR):RRRRHMR8#0_oDFH
O;STRRRRR:FRk0R8#0_oDFH
O;S7RRRRR:HRMR#_08DHFoOS;
RRRBRH:RM#RR0D8_FOoHR;R2
RSR
8CMR_1A7 ww)
;RNs00H0LkC$R#MD_LN_O	LRFGF1VRAw_7wR ):FROlMbFCRM0H0#Rs;kC
NR
sHOE00COkRsCVOkMRRFV17A_w)w R
H#LHCoMb
RsCFO#B#5R),RRR2
RCRLo
HMSHRRVBR5'CCPMN0RMB8RR'=R4R'2m5)R)P'CCRM0NRM8)RR='24'RER0CSM
RRRRH VRR'=R40'RERCMRR
SRRRRRVRHR=)RR''40MEC
RSSRRRRRRRRR<TR=jR''S;
SRRRRDRC#SC
SRRRRRRRRTRRRR<=7R;
RRRRRRRRCRM8H
V;RRRRRMRC8VRH;R
RRMRC8VRH;R
RR8CMRFbsO#C#;M
C8VRRk;MO
-

-============================================================================-
-R_1A7 ww1-R
-============================================================================R

RDRRHNLssH$RC;CC
RRRRCk#RCHCC03#8F_Do_HO4c4n3DND;R
RR#RkCCRHC#C30D8_FOoH_#kMHCoM8D3ND
;
CHM001$RAw_7wR 1HR#
RFRbs50RRR
RRRR RH:RM#RR0D8_FOoHRR:=';]'
RRRRR1R:MRHR0R#8F_Do;HO
RSRT:RRR0FkR0R#8F_Do;HO
RSR7:RRRRHMR8#0_oDFH
O;SBRRRRR:HRMR#_08DHFoO2RR;R
SRM
C8AR1_w7w R1;
0N0skHL0#CR$LM_D	NO_GLFRRFV17A_w1w RO:RFFlbM0CMRRH#0Csk;

RNEsOHO0C0CksRMVkOVRFR_1A7 ww1#RH
oLCHRM
bOsFC5##BRR,1R2
RCRLo
HMSHRRVBR5'CCPMN0RMB8RR'=R4R'2m5)R1P'CCRM0NRM81RR='24'RER0CSM
RRRRH VRR'=R40'RERCMRR
SRRRRRVRHR=1RR''40MEC
RSSRRRRRRRRR<TR=4R''S;
SRRRRDRC#SC
SRRRRRRRRTRRRR<=7R;
RRRRRRRRCRM8H
V;RRRRRMRC8VRH;R
RRMRC8VRH;R
RR8CMRFbsO#C#;M
C8VRRk;MO
-

-============================================================================-
-R_1A7hwwR-
-============================================================================
R
RRHRDLssN$CRHC
C;RRRRkR#CHCCC38#0_oDFH4O_43ncN;DD
RRRRCk#RCHCC03#8F_Do_HOkHM#o8MC3DND;C

M00H$AR1_w7wh#RH
RRRb0FsR
5RSTRRRRR:FRk0R8#0_oDFH
O;S7RRRRR:HRMR#_08DHFoOS;
RRRBRH:RM#RR0D8_FOoHR;R2
RSR
8CMR_1A7hww;NR
0H0sLCk0RM#$_NLDOL	_FFGRVAR1_w7whRR:ObFlFMMC0#RHRk0sCR;

ONsECH0Os0kCkRVMFORVAR1_w7wh#RH
oLCHRM
bOsFC5##BR2
RCRLo
HMSHRRV'RBCMPC0MRN8RRB=jR''ER0CSM
SRRT<7=R;R
RRRRRCRM8H
V;RCRRMb8RsCFO#
#;CRM8RMVkO
;

=--=========================================================================
==-1-RAw_7w)h1R-
-============================================================================
R
RRHRDLssN$CRHC
C;RRRRkR#CHCCC38#0_oDFH4O_43ncN;DD
RRRRCk#RCHCC03#8F_Do_HOkHM#o8MC3DND;C

M00H$AR1_w7whR1)HR#
RFRbs50RRR
RRRR)RH:RM#RR0D8_FOoH;R
SRRTR:kRF0#RR0D8_FOoH;R
SRR7R:MRHR0R#8F_Do;HO
RSRB:RRRRHMR8#0_oDFHROR2S;
RCR
M18RAw_7w)h1;NR
0H0sLCk0RM#$_NLDOL	_FFGRVAR1_w7whR1):FROlMbFCRM0H0#Rs;kC
NR
sHOE00COkRsCVOkMRRFV17A_w1wh)#RH
oLCHRM
bOsFC5##BR2
RCRLo
HMSHRRV'RBCMPC0MRN8RRB=jR''ER0CSM
RRRRRRHV)RR='04'E
CMSRSRRRRRRRRT<'=Rj
';SRSRR#CDCS
SRRRRRRRRT=R<R
7;RRRRRCRRMH8RVR;
RCRRMH8RVR;
RMRC8sRbF#OC#C;
MR8RVOkM;



=--=========================================================================
==-1-RAw_7w1h1R-
-============================================================================
R
RRHRDLssN$CRHC
C;RRRRkR#CHCCC38#0_oDFH4O_43ncN;DD
RRRRCk#RCHCC03#8F_Do_HOkHM#o8MC3DND;S

CHM001$RAw_7w1h1R
H#SRRRb0FsR
5RSRRRRR1R:MRHR0R#8F_Do;HO
RSSRRTR:kRF0#RR0D8_FOoH;S
SRRR7RH:RM#RR0D8_FOoH;S
SRRRBRH:RM#RR0D8_FOoHR;R2
RSSRC
SM18RAw_7w1h1;SR
Ns00H0LkC$R#MD_LN_O	LRFGF1VRAw_7w1h1RO:RFFlbM0CMRRH#0Csk;R
S
sSNO0EHCkO0sVCRkRMOF1VRAw_7w1h1R
H#SoLCHSM
RFbsO#C#5
B2SRRRLHCoMS
SRVRHRCB'P0CMR8NMR=BRR''jRC0EMS
SRRRRRRHV1RR='04'E
CMSRSSRRRRRTRRRR<=';4'
SSSRCRRD
#CSRSSRRRRRTRRRR<=7S;
RRRRRCRRMH8RVS;
RRRRCRM8H
V;SRRRCRM8bOsFC;##
MSC8VRRk;MO

S
-=-==========================================================================-=
-AR1_w7wh
)R-=-==========================================================================
=
RRRRDsHLNRs$HCCC;R
RR#RkCCRHC#C30D8_FOoH_n44cD3NDR;
RkRR#HCRC3CC#_08DHFoOM_k#MHoCN83D
D;
0CMHR0$17A_w)whR
H#RbRRFRs05RR
R)RRRRR:HRMR#_08DHFoOS;
RRRTRF:RkR0R#_08DHFoOS;
RRR7RH:RM#RR0D8_FOoH;R
SRRBR:MRHR0R#8F_DoRHOR
2;S
RRCRM817A_w)wh;NR
0H0sLCk0RM#$_NLDOL	_FFGRVAR1_w7wh:)RRlOFbCFMMH0R#sR0k
C;Rs
NO0EHCkO0sVCRkRMOF1VRAw_7wRh)HL#
CMoH
sRbF#OC#R5B,RR)2R
RRoLCHSM
RVRHR'5BCMPC0MRN8RRB=jR''m2R))R5'CCPMN0RM)8RR'=R4R'2RC0EMR
SRRRRH)VRR'=R4E'0CSM
SRRRRRRRR<TR=jR''S;
SRRRCCD#
RSSRRRRRTRRRR<=7R;
RRRRRMRC8VRH;R
RRMRC8VRH;R
RR8CMRFbsO#C#;M
C8VRRk;MO
-

-============================================================================-
-R_1A7hww1-R
-============================================================================R

RDRRHNLssH$RC;CC
RRRRCk#RCHCC03#8F_Do_HO4c4n3DND;R
RR#RkCCRHC#C30D8_FOoH_#kMHCoM8D3ND
;

0CMHR0$17A_w1whR
H#RbRRFRs05RR
R1RRRRR:HRMR#_08DHFoOS;
RRRTRF:RkR0R#_08DHFoOS;
RRR7RH:RM#RR0D8_FOoH;R
SRRBR:MRHR0R#8F_DoRHOR
2;S
RRCRM817A_w1wh;NR
0H0sLCk0RM#$_NLDOL	_FFGRVAR1_w7wh:1RRlOFbCFMMH0R#sR0k
C;Rs
NO0EHCkO0sVCRkRMOF1VRAw_7wRh1HL#
CMoH
sRbF#OC#R5B,RR12R
RRoLCHSM
RVRHR'5BCMPC0MRN8RRB=jR''m2R)1R5'CCPMN0RM18RR'=R4R'2RC0EMR
SRRRRH1VRR'=R4E'0CSM
SRRRRRRRR<TR=4R''S;
SRRRCCD#
RSSRRRRRTRRRR<=7R;
RRRRRMRC8VRH;R
RRMRC8VRH;R
RR8CMRFbsO#C#;M
C8VRRk;MO
-

-============================================================================-
-R_1A7hww -R
-============================================================================R

RDRRHNLssH$RC;CC
RRRRCk#RCHCC03#8F_Do_HO4c4n3DND;R
RR#RkCCRHC#C30D8_FOoH_#kMHCoM8D3ND
;

0CMHR0$17A_w whR
H#RbRRFRs05RR
R RRRRR:HRMR#_08DHFoO=R:R''];R
SRRTR:kRF0#RR0D8_FOoH;R
SRR7R:MRHR0R#8F_Do;HO
RSRB:RRRRHMR8#0_oDFHROR2S;
RCR
M18RAw_7w;h R0
N0LsHkR0C#_$MLODN	F_LGVRFR_1A7hww RR:ObFlFMMC0#RHRk0sCR;

ONsECH0Os0kCkRVMFORVAR1_w7whH R#C
Lo
HMRFbsO#C#5
B2RLRRCMoH
RSRHBVR'CCPMN0RMB8RR'=RjR'R0MEC
RSRRHRRVRR =4R''C0EMS
SRRRRRRRRT=R<R
7;SRSRR8CMR;HV
RRRR8CMR;HV
RRRCRM8bOsFC;##
8CMRkRVM
O;
-
-============================================================================
R--17A_w wh1
)R-=-==========================================================================
=
RRRRDsHLNRs$HCCC;R
RR#RkCCRHC#C30D8_FOoH_n44cD3NDR;
RkRR#HCRC3CC#_08DHFoOM_k#MHoCN83D
D;
M
C0$H0R_1A7hww R1)HR#
RFRbs50RRR
RRRR RH:RM#RR0D8_FOoHRR:=';]'
RRRRR)R:MRHR0R#8F_Do;HO
RSRT:RRR0FkR0R#8F_Do;HO
RSR7:RRRRHMR8#0_oDFH
O;SBRRRRR:HRMR#_08DHFoO2RR;R
SRM
C8AR1_w7wh) 1;NR
0H0sLCk0RM#$_NLDOL	_FFGRVAR1_w7wh) 1RO:RFFlbM0CMRRH#0Csk;

RNEsOHO0C0CksRMVkOVRFR_1A7hww R1)HL#
CMoH
sRbF#OC#25B
RRRLHCoMR
SRRHVBP'CCRM0NRM8BRR='Rj'0MEC
RSRRVRHR= RR''4RC0EM
RRSRRRRRRRH)VRR'=R4E'0CSM
SRRRRRRRRTRRRR<=';j'
RSSRRRRCCD#
RSSRRRRRRRRR<TR=;R7
RRRRRRRCRM8H
V;RRRRRMRC8VRH;R
RRMRC8VRH;R
RR8CMRFbsO#C#;M
C8VRRk;MO
-

-============================================================================-
-R_1A7hww R11
=--=========================================================================
==
RRRRLDHs$NsRCHCCR;
RkRR#HCRC3CC#_08DHFoO4_4nNc3D
D;RRRRkR#CHCCC38#0_oDFHkO_Mo#HM3C8N;DD



CHM001$RAw_7w1h 1#RH
RRRb0FsR
5RRRRR :RRRRHMR8#0_oDFH:OR=]R''R;
R1RRRRR:HRMR#_08DHFoOS;
RRRTRF:RkR0R#_08DHFoOS;
RRR7RH:RM#RR0D8_FOoH;R
SRRBR:MRHR0R#8F_DoRHOR
2;S
RRCRM817A_w wh1R1;
0N0skHL0#CR$LM_D	NO_GLFRRFV17A_w wh1:1RRlOFbCFMMH0R#sR0k
C;Rs
NO0EHCkO0sVCRkRMOF1VRAw_7w1h 1#RH
oLCHRM
bOsFC5##BR2
RCRLo
HMSHRRV'RBCMPC0MRN8RRB=jR''ER0CSM
RRRRH VRR'=R40'RERCMRR
SRRRRRVRHR=1RR''40MEC
RSSRRRRRRRRR<TR=4R''S;
SRRRRDRC#SC
SRRRRRRRRTRRRR<=7R;
RRRRRMRC8VRH;R
RRRRRCRM8H
V;RRRRCRM8H
V;RCRRMb8RsCFO#
#;CRM8RMVkO
;

=--=========================================================================
==-1-RAw_7w)h R-
-============================================================================
R
RRHRDLssN$CRHC
C;RRRRkR#CHCCC38#0_oDFH4O_43ncN;DD
RRRRCk#RCHCC03#8F_Do_HOkHM#o8MC3DND;


CHM001$RAw_7w)h R
H#RbRRFRs05RR
R RRRRR:HRMR#_08DHFoO=R:R''];R
RRRR)RH:RM#RR0D8_FOoH;R
SRRTR:kRF0#RR0D8_FOoH;R
SRR7R:MRHR0R#8F_Do;HO
RSRB:RRRRHMR8#0_oDFHROR2S;
RCR
M18RAw_7w)h ;NR
0H0sLCk0RM#$_NLDOL	_FFGRVAR1_w7whR ):FROlMbFCRM0H0#Rs;kC
NR
sHOE00COkRsCVOkMRRFV17A_w wh)#RH
oLCHRM
bOsFC5##BRR,)
R2RLRRCMoH
RSRH5VRBP'CCRM0NRM8BRR='2j'RRm)5C)'P0CMR8NMR=)RR''420RRE
CMSRRRRRHV RR='R4'0MECRSR
RRRRRHRRVRR)=4R''C0EMS
SRRRRRRRRRRRT<'=Rj
';SRSRRCRRD
#CSRSRRRRRRRRRT=R<R
7;RRRRRRRRR8CMR;HV
RRRRCRRMH8RVR;
RCRRMH8RVR;
RMRC8sRbF#OC#C;
MR8RVOkM;


-=-==========================================================================-=
-AR1_w7whR 1
=--=========================================================================
==
RRRRLDHs$NsRCHCCR;
RkRR#HCRC3CC#_08DHFoO4_4nNc3D
D;RRRRkR#CHCCC38#0_oDFHkO_Mo#HM3C8N;DD
M
C0$H0R_1A7hww H1R#R
RRsbF0RR5
RRRRR R:MRHR0R#8F_DoRHO:'=R]
';RRRR1:RRRRHMR8#0_oDFH
O;STRRRRR:FRk0R8#0_oDFH
O;S7RRRRR:HRMR#_08DHFoOS;
RRRBRH:RM#RR0D8_FOoHR;R2
RSR
8CMR_1A7hww R1;
0N0skHL0#CR$LM_D	NO_GLFRRFV17A_w wh1RR:ObFlFMMC0#RHRk0sCR;

ONsECH0Os0kCkRVMFORVAR1_w7whR 1HL#
CMoH
sRbF#OC#R5B,2R1
RRRLHCoMR
SRRHV5CB'P0CMR8NMR=BRR''j2)RmR'51CMPC0MRN8RR1=4R''R2R0MEC
RSRRVRHR= RR''4RC0EM
RRSRRRRRRRH1VRR'=R4E'0CSM
SRRRRRRRRTRRRR<=';4'
RSSRRRRCCD#
RSSRRRRRRRRR<TR=;R7
RRRRRRRRMRC8VRH;R
RRRRRCRM8H
V;RRRRCRM8H
V;RCRRMb8RsCFO#
#;CRM8RMVkO
;
-----------------------------------------------------------------------------
-----R-------------------------------------------------------------------------
-----R-------------------------AR1aORHCjRcR-------------------------------------------
R------------------------------------------------------------------------------
-------------------------------------------------------------------------------
-------------------------------------------------------------------------------
-------------------------------------------------------------------------------
-------------------------------------------------------------------------------
-------------------------------------------------------------------------------
C

M00H$AR1_v)q.G6n4HnR#R

RMoCCOsHR
5RRRRRRRRRRQRRh_QajRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QacRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ6a_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QaURR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQga_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QaBRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ7a_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_ :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
"RRRRRRRRRRRRR2
R;RRRRRRRRRFRbsR05
RRRRRRRRRRRRRRRRq)7a:qRR0FkR8#0_oDFHPO_CFO0s45R68RRF0IMF2RjRR;
RRRRRRRRRRRRR)RRBRpiRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRR)RRB piRH:RM#RR0D8_FOoHRR:=';]'
RRRRRRRRRRRRRRRRR) R:RRRRHMR8#0_oDFH:OR=]R''R;
RRRRRRRRRRRRR)RRq)77RH:RM#RR0D8_FOoH_OPC05FsRR(R8MFI0jFR2
R;RRRRRRRRRRRRRRRRWiBpRRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRRWiBp RR:HRMR#_08DHFoO=R:R''];R
RRRRRRRRRRRRRR RWRRRR:MRHR0R#8F_DoRHO:'=R]
';RRRRRRRRRRRRRRRRW7q7)RR:HRMR#_08DHFoOC_POs0F5RR(RI8FMR0Fj;2R
RRRRRRRRRRRRRRRR1vqi:RRRRHMR8#0_oDFHPO_CFO0s45R68RRF0IMF2RjRR;
RRRRRRRRRRRRRWRR7qqaRH:RM#RR0D8_FOoH_OPC05FsRR46RI8FMR0FjR2
RRRRRRRRRRRRR;R2

RRRCR
M18RAq_)vn.6G;4n
s
NO0EHCkO0s1CRAq_)vn.6G_4nq])BRRFV1)A_q6v.nnG4R
H#LHCoMCR
M18RAq_)vn.6G_4nq])B;RRR-R--1)A_q6v.nnG4
-

-------------------------------------S-
-R--1)A_q6v.nnG4h-)
-------------------------------------D-
HNLssQ$R ;  
Ck#R Q  a317m_pt_QB4c4n3DND;#
kC RQ 1 3ap7_mBtQ_1zhQ th7D3NDk;
#QCR 3  #_08DHFoOs_NH30EN;DD
 z1R Q  k3MlHCsO0_#8p3qp
;
CHM001$RAq_)vn.6Gh4n)#RH
R
RoCCMsRHO5RR
RRRRRRRRRhRQQja_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QadRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQca_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQUa_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QaARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQBa_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QawRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"RR
RRRRRRRRR2RRRR;
RRRRRRRRRsbF0
5RRRRRRRRRRRRRRRRR)a7qqRR:FRk0#_08DHFoOC_POs0F56R4RFR8IFM0RRj2;R
RRRRRRRRRRRRRRBR)pRih:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRBR)pRi :MRHR0R#8F_DoRHO:'=R]
';RRRRRRRRRRRRRRRR)R RRRR:HRMR#_08DHFoO=R:R''];R
RRRRRRRRRRRRRRqR)7R7):MRHR0R#8F_Do_HOP0COFRs5(8RRF0IMF2RjRR;
RRRRRRRRRRRRRWRRBRpiRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRRWRRB piRH:RM#RR0D8_FOoHRR:=';]'
RRRRRRRRRRRRRRRRRW R:RRRRHMR8#0_oDFH:OR=]R''R;
RRRRRRRRRRRRRWRRq)77RH:RM#RR0D8_FOoH_OPC05FsRR(R8MFI0jFR2
R;RRRRRRRRRRRRRRRRviq1RRR:HRMR#_08DHFoOC_POs0F56R4RFR8IFM0RRj2;R
RRRRRRRRRRRRRR7RWqRaq:MRHR0R#8F_Do_HOP0COFRs54R6R8MFI0jFR2R
RRRRRRRRRRRRRR
2;RRR
RM
C8AR1_v)q.G6n4)nh;N

sHOE00COkRsC1)A_q6v.nnG4hq)_)RB]F1VRAq_)vn.6Gh4n)#RH
oLCH
MRCRM81)A_q6v.nnG4hq)_);B]R-RR-1-RAq_)vn.6Gh4n)


-------------------------------------
--S---R_1A).qv64nGn
hW-------------------------------------
--DsHLNRs$Q   ;#
kC RQ 1 3ap7_mBtQ_n44cD3NDk;
#QCR 3  1_a7pQmtBh_z1hQt N73D
D;kR#CQ   38#0_oDFHNO_sEH03DND;1
z  RQ M 3kslCH#O_0q83p
p;
0CMHR0$1)A_q6v.nnG4hHWR#R

RMoCCOsHR
5RRRRRRRRRRQRRh_QajRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QacRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ6a_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QaURR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQga_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QaBRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ7a_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_ :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
"RRRRRRRRRRRRR2
R;RRRRRRRRRFRbsR05
RRRRRRRRRRRRRRRRq)7a:qRR0FkR8#0_oDFHPO_CFO0s45R68RRF0IMF2RjRR;
RRRRRRRRRRRRR)RRBRpiRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRR)RRB piRH:RM#RR0D8_FOoHRR:=';]'
RRRRRRRRRRRRRRRRR) R:RRRRHMR8#0_oDFH:OR=]R''R;
RRRRRRRRRRRRR)RRq)77RH:RM#RR0D8_FOoH_OPC05FsRR(R8MFI0jFR2
R;RRRRRRRRRRRRRRRRWiBphRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRRWiBp RR:HRMR#_08DHFoO=R:R''];R
RRRRRRRRRRRRRR RWRRRR:MRHR0R#8F_DoRHO:'=R]
';RRRRRRRRRRRRRRRRW7q7)RR:HRMR#_08DHFoOC_POs0F5RR(RI8FMR0Fj;2R
RRRRRRRRRRRRRRRR1vqi:RRRRHMR8#0_oDFHPO_CFO0s45R68RRF0IMF2RjRR;
RRRRRRRRRRRRRWRR7qqaRH:RM#RR0D8_FOoH_OPC05FsRR46RI8FMR0FjR2
RRRRRRRRRRRRR;R2

RRRCR
M18RAq_)vn.6Xh4nW
;
NEsOHO0C0CksR_1A).qv64nGn_hWq])BRRFV1)A_q6v.nnG4hHWR#C
LoRHM
8CMR_1A).qv64nGn_hWq])B;RRR-R--1)A_q6v.nnG4h
W

-
---------------------------------------
S-1-RAq_)vn.6Gh4n)
hW-------------------------------------
--DsHLNRs$Q   ;#
kC RQ 1 3ap7_mBtQ_n44cD3NDk;
#QCR 3  1_a7pQmtBh_z1hQt N73D
D;kR#CQ   38#0_oDFHNO_sEH03DND;1
z  RQ M 3kslCH#O_0q83p
p;
0CMHR0$1)A_q6v.nnG4hW)hR
H#
oRRCsMCH5ORRR
RRRRRRRRRRQQhaR_j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QanRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ(a_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QaqRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQAa_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQwa_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jjRR
RRRRRRRRRRRR2;R
RRRRRRRRRb0Fs5RR
RRRRRRRRRRRRR)RR7qqaRF:Rk#0R0D8_FOoH_OPC05FsRR46RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRp)Bi:hRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRp)Bi: RRRHMR8#0_oDFH:OR=]R''R;
RRRRRRRRRRRRR)RR RRRRH:RM#RR0D8_FOoHRR:=';]'
RRRRRRRRRRRRRRRR7)q7:)RRRHMR8#0_oDFHPO_CFO0s(5RRFR8IFM0RRj2;R
RRRRRRRRRRRRRRBRWpRih:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRBRWpRi :MRHR0R#8F_DoRHO:'=R]
';RRRRRRRRRRRRRRRRWR RRRR:HRMR#_08DHFoO=R:R''];R
RRRRRRRRRRRRRRqRW7R7):MRHR0R#8F_Do_HOP0COFRs5(8RRF0IMF2RjRR;
RRRRRRRRRRRRRvRRqR1iRH:RM#RR0D8_FOoH_OPC05FsRR46RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRqW7a:qRRRHMR8#0_oDFHPO_CFO0s45R68RRF0IMF2Rj
RRRRRRRRRRRRRRR2R;
RR
R
8CMR_1A).qv64nGnhh)W
;
NEsOHO0C0CksR_1A).qv64nGnhh)W)_qBF]RVAR1_v)q.G6n4)nhhHWR#C
LoRHM
8CMR_1A).qv64nGnhh)W)_qBR];R-R--AR1_v)q.G6n4)nhh
W

---------------------------------------
-S--AR1_v)q6G4.U-
--------------------------------------H
DLssN$ RQ 
 ;kR#CQ   371a_tpmQ4B_43ncN;DD
Ck#R Q  a317m_pt_QBzQh1t7h 3DND;#
kC RQ # 30D8_FOoH_HNs0NE3D
D;zR1 Q   3lMkCOsH_8#03pqp;C

M00H$AR1_v)q6G4.U#RH
R
RoCCMsRHO5RR
RRRRRRRRRhRQQja_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QadRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQca_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQUa_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QaARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQBa_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QawRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"RR
RRRRRRRRR2RRRR;
RRRRRRRRRsbF0
5RRRRRRRRRRRRRRRRR)a7qqRR:FRk0#_08DHFoOC_POs0F5RR(RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRp)Bi:RRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRp)Bi: RRRHMR8#0_oDFH:OR=]R''R;
RRRRRRRRRRRRR)RR RRRRH:RM#RR0D8_FOoHRR:=';]'
RRRRRRRRRRRRRRRR7)q7:)RRRHMR8#0_oDFHPO_CFO0sU5RRFR8IFM0RRj2;R
RRRRRRRRRRRRRRBRWpRiR:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRBRWpRi :MRHR0R#8F_DoRHO:'=R]
';RRRRRRRRRRRRRRRRWR RRRR:HRMR#_08DHFoO=R:R''];R
RRRRRRRRRRRRRRqRW7R7):MRHR0R#8F_Do_HOP0COFRs5U8RRF0IMF2RjRR;
RRRRRRRRRRRRRWRR7qqaRH:RM#RR0D8_FOoH_OPC05FsRR(R8MFI0jFR2R
RRRRRRRRRRRRRR
2;RRR
RM
C8AR1_v)q6G4.U
;
NEsOHO0C0CksR_1A)6qv4U.G_Bq)]VRFR_1A)6qv4U.GR
H#LHCoMCR
M18RAq_)v.64GqU_);B]R-RR-1-RAq_)v.64G
U

-
---------------------------------------
S-1-RAq_)v.64G)Uh
---------------------------------------
LDHs$NsR Q  k;
#QCR 3  1_a7pQmtB4_4nNc3D
D;kR#CQ   371a_tpmQzB_ht1Qh3 7N;DD
Ck#R Q  03#8F_Do_HON0sHED3NDz;
1Q R 3  MCkls_HO#308q;pp
M
C0$H0R_1A)6qv4U.GhH)R#R

RMoCCOsHR
5RRRRRRRRRRQRRh_QajRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QacRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ6a_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QaURR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQga_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QaBRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ7a_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_ :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
"RRRRRRRRRRRRR2
R;RRRRRRRRRFRbsR05
RRRRRRRRRRRRRRRRq)7a:qRR0FkR8#0_oDFHPO_CFO0s(5RRFR8IFM0RRj2;R
RRRRRRRRRRRRRRBR)pRih:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRBR)pRi :MRHR0R#8F_DoRHO:'=R]
';RRRRRRRRRRRRRRRR)R RRRR:HRMR#_08DHFoO=R:R''];R
RRRRRRRRRRRRRRqR)7R7):MRHR0R#8F_Do_HOP0COFRs5U8RRF0IMF2RjRR;
RRRRRRRRRRRRRWRRBRpiRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRRWRRB piRH:RM#RR0D8_FOoHRR:=';]'
RRRRRRRRRRRRRRRRRW R:RRRRHMR8#0_oDFH:OR=]R''R;
RRRRRRRRRRRRRWRRq)77RH:RM#RR0D8_FOoH_OPC05FsRRUR8MFI0jFR2
R;RRRRRRRRRRRRRRRRWa7qqRR:HRMR#_08DHFoOC_POs0F5RR(RI8FMR0FjR2
RRRRRRRRRRRRR;R2

RRRCR
M18RAq_)v.64G)Uh;N

sHOE00COkRsC1)A_q4v6.hGU))_qBF]RVAR1_v)q6G4.URh)HL#
CMoHRM
C8AR1_v)q6G4.U_h)q])B;RRR-R--1)A_q4v6.hGU)



---------------------------------------
-S--AR1_v)q6G4.U
hW-------------------------------------
--DsHLNRs$Q   ;#
kC RQ 1 3ap7_mBtQ_n44cD3NDk;
#QCR 3  1_a7pQmtBh_z1hQt N73D
D;kR#CQ   38#0_oDFHNO_sEH03DND;1
z  RQ M 3kslCH#O_0q83p
p;
0CMHR0$1)A_q4v6.hGUW#RH
R
RoCCMsRHO5RR
RRRRRRRRRhRQQja_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QadRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQca_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQUa_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QaARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQBa_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QawRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"RR
RRRRRRRRR2RRRR;
RRRRRRRRRsbF0
5RRRRRRRRRRRRRRRRR)a7qqRR:FRk0#_08DHFoOC_POs0F5RR(RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRp)Bi:RRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRp)Bi: RRRHMR8#0_oDFH:OR=]R''R;
RRRRRRRRRRRRR)RR RRRRH:RM#RR0D8_FOoHRR:=';]'
RRRRRRRRRRRRRRRR7)q7:)RRRHMR8#0_oDFHPO_CFO0sU5RRFR8IFM0RRj2;R
RRRRRRRRRRRRRRBRWpRih:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRBRWpRi :MRHR0R#8F_DoRHO:'=R]
';RRRRRRRRRRRRRRRRWR RRRR:HRMR#_08DHFoO=R:R''];R
RRRRRRRRRRRRRRqRW7R7):MRHR0R#8F_Do_HOP0COFRs5U8RRF0IMF2RjRR;
RRRRRRRRRRRRRWRR7qqaRH:RM#RR0D8_FOoH_OPC05FsRR(R8MFI0jFR2R
RRRRRRRRRRRRRR
2;RRR
RM
C8AR1_v)q6G4.U;hW
s
NO0EHCkO0s1CRAq_)v.64GWUh_Bq)]VRFR_1A)6qv4U.GhHWR#C
LoRHM
8CMR_1A)6qv4U.GhqW_);B]R-RR-1-RAq_)v.64GWUh
-

-------------------------------------S-
-R--1)A_q4v6.hGU)
hW-------------------------------------
--DsHLNRs$Q   ;#
kC RQ 1 3ap7_mBtQ_n44cD3NDk;
#QCR 3  1_a7pQmtBh_z1hQt N73D
D;kR#CQ   38#0_oDFHNO_sEH03DND;1
z  RQ M 3kslCH#O_0q83p
p;
0CMHR0$1)A_q4v6.hGU)RhWH
#
RCRoMHCsORR5
RRRRRRRRRRRQahQ_:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQna_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QagRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQqa_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ a_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjRj"
RRRRRRRRRRRR;2R
RRRRRRRRbRRF5s0RR
RRRRRRRRRRRRRR7R)qRaq:kRF00R#8F_Do_HOP0COFRs5(8RRF0IMF2RjRR;
RRRRRRRRRRRRR)RRBhpiRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRR)RRB piRH:RM#RR0D8_FOoHRR:=';]'
RRRRRRRRRRRRRRRRR) R:RRRRHMR8#0_oDFH:OR=]R''R;
RRRRRRRRRRRRR)RRq)77RH:RM#RR0D8_FOoH_OPC05FsRRUR8MFI0jFR2
R;RRRRRRRRRRRRRRRRWiBphRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRRWiBp RR:HRMR#_08DHFoO=R:R''];R
RRRRRRRRRRRRRR RWRRRR:MRHR0R#8F_DoRHO:'=R]
';RRRRRRRRRRRRRRRRW7q7)RR:HRMR#_08DHFoOC_POs0F5RRURI8FMR0Fj;2R
RRRRRRRRRRRRRRRRqW7a:qRRRHMR8#0_oDFHPO_CFO0s(5RRFR8IFM0R
j2RRRRRRRRRRRRR2RR;R
R

RRCRM81)A_q4v6.hGU);hW
s
NO0EHCkO0s1CRAq_)v.64G)UhhqW_)RB]F1VRAq_)v.64G)UhhHWR#C
LoRHM
8CMR_1A)6qv4U.GhW)h_Bq)]R;RR---R_1A)6qv4U.GhW)h
-

-------------------------------------S-
-R--1)A_qjv4.ccG
---------------------------------------
LDHs$NsR Q  k;
#QCR 3  1_a7pQmtB4_4nNc3D
D;kR#CQ   371a_tpmQzB_ht1Qh3 7N;DD
Ck#R Q  03#8F_Do_HON0sHED3NDz;
1Q R 3  MCkls_HO#308q;pp
M
C0$H0R_1A)4qvjG.cc#RH
R
RoCCMsRHO5RR
RRRRRRRRRhRQQja_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QadRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQca_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQUa_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QaARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQBa_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QawRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"RR
RRRRRRRRR2RRRR;
RRRRRRRRRsbF0
5RRRRRRRRRRRRRRRRR)a7qqRR:FRk0#_08DHFoOC_POs0F5RRdRI8FMR0Fj;2R
RRRRRRRRRRRRRRRRp)Bi:RRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRp)Bi: RRRHMR8#0_oDFH:OR=]R''R;
RRRRRRRRRRRRR)RR RRRRH:RM#RR0D8_FOoHRR:=';]'
RRRRRRRRRRRRRRRR7)q7:)RRRHMR8#0_oDFHPO_CFO0sg5RRFR8IFM0RRj2;R
RRRRRRRRRRRRRRBRWpRiR:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRBRWpRi :MRHR0R#8F_DoRHO:'=R]
';RRRRRRRRRRRRRRRRWR RRRR:HRMR#_08DHFoO=R:R''];R
RRRRRRRRRRRRRRqRW7R7):MRHR0R#8F_Do_HOP0COFRs5g8RRF0IMF2RjRR;
RRRRRRRRRRRRRWRR7qqaRH:RM#RR0D8_FOoH_OPC05FsRRdR8MFI0jFR2R
RRRRRRRRRRRRRR
2;RRR
RM
C8AR1_v)q4cj.G
c;
ONsECH0Os0kCAR1_v)q4cj.Gqc_)RB]F1VRAq_)v.4jcRGcHL#
CMoHRM
C8AR1_v)q4cj.Gqc_);B]R-RR-1-RAq_)v.4jc
Gc
-

-------------------------------------S-
-R--1)A_qjv4.ccGh-)
-------------------------------------D-
HNLssQ$R ;  
Ck#R Q  a317m_pt_QB4c4n3DND;#
kC RQ 1 3ap7_mBtQ_1zhQ th7D3NDk;
#QCR 3  #_08DHFoOs_NH30EN;DD
 z1R Q  k3MlHCsO0_#8p3qp
;
CHM001$RAq_)v.4jchGc)#RH
R
RoCCMsRHO5RR
RRRRRRRRRhRQQja_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QadRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQca_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQUa_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QaARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQBa_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QawRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"RR
RRRRRRRRR2RRRR;
RRRRRRRRRsbF0
5RRRRRRRRRRRRRRRRR)a7qqRR:FRk0#_08DHFoOC_POs0F5RRdRI8FMR0Fj;2R
RRRRRRRRRRRRRRRRp)Bi:hRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRp)Bi: RRRHMR8#0_oDFH:OR=]R''R;
RRRRRRRRRRRRR)RR RRRRH:RM#RR0D8_FOoHRR:=';]'
RRRRRRRRRRRRRRRR7)q7:)RRRHMR8#0_oDFHPO_CFO0sg5RRFR8IFM0RRj2;R
RRRRRRRRRRRRRRBRWpRiR:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRBRWpRi :MRHR0R#8F_DoRHO:'=R]
';RRRRRRRRRRRRRRRRWR RRRR:HRMR#_08DHFoO=R:R''];R
RRRRRRRRRRRRRRqRW7R7):MRHR0R#8F_Do_HOP0COFRs5g8RRF0IMF2RjRR;
RRRRRRRRRRRRRWRR7qqaRH:RM#RR0D8_FOoH_OPC05FsRRdR8MFI0jFR2R
RRRRRRRRRRRRRR
2;RRR
RM
C8AR1_v)q4cj.G)ch;N

sHOE00COkRsC1)A_qjv4.ccGhq)_)RB]F1VRAq_)v.4jchGc)#RH
oLCH
MRCRM81)A_qjv4.ccGhq)_);B]R-RR-1-RAq_)v.4jchGc)


-------------------------------------
--S---R_1A)4qvjG.cc
hW-------------------------------------
--DsHLNRs$Q   ;#
kC RQ 1 3ap7_mBtQ_n44cD3NDk;
#QCR 3  1_a7pQmtBh_z1hQt N73D
D;kR#CQ   38#0_oDFHNO_sEH03DND;1
z  RQ M 3kslCH#O_0q83p
p;
0CMHR0$1)A_qjv4.ccGhHWR#R

RMoCCOsHR
5RRRRRRRRRRQRRh_QajRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QacRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ6a_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QaURR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQga_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QaBRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ7a_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_ :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
"RRRRRRRRRRRRR2
R;RRRRRRRRRFRbsR05
RRRRRRRRRRRRRRRRq)7a:qRR0FkR8#0_oDFHPO_CFO0sd5RRFR8IFM0RRj2;R
RRRRRRRRRRRRRRBR)pRiR:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRBR)pRi :MRHR0R#8F_DoRHO:'=R]
';RRRRRRRRRRRRRRRR)R RRRR:HRMR#_08DHFoO=R:R''];R
RRRRRRRRRRRRRRqR)7R7):MRHR0R#8F_Do_HOP0COFRs5g8RRF0IMF2RjRR;
RRRRRRRRRRRRRWRRBhpiRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRRWRRB piRH:RM#RR0D8_FOoHRR:=';]'
RRRRRRRRRRRRRRRRRW R:RRRRHMR8#0_oDFH:OR=]R''R;
RRRRRRRRRRRRRWRRq)77RH:RM#RR0D8_FOoH_OPC05FsRRgR8MFI0jFR2
R;RRRRRRRRRRRRRRRRWa7qqRR:HRMR#_08DHFoOC_POs0F5RRdRI8FMR0FjR2
RRRRRRRRRRRRR;R2

RRRCR
M18RAq_)v.4jchGcW
;
NEsOHO0C0CksR_1A)4qvjG.cc_hWq])BRRFV1)A_qjv4.ccGhHWR#C
LoRHM
8CMR_1A)4qvjG.cc_hWq])B;RRR-R--1)A_qjv4.ccGh
W

---------------------------------------
-S--AR1_v)q4cj.G)chh-W
-------------------------------------D-
HNLssQ$R ;  
Ck#R Q  a317m_pt_QB4c4n3DND;#
kC RQ 1 3ap7_mBtQ_1zhQ th7D3NDk;
#QCR 3  #_08DHFoOs_NH30EN;DD
 z1R Q  k3MlHCsO0_#8p3qp
;
CHM001$RAq_)v.4jchGc)RhWH
#
RCRoMHCsORR5
RRRRRRRRRRRQahQ_:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQna_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QagRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQqa_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ a_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjRj"
RRRRRRRRRRRR;2R
RRRRRRRRbRRF5s0RR
RRRRRRRRRRRRRR7R)qRaq:kRF00R#8F_Do_HOP0COFRs5d8RRF0IMF2RjRR;
RRRRRRRRRRRRR)RRBhpiRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRR)RRB piRH:RM#RR0D8_FOoHRR:=';]'
RRRRRRRRRRRRRRRRR) R:RRRRHMR8#0_oDFH:OR=]R''R;
RRRRRRRRRRRRR)RRq)77RH:RM#RR0D8_FOoH_OPC05FsRRgR8MFI0jFR2
R;RRRRRRRRRRRRRRRRWiBphRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRRWiBp RR:HRMR#_08DHFoO=R:R''];R
RRRRRRRRRRRRRR RWRRRR:MRHR0R#8F_DoRHO:'=R]
';RRRRRRRRRRRRRRRRW7q7)RR:HRMR#_08DHFoOC_POs0F5RRgRI8FMR0Fj;2R
RRRRRRRRRRRRRRRRqW7a:qRRRHMR8#0_oDFHPO_CFO0sd5RRFR8IFM0R
j2RRRRRRRRRRRRR2RR;R
R

RRCRM81)A_qjv4.ccGhW)h;N

sHOE00COkRsC1)A_qjv4.ccGhW)h_Bq)]VRFR_1A)4qvjG.cchh)W#RH
oLCH
MRCRM81)A_qjv4.ccGhW)h_Bq)]R;RR---R_1A)4qvjG.cchh)W


-------------------------------------
--S---R_1A).qvjGcU.-
--------------------------------------H
DLssN$ RQ 
 ;kR#CQ   371a_tpmQ4B_43ncN;DD
Ck#R Q  a317m_pt_QBzQh1t7h 3DND;#
kC RQ # 30D8_FOoH_HNs0NE3D
D;zR1 Q   3lMkCOsH_8#03pqp;C

M00H$AR1_v)q.UjcGH.R#R

RMoCCOsHR
5RRRRRRRRRRQRRh_QajRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QacRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ6a_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QaURR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQga_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QaBRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ7a_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_ :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
"RRRRRRRRRRRRR2
R;RRRRRRRRRFRbsR05
RRRRRRRRRRRRRRRRq)7a:qRR0FkR8#0_oDFHPO_CFO0s45RRFR8IFM0RRj2;R
RRRRRRRRRRRRRRBR)pRiR:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRBR)pRi :MRHR0R#8F_DoRHO:'=R]
';RRRRRRRRRRRRRRRR)R RRRR:HRMR#_08DHFoO=R:R''];R
RRRRRRRRRRRRRRqR)7R7):MRHR0R#8F_Do_HOP0COFRs54RjR8MFI0jFR2
R;RRRRRRRRRRRRRRRRWiBpRRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRRWiBp RR:HRMR#_08DHFoO=R:R''];R
RRRRRRRRRRRRRR RWRRRR:MRHR0R#8F_DoRHO:'=R]
';RRRRRRRRRRRRRRRRW7q7)RR:HRMR#_08DHFoOC_POs0F5jR4RFR8IFM0RRj2;R
RRRRRRRRRRRRRR7RWqRaq:MRHR0R#8F_Do_HOP0COFRs548RRF0IMF2Rj
RRRRRRRRRRRRRRR2R;
RR
R
8CMR_1A).qvjGcU.
;
NEsOHO0C0CksR_1A).qvjGcU.)_qBF]RVAR1_v)q.UjcGH.R#C
LoRHM
8CMR_1A).qvjGcU.)_qBR];R-R--AR1_v)q.UjcG
.

---------------------------------------
-S--AR1_v)q.UjcG).h
---------------------------------------
LDHs$NsR Q  k;
#QCR 3  1_a7pQmtB4_4nNc3D
D;kR#CQ   371a_tpmQzB_ht1Qh3 7N;DD
Ck#R Q  03#8F_Do_HON0sHED3NDz;
1Q R 3  MCkls_HO#308q;pp
M
C0$H0R_1A).qvjGcU.Rh)H
#
RCRoMHCsORR5
RRRRRRRRRRRQahQ_:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQna_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QagRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQqa_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ a_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjRj"
RRRRRRRRRRRR;2R
RRRRRRRRbRRF5s0RR
RRRRRRRRRRRRRR7R)qRaq:kRF00R#8F_Do_HOP0COFRs548RRF0IMF2RjRR;
RRRRRRRRRRRRR)RRBhpiRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRR)RRB piRH:RM#RR0D8_FOoHRR:=';]'
RRRRRRRRRRRRRRRRR) R:RRRRHMR8#0_oDFH:OR=]R''R;
RRRRRRRRRRRRR)RRq)77RH:RM#RR0D8_FOoH_OPC05FsRR4jRI8FMR0Fj;2R
RRRRRRRRRRRRRRRRpWBi:RRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRpWBi: RRRHMR8#0_oDFH:OR=]R''R;
RRRRRRRRRRRRRWRR RRRRH:RM#RR0D8_FOoHRR:=';]'
RRRRRRRRRRRRRRRR7Wq7:)RRRHMR8#0_oDFHPO_CFO0s45Rj8RRF0IMF2RjRR;
RRRRRRRRRRRRRWRR7qqaRH:RM#RR0D8_FOoH_OPC05FsRR4R8MFI0jFR2R
RRRRRRRRRRRRRR
2;RRR
RM
C8AR1_v)q.UjcG).h;N

sHOE00COkRsC1)A_qjv.c.UGhq)_)RB]F1VRAq_)vc.jUhG.)#RH
oLCH
MRCRM81)A_qjv.c.UGhq)_);B]R-RR-1-RAq_)vc.jUhG.)


-------------------------------------
--S---R_1A).qvjGcU.
hW-------------------------------------
--DsHLNRs$Q   ;#
kC RQ 1 3ap7_mBtQ_n44cD3NDk;
#QCR 3  1_a7pQmtBh_z1hQt N73D
D;kR#CQ   38#0_oDFHNO_sEH03DND;1
z  RQ M 3kslCH#O_0q83p
p;
0CMHR0$1)A_qjv.c.UGhHWR#R

RMoCCOsHR
5RRRRRRRRRRQRRh_QajRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QacRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ6a_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QaURR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQga_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QaBRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ7a_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_ :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
"RRRRRRRRRRRRR2
R;RRRRRRRRRFRbsR05
RRRRRRRRRRRRRRRRq)7a:qRR0FkR8#0_oDFHPO_CFO0s45RRFR8IFM0RRj2;R
RRRRRRRRRRRRRRBR)pRiR:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRBR)pRi :MRHR0R#8F_DoRHO:'=R]
';RRRRRRRRRRRRRRRR)R RRRR:HRMR#_08DHFoO=R:R''];R
RRRRRRRRRRRRRRqR)7R7):MRHR0R#8F_Do_HOP0COFRs54RjR8MFI0jFR2
R;RRRRRRRRRRRRRRRRWiBphRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRRWiBp RR:HRMR#_08DHFoO=R:R''];R
RRRRRRRRRRRRRR RWRRRR:MRHR0R#8F_DoRHO:'=R]
';RRRRRRRRRRRRRRRRW7q7)RR:HRMR#_08DHFoOC_POs0F5jR4RFR8IFM0RRj2;R
RRRRRRRRRRRRRR7RWqRaq:MRHR0R#8F_Do_HOP0COFRs548RRF0IMF2Rj
RRRRRRRRRRRRRRR2R;
RR
R
8CMR_1A).qvjGcU.;hW
s
NO0EHCkO0s1CRAq_)vc.jUhG.W)_qBF]RVAR1_v)q.UjcGW.hR
H#LHCoMCR
M18RAq_)vc.jUhG.W)_qBR];R-R--AR1_v)q.UjcGW.h
-

-------------------------------------S-
-R--1)A_qjv.c.UGhW)h
---------------------------------------
LDHs$NsR Q  k;
#QCR 3  1_a7pQmtB4_4nNc3D
D;kR#CQ   371a_tpmQzB_ht1Qh3 7N;DD
Ck#R Q  03#8F_Do_HON0sHED3NDz;
1Q R 3  MCkls_HO#308q;pp
M
C0$H0R_1A).qvjGcU.hh)W#RH
R
RoCCMsRHO5RR
RRRRRRRRRhRQQja_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QadRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQca_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQUa_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QaARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQBa_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QawRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"RR
RRRRRRRRR2RRRR;
RRRRRRRRRsbF0
5RRRRRRRRRRRRRRRRR)a7qqRR:FRk0#_08DHFoOC_POs0F5RR4RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRp)Bi:hRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRp)Bi: RRRHMR8#0_oDFH:OR=]R''R;
RRRRRRRRRRRRR)RR RRRRH:RM#RR0D8_FOoHRR:=';]'
RRRRRRRRRRRRRRRR7)q7:)RRRHMR8#0_oDFHPO_CFO0s45Rj8RRF0IMF2RjRR;
RRRRRRRRRRRRRWRRBhpiRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRRWRRB piRH:RM#RR0D8_FOoHRR:=';]'
RRRRRRRRRRRRRRRRRW R:RRRRHMR8#0_oDFH:OR=]R''R;
RRRRRRRRRRRRRWRRq)77RH:RM#RR0D8_FOoH_OPC05FsRR4jRI8FMR0Fj;2R
RRRRRRRRRRRRRRRRqW7a:qRRRHMR8#0_oDFHPO_CFO0s45RRFR8IFM0R
j2RRRRRRRRRRRRR2RR;R
R

RRCRM81)A_qjv.c.UGhW)h;N

sHOE00COkRsC1)A_qjv.c.UGhW)h_Bq)]VRFR_1A).qvjGcU.hh)W#RH
oLCH
MRCRM81)A_qjv.c.UGhW)h_Bq)]R;RR---R_1A).qvjGcU.hh)W


-------------------------------------
--S---R_1A)cqvji_c
---------------------------------------
LDHs$NsR Q  k;
#QCR 3  1_a7pQmtB4_4nNc3D
D;kR#CQ   371a_tpmQzB_ht1Qh3 7N;DD
Ck#R Q  03#8F_Do_HON0sHED3NDz;
1Q R 3  MCkls_HO#308q;pp
M
C0$H0R_1A)cqvji_cR
H#
oRRCsMCH5ORRR
RSRRRWa)Q m_v7: RRs#0HRMo:"=R.X6n4;n"R-R-RMONRRLC.X6n4FnRs4R6.RXUF4sRjX.ccsRFRc.jU
X.RRRSR R)qv7_mR7 R#:R0MsHo=R:R6".nnX4"R;R-O-RNLMRC6R.nnX4RRFs6X4.UsRFR.4jcRXcF.sRjXcU.R
RRRRRRRRRRQQhaR_j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QanRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ(a_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QaqRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQAa_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQwa_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jjRR
RRRRRRRRRRRR2;R
RRRRRRRRRb0Fs5RR
RRRRRRRRRRRRR)RR7qqaRF:Rk#0R0D8_FOoH_OPC05FsRR46RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRp)Bi:RRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRp)Bi: RRRHMR8#0_oDFH:OR=]R''R;
RRRRRRRRRRRRR)RR RRRRH:RM#RR0D8_FOoHRR:=';]'
RRRRRRRRRRRRRRRR7)q7:)RRRHMR8#0_oDFHPO_CFO0s45Rj8RRF0IMF2RjRR;
RRRRRRRRRRRRRWRRBRpiRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRRWRRB piRH:RM#RR0D8_FOoHRR:=';]'
RRRRRRRRRRRRRRRRRW R:RRRRHMR8#0_oDFH:OR=]R''R;
RRRRRRRRRRRRRWRRq)77RH:RM#RR0D8_FOoH_OPC05FsRR4jRI8FMR0Fj;2R
RRRRRRRRRRRRRRRR1vqi:RRRRHMR8#0_oDFHPO_CFO0s45R68RRF0IMF2RjRR;
RRRRRRRRRRRRRWRR7qqaRH:RM#RR0D8_FOoH_OPC05FsRR468MFI0jFR2R
RRRRRRRRRRRRRR
2;RRR
RM
C8AR1_v)qccj_i
;
NEsOHO0C0CksR_1A)cqvji_c_FeRVAR1_v)qccj_i#RH
oLCH
MRCRM81)A_qjvc__cieR;RR---R_1A)cqvji_c
-

-------------------------------------S-
-R--1)A_qjvc_hci)-
--------------------------------------H
DLssN$ RQ 
 ;kR#CQ   371a_tpmQ4B_43ncN;DD
Ck#R Q  a317m_pt_QBzQh1t7h 3DND;#
kC RQ # 30D8_FOoH_HNs0NE3D
D;zR1 Q   3lMkCOsH_8#03pqp;C

M00H$AR1_v)qccj_iRh)H
#
RCRoMHCsORR5
SRRRWRR) Qa_7vm RR:#H0sM:oR=.R"64nXnR";RR--ORNML.CR64nXnsRFR.64XFURsjR4.ccXRRFs.UjcXR.
RRSRRq) 7m_v7R R:0R#soHMRR:="n.6X"4n;-RR-NROMCRLRn.6XR4nF6sR4U.XRRFs4cj.XFcRsjR.c.UX
RRRRRRRRRRRQahQ_:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQna_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QagRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQqa_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ a_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjRj"
RRRRRRRRRRRR;2R
RRRRRRRRbRRF5s0RR
RRRRRRRRRRRRRR7R)qRaq:kRF00R#8F_Do_HOP0COFRs54R6R8MFI0jFR2
R;RRRRRRRRRRRRRRRR)iBphRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRR)iBp RR:HRMR#_08DHFoO=R:R''];R
RRRRRRRRRRRRRR R)RRRR:MRHR0R#8F_DoRHO:'=R]
';RRRRRRRRRRRRRRRR)7q7)RR:HRMR#_08DHFoOC_POs0F5jR4RFR8IFM0RRj2;R
RRRRRRRRRRRRRRBRWpRiR:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRBRWpRi :MRHR0R#8F_DoRHO:'=R]
';RRRRRRRRRRRRRRRRWR RRRR:HRMR#_08DHFoO=R:R''];R
RRRRRRRRRRRRRRqRW7R7):MRHR0R#8F_Do_HOP0COFRs54RjR8MFI0jFR2
R;RRRRRRRRRRRRRRRRviq1RRR:HRMR#_08DHFoOC_POs0F56R4RFR8IFM0RRj2;R
RRRRRRRRRRRRRR7RWqRaq:MRHR0R#8F_Do_HOP0COFRs5486RF0IMF2Rj
RRRRRRRRRRRRRRR2R;
RR
R
8CMR_1A)cqvji_ch
);
ONsECH0Os0kCAR1_v)qccj_i_h)eVRFR_1A)cqvji_chH)R#C
LoRHM
8CMR_1A)cqvji_che)_;RRR-R--1)A_qjvc_hci)


-------------------------------------
--S---R_1A)cqvji_ch-W
-------------------------------------D-
HNLssQ$R ;  
Ck#R Q  a317m_pt_QB4c4n3DND;#
kC RQ 1 3ap7_mBtQ_1zhQ th7D3NDk;
#QCR 3  #_08DHFoOs_NH30EN;DD
 z1R Q  k3MlHCsO0_#8p3qp
;
CHM001$RAq_)v_cjcWihR
H#
oRRCsMCH5ORRR
RSRRRWa)Q m_v7: RRs#0HRMo:"=R.X6n4;n"R-R-RMONRRLC.X6n4FnRs4R6.RXUF4sRjX.ccsRFRc.jU
X.RRRSR R)qv7_mR7 R#:R0MsHo=R:R6".nnX4"R;R-O-RNLMRC6R.nnX4RRFs6X4.UsRFR.4jcRXcF.sRjXcU.R
RRRRRRRRRRQQhaR_j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QanRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ(a_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QaqRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQAa_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQwa_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jjRR
RRRRRRRRRRRR2;R
RRRRRRRRRb0Fs5RR
RRRRRRRRRRRRR)RR7qqaRF:Rk#0R0D8_FOoH_OPC05FsRR46RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRp)Bi:RRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRp)Bi: RRRHMR8#0_oDFH:OR=]R''R;
RRRRRRRRRRRRR)RR RRRRH:RM#RR0D8_FOoHRR:=';]'
RRRRRRRRRRRRRRRR7)q7:)RRRHMR8#0_oDFHPO_CFO0s45Rj8RRF0IMF2RjRR;
RRRRRRRRRRRRRWRRBhpiRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRRWRRB piRH:RM#RR0D8_FOoHRR:=';]'
RRRRRRRRRRRRRRRRRW R:RRRRHMR8#0_oDFH:OR=]R''R;
RRRRRRRRRRRRRWRRq)77RH:RM#RR0D8_FOoH_OPC05FsRR4jRI8FMR0Fj;2R
RRRRRRRRRRRRRRRR1vqi:RRRRHMR8#0_oDFHPO_CFO0s45R68RRF0IMF2RjRR;
RRRRRRRRRRRRRWRR7qqaRH:RM#RR0D8_FOoH_OPC05FsRR468MFI0jFR2R
RRRRRRRRRRRRRR
2;RRR
RM
C8AR1_v)qccj_i;hW
s
NO0EHCkO0s1CRAq_)v_cjcWih_FeRVAR1_v)qccj_iRhWHL#
CMoHRM
C8AR1_v)qccj_i_hWeR;RR---R_1A)cqvji_ch
W

---------------------------------------
-S--AR1_v)qccj_ihh)W-
--------------------------------------H
DLssN$ RQ 
 ;kR#CQ   371a_tpmQ4B_43ncN;DD
Ck#R Q  a317m_pt_QBzQh1t7h 3DND;#
kC RQ # 30D8_FOoH_HNs0NE3D
D;zR1 Q   3lMkCOsH_8#03pqp;C

M00H$AR1_v)qccj_ihh)W#RH
R
RoCCMsRHO5RR
RRSRRQW)av _mR7 :0R#soHMRR:="n.6X"4n;-RR-NROMCRLRn.6XR4nF6sR4U.XRRFs4cj.XFcRsjR.c.UX
SRRR)RR _q7v m7RRR:#H0sM:oR=.R"64nXnR";RR--ORNML.CR64nXnsRFR.64XFURsjR4.ccXRRFs.UjcXR.
RRRRRRRRRhRQQja_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QadRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQca_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQUa_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QaARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQBa_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QawRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"RR
RRRRRRRRR2RRRR;
RRRRRRRRRsbF0
5RRRRRRRRRRRRRRRRR)a7qqRR:FRk0#_08DHFoOC_POs0F56R4RFR8IFM0RRj2;R
RRRRRRRRRRRRRRBR)pRih:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRBR)pRi :MRHR0R#8F_DoRHO:'=R]
';RRRRRRRRRRRRRRRR)R RRRR:HRMR#_08DHFoO=R:R''];R
RRRRRRRRRRRRRRqR)7R7):MRHR0R#8F_Do_HOP0COFRs54RjR8MFI0jFR2
R;RRRRRRRRRRRRRRRRWiBphRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRRWiBp RR:HRMR#_08DHFoO=R:R''];R
RRRRRRRRRRRRRR RWRRRR:MRHR0R#8F_DoRHO:'=R]
';RRRRRRRRRRRRRRRRW7q7)RR:HRMR#_08DHFoOC_POs0F5jR4RFR8IFM0RRj2;R
RRRRRRRRRRRRRRqRv1RiR:MRHR0R#8F_Do_HOP0COFRs54R6R8MFI0jFR2
R;RRRRRRRRRRRRRRRRWa7qqRR:HRMR#_08DHFoOC_POs0F56R4RI8FMR0FjR2
RRRRRRRRRRRRR;R2

RRRCR
M18RAq_)v_cjc)ihh
W;
ONsECH0Os0kCAR1_v)qccj_ihh)WR_eF1VRAq_)v_cjc)ihhHWR#C
LoRHM
8CMR_1A)cqvji_chW)h_Re;R-R--AR1_v)qccj_ihh)W


DsHLNRs$HCCC;#
kCCRHC#C30D8_FOoH_n44cD3NDk;
#HCRC3CC#_08DHFoOs_NH30EN;DD
Ck#RCHCC03#8F_Do_HOkHM#o8MC3DND;C

M00H$sSbCF_HS
H#
FSbs50S
SSSLC#_M:SSSSHM#_08DHFoOS;S-a-KqCtRMDNLCRRRRRRRRRRR
SSS#VEH0:SSSSHM#_08DHFoOS;S-a-Kq#tRE0HVRRRRRRRRRRRR
SSS0	ODSSS:H#MS0D8_FOoH;-SS-qKatDROFRO	RRRRRRRRR
RRSkSSb08NC:SSSSHM#_08DHFoOS;S-a-KqktRb08NCRRRRRRRRRRR
SSS#S8HSSS:H#MS0D8_FOoH;-SS-qKatCR#sDHNR08NNMRHR
RRSlSSFS8CSH:SM0S#8F_Do;HOS-S-KtaqR8lFCRRRRRRRRRRRRSR
SHSExS_LSH:SM0S#8F_Do;HOS-S-KtaqRoEHERRXO0FMsRFDRSR
S8S#FSSS:kSF00S#8F_Do;HOS-S-KtaqRs#CHRND8NN0R0FkRSR
SFS8kS04SF:Sk#0S0D8_FOoH;-SS-shFlRNDQkMb0CRODFDRkk0b0
R4S8SSFjk0SSS:FSk0#_08DHFoOS;S-F-hsDlNRbQMkO0RCRDDFbk0kj0R
SSS848sSSS:H#MS0D8_FOoH;-SS-shFlRNDmbk0kO0RCRDDHkMb0
R4S8SS8SsjSH:SM0S#8F_Do;HOS-S-hlFsNmDRkk0b0CRODHDRM0bkRSj
SCSFbSHMSH:SM0S#8F_Do;HOS-S-hlFsNmDRk0bk-N MLRDCRRRRRSR
SFSEDS8S:MSHS8#0_oDFHSO;Sh--FNslDMRQbRk0ODCDRMOF0DsFRS
SS0s#HSFS:MSHS8#0_oDFHSO;Sh--FNslDMRQbRk0ODCDR#sCCR0RRS
SSOHMDS	S:MSHS8#0_oDFHSO;Sh--FNslDMRQbRk0ODCDRFODOR	RRS
SS0FkOSD	SH:SM0S#8F_Do;HOS-S-hlFsNmDRkk0b0CRODODRD	FORSR
SLSOHS0S:MSHS8#0_oDFHPO_CFO0s6R5RI8FMR0FjS2;-F-BMoVHkFsHMHRL0R#RRS
SS8bNHSMS:MSHS8#0_oDFHSO;Su--qH7RM0bkRRRRRRRRRSR
SNSb80FkSSS:FSk0#_08DHFoOS;S-q-u7kRF00bkRRRRRRRRRS
SS8bNFSCMSF:Sk#0S0D8_FOoHR-SS-7uqR0FkbRk0CLMNDRCR
SSS2
;
CRM8b_sCH
F;
ONsECH0Os0kCsRbCF_H_FPRVsRbCF_HR
H#So#HMSNDbHN8M4_M,OHMDM	_.N,b8_HMM:dSS8#0_oDFH
O;So#HMSNDHvM_zMX_cSS:#_08DHFoOS;
#MHoNEDSF_D8q.h7S#:S0D8_FOoH;#
SHNoMD8S8sMj_4:4SS8#0_oDFH
O;So#HMSNDFOk0DM	_4:.SS8#0_oDFH
O;So#HMSND848s_dM4S#:S0D8_FOoH;#
SHNoMD4SMcSSS:0S#8F_Do;HO
HS#oDMNSk8F0C_so__jMSS:#_08DHFoOS;
#MHoN)DSCFo_sH_WshC_4:(SS8#0_oDFH
O;So#HMSNDMS4USSS:#_08DHFoOS;
#MHoNMDS4SgSS#:S0D8_FOoH;#
SHNoMDsS0HN#00:CSS8#0_oDFH
O;So#HMSNDFOk0DM	_.:.SS8#0_oDFH
O;So#HMSNDMS.nSSS:#_08DHFoOS;
#MHoNFDSCMM__cM.S#:S0D8_FOoH;#
SHNoMD0S[Nko_b08NCd_MjSS:#_08DHFoOS;
#MHoN8DSHsM_Cjo_S#:S0D8_FOoH;#
SHNoMD8RRHsM_C4o_S#:S0D8_FOoH;#
SHNoMDFS8ks0_Cjo_S#:S0D8_FOoH;#
SHNoMDFS8ks0_C4o_S#:S0D8_FOoH;#
SHNoMDsS0HN#00JC_S#:S0D8_FOoH;#
SHNoMD0S[NFo_CC_soSS:#_08DHFoOS;
#MHoN0DSC4lb,l0CbS.S:0S#8F_Do_HOP0COF5sR4FR8IFM0R;j2
HS#oDMNSk8F0S_jS#:S0D8_FOoH;-SS-HSIsVCRFbsRFRs0#MHoNkDR#CNo
oLCHSM
[o0N_8kbN_0CMSdj<M=SF50SLC#_MMRN8MR5Fk0Rb08NC;22
SS
#S8FSS<=8_HMs_CojS;
80Fk4<RS=8RSHsM_C4o_;-
-------------------------------------------------------------Sb
SNM8H__M4HSS:bOsFCS##5k8F0C_so,_jR8bNHRM,#VEH0S2
SLSSCMoH
SSSSVSHSE5#H=V0'24'SC0EMS
SSSSSbHN8M4_MSS<=80Fk_osC_
j;SSSSS#CDCS
SSSSSbHN8M4_MSS<=bHN8MS;
SSSSCRM8H
V;SSSSCSM8bOsFC;##
SS
HDMO	._M_:HSSFbsO#C#S#5L_,CMRD0O	H,RM	OD2S
SSCSLo
HMSSSSSSHV5_L#C'M=4S'20MEC
SSSSHSSM	OD_SM.<0=SO;D	
SSSSDSC#SC
SSSSSOHMDM	_.=S<SOHMD
	;SSSSS8CMR;HV
SSSS8CMRFbsO#C#;S

8_HMs_CojS_H:sSbF#OC#HS5M	OD_,M.R0s#H
F2SSSSLHCoMS
SSHSSVsS5#F0H=''42ES0CSM
SSSSSM8H_osC_<jS=jS''S;
SSSSCHD#VHS5M	OD_RM.'CCPMN0RMH8RM	OD_=M.'24'RC0EMS
SSSSS8_HMs_Coj=S<S8bNHMM_4S;
SSSSCRM8H
V;SSSSCRM8bOsFC;##
------------------------------------------------------------S-SSSS
bHN8Md_M_:HSSFbsO#C#S#5L_,CMRM8H_osC_Rj,bHN8MS2
SLSSCMoH
SSSSVSHS#5L_=CM'24'SC0EMS
SSSSSbHN8Md_MSS<=8_HMs_CojS;
SSSSCCD#
SSSSbSSNM8H_SMd<b=SNM8H;S
SSCSSMH8RVS;
SCSSMb8SsCFO#
#;S8
SHsM_C4o__:HSSFbsO#C#SM5HO_D	MR.,sH#0FS2
SLSSCMoH
SSSSVSHS#5s0=HF'24'SC0EMS
SSSSS8_HMs_Co4=S<S''j;S
SSCSSDV#HSM5HO_D	M'.RCMPC0MRN8MRHO_D	M'.=jR'20MEC
SSSSHSSV[S50_NokNb80MC_d'j=4S'20MEC
SSSSSSS8_HMs_Co4=S<S8bNHMM_dS;
SSSSS8CMR;HV
SSSSMSC8VRH;S
SSMSC8sRbF#OC#-;
-------------------------------------------------------------SS
E8FD_7qh.=R<RHOL0254R8NMRDEF8
;
RSRR-M-QbRk0vRzXR
RSSl0Cb<4S=FSEDq8_hR7.&LROHj052
;
S_HMv_zXMHc_Sb:SsCFO#5#S0bCl48,RF_k0j8,RHsM_Cjo_,NRb82HM
RRRSSSSLHCoMR
RRSSSSNSO#0CSC4lbR
H#RSRRSSSSIMECSj"j">S=
RRRSSSSSMSH_Xvz_RMc<8=RHsM_Cjo_;R
RRSSSSESIC"MSjS4"=R>
RSRSSSSSHvM_zMX_c=R<R8bNH
M;RSRRSSSSIMECSj"4">S=
RRRSSSSSMSH_Xvz_RMc<8=RF_k0jR;
RSRSSISSESCM""44S
=>RSRRSSSSS_HMv_zXM<cR=FR8kj0_;R
RRSSSSESICFMR0sEC#=RS>R
RRSSSSHSSMz_vXc_MRR<=';j'
RRRSSSSS8CMR#ONCR;
RSRSSMSC8sRbF#OC#
;
------------------------80FkjCRoMNCs0-C-----------------------------
FS8kj0__:HSSFbsO#C#SF5l8RC,8_HMs_Co4H,RMz_vXc_M2S
SSoLCHSM
SHSSVlS5F=8C'24'SC0EMS
SS8SSF_k0j=S<SM8H_osC_
4;SSSSCCD#
SSSSFS8kj0_SS<=HvM_zMX_cS;
SCSSMH8RVS;
SMSC8sRbF#OC#S;

FS8kS0j<8=SF_k0j-;
-----------------------------------------------------------------S--
-S-mbk0k)0RC#oH0
CsS8
SF_k0s_CojS_H:sSbF#OC#FS5kD0O	4_M.s,R#F0H2S
SSCSLo
HMSSSSSSHV50s#H'F=4S'20MEC
SSSS8SSF_k0s_Coj=S<S''j;S
SSCSSDV#HSk5F0	OD_.M4RP'CCRM0NRM8FOk0DM	_4'.=4R'20MEC
SSSS8SSF_k0s_Coj=S<Ss88j4_M4S;
SSSSCRM8H
V;SSSSCRM8bOsFC;##
-
S-GvkCV#RFmsRkk0b0CRso0H#C
s#S8
SF_k0s_CojR_MSR<=MRF080Fk_osC_
j;SgM4RSSS<M=RF50RFOk0DM	_4F.RsLROH.052
2;S)
SCFo_sH_WshC_4H(_Sb:SsCFO#5#SO0LH5,.2Rk8F0C_so__jM8,R82sj
SSSSCSLo
HMSSSSSVSHSL5OH.0524=''02SE
CMSSSSS)SSCFo_sH_WshC_4<(S=FS8ks0_Cjo__
M;SSSSSDSC#SC
SSSSSCS)os_F_sWHC4_h(=S<Ss88jS;
SSSSS8CMR;HV
SSSSMSC8sRbF#OC#S;

4SMUS_HS:SSSFbsO#C#S45Mg8,RF_k0s_Co48,RF_k0s_CojS2
SSSSLHCoMS
SSSSSH5VSM=4g'24'SC0EMS
SSSSSSUM4SS<=80Fk_osC_
4;SSSSSDSC#SC
SSSSS4SMU=S<Sk8F0C_so;_j
SSSSCSSMH8RVS;
SSSSCRM8bOsFC;##
M
S4Hc_SSSS:sSbF#OC#OS5L5H0dR2,)_CoFWs_H_sCh,4(RUM42SS
SSSSLHCoMS
SSSSSH5VSO0LH5=d2'24'SC0EMS
SSSSSScM4SS<=)_CoFWs_H_sCh;4(
SSSSCSSD
#CSSSSSMSS4<cS=4SMUS;
SSSSS8CMR;HV
SSSSMSC8sRbF#OC#S;
SSSS
NSb80Fk_SHSSb:SsCFO#5#SlCF8,FR8ks0_C4o_,4RMcS2
SSSSLHCoMS
SSSSSH5VSlCF8=''42ES0CSM
SSSSSNSb80FkSS<=80Fk_osC_
4;SSSSSDSC#SC
SSSSSNSb80FkSS<=M;4c
SSSSCSSMH8RVS;
SSSSCRM8bOsFC;##
-
S-qKat#Rq#MHo#

SSs88j4_M4S_HSb:SsCFO#5#S#VEH00,Rs0H#N_0CJ8,R82sj
SSSSCSLo
HMSSSSSVSHSE5#H=V0'24'SC0EMS
SSSSSSs88j4_M4=S<SH0s#00NC;_J
SSSSCSSD
#CSSSSS8SS8_sjMS44<8=S8;sj
SSSSCSSMH8RVS;
SSSSCRM8bOsFC;##
F
SkD0O	4_M.S_HSb:SsCFO#5#SLC#_M0,RO,D	R0FkO2D	
SSSSCSLo
HMSSSSSVSHS#5L_=CM'24'SC0EMS
SSSSSS0FkO_D	MS4.<0=SO;D	
SSSSCSSD
#CSSSSSFSSkD0O	4_M.=S<S0FkO;D	
SSSSCSSMH8RVS;
SSSSCRM8bOsFC;##
SSSSSS
848s_dM4_SHS:sSbF#OC#LS5#M_C,FR8ks0_Cjo_,8R8s
42SSSSSoLCHSM
SSSSSSHV5_L#C'M=4S'20MEC
SSSSSSS848s_dM4SS<=80Fk_osC_
j;SSSSSDSC#SC
SSSSS8S8sM4_4<dS=8S8s
4;SSSSSMSC8VRH;S
SSCSSMb8RsCFO#
#;
-S-KtaqRosCHC#0sSR
80Fk_osC_H4_SSS:bOsFCS##50FkO_D	M,4.R0s#H
F2SSSSSoLCHSM
SSSSSSHV50s#H'F=4S'20MEC
SSSSSSS80Fk_osC_<4S=jS''S;
SSSSS#CDH5VSFOk0DM	_4'.RCMPC0MRN8kRF0	OD_.M4=''j2ER0CSM
SSSSSFS8ks0_C4o_SS<=848s_dM4;S
SSSSSCRM8H
V;SSSSS8CMRFbsO#C#;S
SS
SS----------------------------------------------------------------------------

---m-Skk0b0MR NCLDRopFH-O
--
--------------------------------------------------------------------------
--Sm-- sRaHN#00)CRC#oH0
CsSH0s#00NCS_H:sSbF#OC##S5E0HV,8R#HF,RCMbH2S
SSCSLo
HMSSSSSSHV5H#EV'0=4S'20MEC
SSSS0SSs0H#NS0C<#=S8
H;SSSSS#CDCS
SSSSS0#sH0CN0SS<=FHCbMS;
SSSSCRM8H
V;SSSSCRM8bOsFC;##
0
Ss0H#N_0CJS_H:sSbF#OC#FS5kD0O	._M.s,R#F0H2S
SSCSLo
HMSSSSSSHV50s#H'F=4S'20MEC
SSSS0SSs0H#N_0CJ=S<S''j;S
SSCSSDV#HSk5F0	OD_.M.RP'CCRM0NRM8FOk0DM	_.=.RR''42ER0CSM
SSSSSH0s#00NCS_J<0=Ss0H#N;0C
SSSSMSC8VRH;S
SSMSC8sRbF#OC#S;
S
SSSK--aRqtsHCo#s0C
kSF0	OD_.M._:HSSFbsO#C#S#5L_,CMRD0O	F,RkD0O	S2
SLSSCMoH
SSSSVSHS#5L_=CM'24'SC0EMS
SSSSSFOk0DM	_.<.S=OS0D
	;SSSSS#CDCS
SSSSSFOk0DM	_.<.S=kSF0	OD;S
SSCSSMH8RVS;
SCSSMb8RsCFO#
#;S[
S0_NoFsC_CHo_Sb:SsCFO#5#SFOk0DM	_.R.,sH#0FS2
SLSSCMoH
SSSSVSHS#5s0=HF'24'SC0EMS
SSSSS[o0N__FCsSCo<'=Sj
';SSSSS#CDH5VSFOk0DM	_.'.RCMPC0MRN8kRF0	OD_.M.Rj=''02RE
CMSSSSSVSHS05[Nko_b08NCd_Mj4=''02SE
CMSSSSS[SS0_NoFsC_C<oS=NSb8_HMM
d;SSSSSMSC8VRH;S
SSCSSMH8RVS;
SCSSMb8RsCFO#
#;SR
RRCS0lSb.<O=SL5H06&2RRHOL025c;RR
R-S-SMFC_MM_.Hc_Sb:SsCFO#5#SO0LH5,62O0LH5,c2RbFCHRM,0#sH0CN0_RJ2
SRRF_CMM._McS_H:sSbF#OC#0S5C.lb,CRFb,HMRH0s#00NC2_JRR
RSSSSSoLCH
MRRSRSSSSS-N-O#OCSL5H06&2RRHOL025cRRH#
SRRSSSSS#ONCCS0lRb.H
#RRSRSSSSSSCIEMjS"j="S>RR
RSSSSSSSF_CMM._Mc=S<S''j;RR
RSSSSSSSIMECS4"j">S=RR
RSSSSSFSSCMM__cM.SS<=';4'RR
RSSSSSISSESCM""4jSR=>
SRRSSSSSCSFM__MMS.c<F=SCMbH;RR
RSSSSSSSIMECS4"4">S=
RRRSSSSSFSSCMM__cM.SS<=0#sH0CN0_RJ;
RRRSSSSSISSERCMFC0EsS#S=
>RRSRRSSSSSCSFM__MMS.c<'=SjR';
RRRSSSSSMSC8NRO#RC;
RRRSSSSS8CMRFbsO#C#;

SSnM._SHSSb:SsCFO#5#SlCF8,0R[NFo_CC_soF,RCMM__cM.2S
SSCSLo
HMSSSSSSHV58lFC4=''02SE
CMSSSSS.SMn=S<SN[0oC_F_osC;S
SSCSSD
#CSSSSS.SMn=S<SMFC_MM_.
c;SSSSS8CMR;HV
SSSS8CMRFbsO#C#;S

bFN8C<MR=FRM0ER5HLx_R8NMRnM.2S;

8CMRCbs__HFP
;
------------------------------------------------------------------------
S--SSSS1QA_m-
----------------------------------------------------------------------
-
DsHLNRs$HCCC;#
kCCRHC#C30D8_FOoH_n44cD3NDk;
#HCRC3CC#_08DHFoOs_NH30EN;DD
Ck#RCHCC03#8F_Do_HOkHM#o8MC3DND;-
-DsHLNSs$I	Fs;#
kCFSIs#	30D8_FOoH_a1A3DND;C

M00H$AS1_RQmH
#
SMoCCOsHRS5
S Sht)_aQ tt)RR:LSH0SSSSSS:=';j'
SSSu_Qha YuSL:RHP0_CFO0s6R5RI8FMR0Fj:2S=jS"jjjjj
";SuSSzzppu:SSR0LHSSSSS=S:S''j;S
SS_Qm1haq77q)S#:R0MsHoSSSS=S:SA"1_Bpev"m1
SSS2S;
b0FsRS
S5S
S7z_maR_4SRSRRRR:H#MR0D8_FOoH;S
S7z_maR_jSRSRRRR:H#MR0D8_FOoH;S
SBBpmih_ q ApSRS:H#MR0D8_FOoH;S
SpBqa]h_Qu_zaezqp RS:H#MR0D8_FOoH;S
SQzhuap_BiSSS:MRHR8#0_oDFH
O;SSS
SQ7_hS_4S:SSR0FkR8#0_oDFH
O;S_S7Qjh_SSSS:kRF00R#8F_Do;HO
mSSzzauah_ q ApSRS:H#MR0D8_FOoHS':=]
';SzSmaauz_iBpS:SSRRHM#_08DHFoOS;
SBuqi qt_huQS:SSRFHMk#0S0k8_DHFoOS
S2
;RSCS
M18RAm_QRN;
0H0sLCk0RM#$_NLDOL	_FFGRVAR1_RQm:FROlMbFCRM0H0#Rs;kC
s
NO0EHCkO0s1CRAm_Q_FeRVAR1_RQmH
#
SlOFbCFMMb0SsHC_Fb
SFSs05S
SSDEF8SS:HSMR#_08DHFoOS;
S#Ss0SHF:MSHS8#0_oDFH
O;SLSS#M_CSH:SM0S#8F_Do;HO
SSS#VEH0SS:H#MS0D8_FOoH;S
SSD0O	SS:H#MS0D8_FOoH;S
SSOHMD:	SSSHM#_08DHFoOS;
SkSF0	ODSH:SM0S#8F_Do;HO
SSSkNb80:CSSSHM#_08DHFoOS;
SCSFbSHM:MSHS8#0_oDFH
O;S#SS8SHS:MSHS8#0_oDFH
O;SlSSFS8C:MSHS8#0_oDFH
O;SESSHLx_SH:SM0S#8F_Do;HO
SSS#S8FSF:Sk#0S0D8_FOoH;S
SSk8F0:4SS0FkS8#0_oDFH
O;S8SSFjk0SF:Sk#0S0D8_FOoH;S
SSs884SS:H#MS0D8_FOoH;S
SSs88jSS:H#MS0D8_FOoH;S
SS8bNH:MSSSHM#_08DHFoOS;
SNSb80FkSF:Sk#0S0D8_FOoH;S
SS8bNFSCM:kSF00S#8F_Do;HO
SSSO0LHSH:SM0S#8F_Do_HOP0COF5sS6FR8IFM0R
j2S2SS;C
SMO8RFFlbM0CM;S

#MHoNHDSM	OD_RM,FOk0DM	_,MRHO,D	R0FkO,D	#S8F:0S#8F_Do;HO
SS
#MHoNLDS#M_CS#:S0D8_FOoHS':=jS';-F-AkNM8s#$RORNMCLMNDRCRRRRRRRRRR#
SHNoMDES#HSV0:0S#8F_DoSHO:j=''-;S-kAFMs8N$OR#N#MRE0HVRRRRRRRRRRRR
HS#oDMNSD0O	SS:#_08DHFoO=S:';j'SA--F8kMNRs$#MONRFODOR	RRRRRRRRRRSR
#MHoNkDSb08NCSS:#_08DHFoO=S:';j'SA--F8kMNRs$#MONR8kbNR0CRRRRRRRRRSR
#MHoN#DS8SHS:0S#8F_DoSHO:j=''-;S-kAFMs8N$OR#N#MRCNsHDNR80HNRMRRR
HS#oDMNS8lFCSS:#_08DHFoO=S:';j'SA--F8kMNRs$#MONR8lFCRRRRRRRRRRRRSR
#MHoNEDSHLx_S#:S0D8_FOoHS':=4S';-F-AkNM8s#$RORNMa#sH0CN0RMOF0DsFR

SSo#HMSNDb_HMO0LH:0S#8F_Do_HOP0COF6s5RI8FMR0Fj
2;So#HMSNDM_Co0osH:0S#8F_Do;HO
HS#oDMNSDbkDb_kS#:S0D8_FOoH;#
SHNoMDFSEDF8,CMbH,8bNF,CMbFN8kb0,NM8HS#:S0D8_FOoH;C
Lo
HMSb
SHOM_LSH0<a=Sma_17tpmQ BeB)amSQ5uhY_au; 2
CSMos_0H<oS=mSa_71apQmtBhS5 at_)tQt ;)2
kSbDkD_b<SS=mSa_71apQmtBuS5zzppu
2;
MSHO_D	M=S<RhSQu_zaBRpiGRFsM_Co0osH;F
SkD0O	<_M=zSmaauz_iBpRsGFRoMC_H0soS;
HDMO	=S<SOHMDM	_R8NMRmBpB i_hpqA S;
FOk0D<	S=kSF0	OD_NMRMB8RpimB_q hA;p 
SS
E8FDSS<=pBqa]h_Qu_zaezqp S;
FHCbM=S<Samzu_za Ahqp
 ;Su
SqqBitu _QHh_Sb:SsCFO#5#SbFN8CRM,bFN8kR0,uiqBq_t u2Qh
CSLo
HMSNSb8SHM<u=SqqBitu _Q
h;SVSHSN5b8MFC=''42ER0CSM
SqSuBtiq Q_uh=S<S''Z;S
SCCD#
SSSuiqBq_t uSQh<b=SNk8F0S;
S8CMR;HV
MSC8sRbF#OC#-;
----------------------------------------------------------------Sb
SsHC_FS_H:sSbCF_H
FSbsl0RN5bS
SSSSDEF8>S=SDEF8S,
SsSS#F0HSS=>',j'
SSSS_L#C=MS>#SL_,CM
SSSSH#EV=0S>ES#H,V0
SSSSD0O	>S=SD0O	S,
SHSSM	ODSS=>HDMO	S,
SFSSkD0O	>S=S0FkO,D	
SSSS8kbNS0C=k>Sb08NCS,
SFSSCMbHSS=>FHCbMS,
S#SS8SHS=#>S8
H,SSSSlCF8SS=>lCF8,S
SSHSExS_L=E>SHLx_,S
SS8S#F=SS>8S#FS,
S8SSF4k0SS=>7h_Q_
4,SSSS80Fkj>S=SQ7_h,_j
SSSSs884>S=Sm7_z4a_,S
SS8S8s=jS>_S7m_zajS,
SbSSNM8HSS=>bHN8MS,
SbSSNk8F0>S=S8bNF,k0
SSSS8bNFSCM=b>SNC8FMS,
SOSSLSH0=b>SHOM_L
H0SSSS2C;
M18SAm_Q_
e;
--------------------------------------------------------------------
---S-SS1SSAA_t_
Qm---------------------------------------------------------------------
-
DsHLNRs$HCCC;#
kCCRHC#C30D8_FOoH_n44cD3NDk;
#HCRC3CC#_08DHFoOs_NH30EN;DD
Ck#RCHCC03#8F_Do_HOkHM#o8MC3DND;-
-DsHLNSs$I	Fs;#
kCFSIs#	30D8_FOoH_a1A3DND;C

M00H$AS1__tAQHmR#o
SCsMCH5OS
SSSh_ tat)QtR ):HRL0SSSS:SS=jS''S;
SQSuhY_au: SR0LH_OPC0RFs586RF0IMF2RjSS:="jjjj"jj;S
SSpuzpSzuSL:RHS0SSSSS:'=Sj
';SQSSma_1qqh7):7SRs#0HSMoSSSS:"=S1pA_emBv1S"
S;S2
SSS
FSbs50S
SSSuiqBq_t uSQhSSS:HkMF00S#8D_kFOoH;S
SSapqBQ]_hauz_peqz: SSSHMS8#0_oDFH
O;SBSSpimB_q hARp RRRRR:RRSSHMS8#0_oDFH
O;SQSShauz_iBpRRRRRRRRR:RRSSHMS8#0_oDFH
O;SmSSzzauap_BiRRRRRRRR:RRSSHMS8#0_oDFH
O;SmSSzzauah_ q ApSRS:H#MR0D8_FOoHS':=]
';S7SS_amz_R4RRRRRRRRRR:RRSSHMS8#0_oDFH
O;S7SS_amz_RjRRRRRRRRRR:RRSSHMS8#0_oDFH
O;S7SS__Qh4RRRRRRRRRRRR:RRS0FkS0S#8F_Do;HO
SSS7h_Q_RjRRRRRRRRRRRRR:kSF0#SS0D8_FOoH;S
SSmtpA_qpAwzw m)_zzauaF:SkS0S#_08DHFoOS
SS
2;CRM81tA_Am_Q;0
N0LsHkR0C#_$MLODN	F_LGVRFR_1AtQA_mRR:ObFlFMMC0#RHRk0sC
;
NEsOHO0C0CksR_1AtQA_mR_eF1VRAA_t_RQmH
#
SlOFbCFMMb0SsHC_Fb
SFSs05S
SSDEF8SS:HSMR#_08DHFoOS;
S#Ss0SHF:MSHS8#0_oDFH
O;SLSS#M_CSH:SM0S#8F_Do;HO
SSS#VEH0SS:H#MS0D8_FOoH;S
SSD0O	SS:H#MS0D8_FOoH;S
SSOHMD:	SSSHM#_08DHFoOS;
SkSF0	ODSH:SM0S#8F_Do;HO
SSSkNb80:CSSSHM#_08DHFoOS;
SCSFbSHM:MSHS8#0_oDFH
O;S#SS8SHS:MSHS8#0_oDFH
O;SlSSFS8C:MSHS8#0_oDFH
O;SESSHLx_SH:SM0S#8F_Do;HO
SSS#S8FSF:Sk#0S0D8_FOoH;S
SSk8F0:4SS0FkS8#0_oDFH
O;S8SSFjk0SF:Sk#0S0D8_FOoH;S
SSs884SS:H#MS0D8_FOoH;S
SSs88jSS:H#MS0D8_FOoH;S
SS8bNH:MSSSHM#_08DHFoOS;
SNSb80FkSF:Sk#0S0D8_FOoH;S
SS8bNFSCM:kSF00S#8F_Do;HO
SSSO0LHSH:SM0S#8F_Do_HOP0COF5sS6FR8IFM0R
j2S2SS;C
SMO8RFFlbM0CM;

SSo#HMSNDHDMO	,_MFOk0DM	_,OHMDF	,kD0O	8,#FSS:#_08DHFoOS;

HS#oDMNS_L#C:MSS8#0_oDFH:OS=''j;-S-AMFk8$NsRN#OMMRCNCLDRRRRRRRRR
RRSo#HMSND#VEH0SS:#_08DHFoO=S:';j'SA--F8kMNRs$#MONRH#EVR0RRRRRRRRRRSR
#MHoN0DSOSD	:0S#8F_DoSHO:j=''-;S-kAFMs8N$OR#NOMRD	FORRRRRRRRRRRR
HS#oDMNS8kbNS0C:0S#8F_DoSHO:j=''-;S-kAFMs8N$OR#NkMRb08NCRRRRRRRRRRR
HS#oDMNSH#8SSS:#_08DHFoO=S:';j'SA--F8kMNRs$#MONRs#CHRND8NN0RRHMRSR
#MHoNlDSFS8C:0S#8F_DoSHO:j=''-;S-kAFMs8N$OR#NlMRFR8CRRRRRRRRRRRR
HS#oDMNSxEH_:LSS8#0_oDFH:OS=''4;-S-AMFk8$NsRN#OMsRaHN#00OCRFsM0F
DRS#
SHNoMDFSEDF8,CMbH,8bNF,CMbFN8kb0,NM8HS#:S0D8_FOoH;

SSo#HMSNDM_Co0osH:0S#8F_Do;HO
HS#oDMNSDbkDb_kS#:S0D8_FOoH;#
SHNoMDHSbML_OHS0:#_08DHFoOC_POs0F586RF0IMF2Rj;

SLHCoM

SSoMC_H0so=S<S_am1pa7mBtQS 5ht)_aQ tt)
2;SMbH_HOL0=S<S_am1pa7mBtQea Bm5)Su_Qha Yu2S;
bDkD_SkbSS<=a1m_am7ptSQB5puzp2zu;S

HDMO	S_M<S=RQzhuap_BiFRGsCRMos_0H
o;S0FkO_D	M=S<Samzu_zaBRpiGRFsM_Co0osH;H
SM	ODSS<=HDMO	R_MNRM8BBpmih_ q Ap;F
SkD0O	=S<S0FkO_D	MMRN8pRBm_Bi Ahqp
 ;SE
SFSD8<p=Sq]aB_uQhzea_q pz;F
SCMbHSS<=muzaz a_hpqA S;

qSuBtiq Q_uhS_H:sSbF#OC#bS5NC8FMb,RNk8F0u,RqqBitu _Q
h2SoLCHSM
S8bNH<MS=qSuBtiq Q_uhS;
SSHV58bNF=CM'24'RC0EMS
SSBuqi qt_huQSS<=';Z'
CSSD
#CSuSSqqBitu _Q<hS=NSb80Fk;S
SCRM8H
V;S8CMRFbsO#C#;

SSmtpA_qpAwzw m)_zzaua=S<S8bNH
M;-----------------------------------------------------------------
S
SCbs__HFHSS:b_sCHSF
b0FsRblNSS5
SESSFSD8=E>SF,D8
SSSS0s#H=FS>jS''S,
SLSS#M_CSS=>LC#_MS,
S#SSE0HVSS=>#VEH0S,
S0SSOSD	=0>SO,D	
SSSSOHMD=	S>MSHO,D	
SSSS0FkOSD	=F>SkD0O	S,
SkSSb08NC>S=S8kbN,0C
SSSSbFCH=MS>CSFb,HM
SSSSH#8S>S=SH#8,S
SSFSl8=CS>FSl8
C,SSSSE_HxL>S=SxEH_
L,SSSS#S8FSS=>#,8F
SSSSk8F0=4S>_S7Q4h_,S
SSFS8kS0j=7>S__QhjS,
S8SS8Ss4=7>S_amz_
4,SSSS8j8sSS=>7z_ma,_j
SSSS8bNH=MS>NSb8,HM
SSSS8bNFSk0=b>SNk8F0S,
SbSSNC8FM>S=S8bNF,CM
SSSSHOL0>S=SMbH_HOL0S
SS;S2
8CMS_1AtQA_m;_e
-
--------------------------------------------------------------
---S-SS1SSAA_t
----------------------------------------------------------------
-
DsHLNRs$HCCC;#
kCCRHC#C30D8_FOoH_n44cD3NDk;
#HCRC3CC#_08DHFoOs_NH30EN;DD
Ck#RCHCC03#8F_Do_HOkHM#o8MC3DND;-
-DsHLNSs$I	Fs;#
kCFSIs#	30D8_FOoH_a1A3DND;C

M00H$AS1_StAH
#
b0FsSS5
SmtpA_qpAwzw m)_zzauaSSS:kSF00S#8F_Do;HO
zSS1_ )1hQtqap_mp_tmpAq_wAzwS ):MSHS8#0_oDFHSO
S
2;
8CMS_1At
A;Ns00H0LkC$R#MD_LN_O	LRFGF1VRAA_tRO:RFFlbM0CMRRH#0Csk;N

sHOE00COkSsC1tA_AR_eF1VRAA_tR
H#LHCoMt
SpqmApz_Aw)w _amzuSza<z=S1_ )1hQtqap_mp_tmpAq_wAzw; )
8CMR_1AteA_;



H
DLssN$CRHC
C;kR#CHCCC38#0_oDFH4O_43ncN;DD
Ck#RCHCC03#8F_Do_HON0sHED3NDk;
#HCRC3CC#_08DHFoOM_k#MHoCN83D
D;
0CMHS0$1WA_qA)vmSmaHb#
FSs05S
SAammSH:SM0S#8F_Do;HO
1SS4:SSSSHM#_08DHFoOS;
SS1jSH:SM0S#8F_Do;HO
2SS;C

M18RAq_W)mvAm
a;Ns00H0LkC$R#MD_LN_O	LRFGF1VRAq_W)mvAm:aRRlOFbCFMMH0R#sR0k
C;Ns00H0LkC$R#MF_MbMskCVRFR_1AWvq)AammRO:RFFlbM0CMRRH#0Csk;-

-----------------------------------------------------------
-SSSS_1AQ7m_1-
----------------------------------------------------------
-
DsHLNRs$HCCC;#
kCCRHC#C30D8_FOoH_n44cD3NDk;
#HCRC3CC#_08DHFoOs_NH30EN;DD
Ck#RCHCC03#8F_Do_HOkHM#o8MC3DND;-
-DsHLNSs$I	Fs;#
kCFSIs#	30D8_FOoH_a1A3DND;S

-H-7VsVCCHM0N#DRHNoMDoHMR
QmCHM001$SAm_Q_S71HS#
oCCMsSHO5S
SSth _Qa)t)t RL:RHS0SSSSS:'=Sj
';SuSSQah_YSu :HRL0C_POs0FRR568MFI0jFR2=S:Sj"jjjjj"S;
SmSQ_q1ah)7q7RS:#H0sMSoSS:SS=1S"Ae_p7m1_zzauaS"
S;S2
b
SFSs05S
SSm7_z4a_S:SSSSHM#_08DHFoO-;S-MRQbRk0Fbk0k40RRS
SSm7_zja_S:SSSSHM#_08DHFoO-;S-MRQbRk0Fbk0kj0RRS
SSmBpB i_hpqA SS:H#MS0D8_FOoH;-S-RFBDOC	RMDNLCh#R -WRRlOFlRFM0HFRMk/F0DROF#O	RS
SSQ7_hS_4SSS:FSk0#_08DHFoO-;S-kRm00bkRbHMk40R
SSS7h_Q_SjSSF:Sk#0S0D8_FOoH;-S-R0mkbRk0HkMb0
RjSmSSzzauah_ q ApSRS:H#MR0D8_FOoHS':=]S';-m-Rk0bk-N MLRDC
SSSpBqa]h_Qu_zaezqp SS:H#MS0D8_FOoH;-S-RbQMkO0RFsM0F
DRSQSShauz_iBpSSS:H#MS0D8_FOoH;-S-RbQMkO0RD	FORS
SSamzu_zaBSpiSH:SM0S#8F_Do;HOR-R-R0mkbRk0OODF	S
SSBuqi qt_huQSSS:HkMF00S#8D_kFOoH;-S-RCz#sR'#b	NONRoCbRHM-uR'qR7'Fbk0kR0R
SSSuiqBq_t u_QhASS:HkMF00S#8D_kFOoHSR--zs#C'b#RNNO	obCRH-MRRq'u7F'Rkk0b0
RRS2SS;C

M18RAm_Q_;71
0N0skHL0#CR$LM_D	NO_GLFRRFV1QA_m1_7RO:RFFlbM0CMRRH#0Csk;N

sHOE00COkRsC1QA_m1_7_FeRVAR1__Qm7H1R#-
S-HS#oDMN#-
------------------
--So#HMSNDHDMO	,_MFOk0DM	_,OHMDF	,kD0O	8,#FSS:#_08DHFoOS;

HS#oDMNS_L#C:MSS8#0_oDFH:OS=''j;-S-AMFk8$NsRN#OMMRCNCLDRRRRRRRRR
RRSo#HMSND#VEH0SS:#_08DHFoO=S:';j'SA--F8kMNRs$#MONRH#EVR0RRRRRRRRRRSR
#MHoN0DSOSD	:0S#8F_DoSHO:j=''-;S-kAFMs8N$OR#NOMRD	FORRRRRRRRRRRR
HS#oDMNS8kbNS0C:0S#8F_DoSHO:j=''-;S-kAFMs8N$OR#NkMRb08NCRRRRRRRRRRR
HS#oDMNSH#8SSS:#_08DHFoO=S:';j'SA--F8kMNRs$#MONRs#CHRND8NN0RRHMRSR
#MHoNlDSFS8C:0S#8F_DoSHO:j=''-;S-kAFMs8N$OR#NlMRFR8CRRRRRRRRRRRR
HS#oDMNSxEH_:LSS8#0_oDFH:OS=''4;-S-AMFk8$NsRN#OMsRaHN#00OCRFsM0F
DRS#
SHNoMDFSEDF8,CMbHS#:S0D8_FOoH;-S-aRECskCJH8sCRObN	CNoRMbHRb0$CkRl#L0RCCR#0ERICHMRFN_lORsFHH#RMN#0MN0H03C8
HS#oDMNS8bNF,CMR8bNF,k0R8bNH:MSS8#0_oDFH
O;S#
SHNoMDHSbML_OHS0:#_08DHFoOC_POs0F586RF0IMF2Rj;#
SHNoMDCSMos_0HSo:#_08DHFoOS;

-S-SlOFbCFMMb0RsHC_FO
SFFlbM0CMSCbs_
HFSsbF0
S5SESSFSD8:MSHR0S#8F_Do;HO
SSSsH#0FSS:H#MS0D8_FOoH;S
SS_L#C:MSSSHM#_08DHFoOS;
SES#HSV0:MSHS8#0_oDFH
O;S0SSOSD	:MSHS8#0_oDFH
O;SHSSM	ODSH:SM0S#8F_Do;HO
SSSFOk0D:	SSSHM#_08DHFoOS;
SbSk8CN0SH:SM0S#8F_Do;HO
SSSFHCbMSS:H#MS0D8_FOoH;S
SSH#8SSS:H#MS0D8_FOoH;S
SS8lFCSS:H#MS0D8_FOoH;S
SSxEH_:LSSSHM#_08DHFoOS;
S8S#F:SSS0FkS8#0_oDFH
O;S8SSF4k0SF:Sk#0S0D8_FOoH;S
SSk8F0:jSS0FkS8#0_oDFH
O;S8SS8Ss4:MSHS8#0_oDFH
O;S8SS8Ssj:MSHS8#0_oDFH
O;SbSSNM8HSH:SM0S#8F_Do;HO
SSSbFN8k:0SS0FkS8#0_oDFH
O;SbSSNC8FMSS:FSk0#_08DHFoOS;
SLSOH:0SSSHM#_08DHFoOC_POs0FSR568MFI0jFR2S
SS
2;S8CMRlOFbCFMM
0;
oLCHSM
M_Co0osHSS<=a1m_am7ptSQB5th _Qa)t)t 2S;
b_HMO0LHSS<=a1m_am7pteQB mBa)uS5Qah_Y2u ;

S
MSHO_D	M=S<RhSQu_zaBRpiGRFsM_Co0osH;F
SkD0O	S_M<m=Szzauap_BiFRGsCRMos_0H
o;SOHMD<	S=MSHO_D	MMRN8pRBm_Bi Ahqp
 ;S0FkOSD	<F=SkD0O	R_MNRM8BBpmih_ q Ap;

SSDEF8=S<SapqBQ]_hauz_peqz
 ;SbFCH<MS=zSmaauz_q hA;p 
SS
uiqBq_t u_QhHSS:bOsFCS##58bNF,CMR8bNF2k0
CSLo
HMSVSHSN5b8MFC=''42ER0CSM
SqSuBtiq Q_uh=S<S''Z;S
SCCD#
SSSuiqBq_t uSQh<b=SNk8F0S;
S8CMR;HV
MSC8sRbF#OC#S;

NSb8RHM<u=RqqBitu _Q;hR
SS
uiqBq_t u_QhAS_H:sSbF#OC#bS5NC8FMb,RNk8F0S2
LHCoMS
SH5VSbFN8C'M=4R'20MEC
SSSuiqBq_t u_QhA=S<S''Z;S
SCCD#
SSSuiqBq_t u_QhA=S<S0MFR8bNF;k0
CSSMH8RVS;
CRM8bOsFC;##
E
SFSD8<p=Rq]aB_uQhzea_q pz;F
SCMbHR=S<Ramzu_za Ahqp
 ;
S--b_sCHHF_
sSbCF_H_:HSSCbs_
HFSsbF0NRlb
S5SSSSE8FDSS=>E8FD,S
SS#Ss0SHF='>Sj
',SSSSLC#_M>S=S_L#C
M,SSSS#VEH0>S=SH#EV
0,SSSS0	ODSS=>0	OD,S
SSMSHOSD	=H>SM	OD,S
SSkSF0	ODSS=>FOk0D
	,SSSSkNb80=CS>bSk8CN0,S
SSCSFbSHM=F>SCMbH,S
SS8S#H=SS>8S#HS,
SlSSFS8C=l>SF,8C
SSSSxEH_=LS>HSEx,_L
SSSSF#8S>S=SF#8,S
SSFS8kS04=7>S__Qh4S,
S8SSFjk0SS=>7h_Q_
j,SSSS848sSS=>7z_ma,_4
SSSSs88j>S=Sm7_zja_,S
SSNSb8SHM=b>SNM8H,S
SSNSb80FkSS=>bFN8k
0,SSSSbFN8C=MS>NSb8MFC,S
SSLSOH=0S>HSbML_OHS0
S2SS;C

M18RAm_Q__71e
;
--------------------------------------------------------------
-SSSSS7th
------------------------------------------------------------
-
DsHLNRs$HCCC;#
kCCRHC#C30D8_FOoH_n44cD3NDk;
#HCRC3CC#_08DHFoOs_NH30EN;DD
Ck#RCHCC03#8F_Do_HOkHM#o8MC3DND;C

M00H$hSt7#SH
sbF0
S5SSSY:kSF00S#8F_Do
HOS;S2
M
C8hRt7N;
0H0sLCk0RM#$_NLDOL	_FFGRVhRt7RR:ObFlFMMC0#RHRk0sC
;
NEsOHO0C0CksR7th_FeRVhRt7#RH
oLCHSM
Y=S<S''j;M
C8hRt7;_e
-
----------------------------------------------------------
---S-SSeSSB-B
------------------------------------------------------------
H
DLssN$CRHC
C;kR#CHCCC38#0_oDFH4O_43ncN;DD
Ck#RCHCC03#8F_Do_HON0sHED3NDk;
#HCRC3CC#_08DHFoOM_k#MHoCN83D
D;
0CMHS0$eSBBHb#
FSs05S
SYSS:FSk0#_08DHFoOS
S2
;
CRM8e;BB
0N0skHL0#CR$LM_D	NO_GLFRRFVeRBB:FROlMbFCRM0H0#Rs;kC
s
NO0EHCkO0seCRBeB_RRFVeRBBHL#
CMoH
SSY<'=S4
';CRM8e_BBe
;

-
-/////////////////////////////////////-R---
S-Q-RBj cv)]RquvRsHHl0CHP#-R---
-/////////////////////////////////////-R--


-------------------------------------
--S---R_1A)4qvjG.c4-n
-------------------------------------D-
HNLssQ$R ;  
Ck#R Q  a317m_pt_QB4c4n3DND;#
kC RQ 1 3ap7_mBtQ_1zhQ th7D3NDk;
#QCR 3  #_08DHFoOs_NH30EN;DD
 z1R Q  k3MlHCsO0_#8p3qp
;
CHM001$RAq_)v.4jcnX4R
H#
oRRCsMCH5ORRR
RRRRRRRRRRQQhaR_j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QanRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ(a_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QaqRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQAa_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQwa_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R

RRRRRRRRRhRQQ4a_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;R
RRRRRRRRRRRQahQ_R.j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R..:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R. :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"RR

RRRRRRRRRhRQQda_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"RR
RRRRRRRRR2RRR
;
RRRRRRRRRFRbsR05
RRRRRRRRRRRRRRRRq)7a:qRR0FkR8#0_oDFHPO_CFO0s45R68RRF0IMF2RjRR;
RRRRRRRRRRRRR)RRBRpiRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRR)RRB piRH:RM#RR0D8_FOoHRR:=';]'
RRRRRRRRRRRRRRRRR) R:RRRRHMR8#0_oDFH:OR=]R''R;
RRRRRRRRRRRRR)RRq)77RH:RM#RR0D8_FOoH_OPC05FsRRgR8MFI0jFR2
R;RRRRRRRRRRRRRRRRWiBpRRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRRWiBp RR:HRMR#_08DHFoO=R:R''];R
RRRRRRRRRRRRRR RWRRRR:MRHR0R#8F_DoRHO:'=R]
';RRRRRRRRRRRRRRRRW7q7)RR:HRMR#_08DHFoOC_POs0F5RRgRI8FMR0Fj;2R
RRRRRRRRRRRRRRRR1vqi:RRRRHMR8#0_oDFHPO_CFO0s45R68RRF0IMF2RjRR;
RRRRRRRRRRRRRWRR7qqaRH:RM#RR0D8_FOoH_OPC05FsRR46RI8FMR0FjR2
RRRRRRRRRRRRR;R2

RRRCR
M18RAq_)v.4jcnX4;N

sHOE00COkRsC1)A_qjv4.4cXn)_qBF]RVAR1_v)q4cj.XR4nHL#
CMoHRM
C8AR1_v)q4cj.X_4nq])B;RRR-R--1)A_qjv4.4cXn


-------------------------------------
--S---R_1A)4qvjG.c4)nh
---------------------------------------
LDHs$NsR Q  k;
#QCR 3  1_a7pQmtB4_4nNc3D
D;kR#CQ   371a_tpmQzB_ht1Qh3 7N;DD
Ck#R Q  03#8F_Do_HON0sHED3NDz;
1Q R 3  MCkls_HO#308q;pp
M
C0$H0R_1A)4qvjG.c4)nhR
H#
oRRCsMCH5ORRR
RRRRRRRRRRQQhaR_j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QanRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ(a_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QaqRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQAa_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQwa_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;
R
RRRRRRRRRQRRh_Qa4:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjR";
R
RRRRRRRRRRQQhaj_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha4_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha._.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhad_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhac_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha6_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhan_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha(_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaU_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhag_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaq_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaA_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaB_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha7_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha _.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaw_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;
R
RRRRRRRRRQRRh_Qad:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
"RRRRRRRRRRRRR2
R;RRRRRRRRRFRbsR05
RRRRRRRRRRRRRRRRq)7a:qRR0FkR8#0_oDFHPO_CFO0s45R68RRF0IMF2RjRR;
RRRRRRRRRRRRR)RRBhpiRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRR)RRB piRH:RM#RR0D8_FOoHRR:=';]'
RRRRRRRRRRRRRRRRR) R:RRRRHMR8#0_oDFH:OR=]R''R;
RRRRRRRRRRRRR)RRq)77RH:RM#RR0D8_FOoH_OPC05FsRRgR8MFI0jFR2
R;RRRRRRRRRRRRRRRRWiBpRRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRRWiBp RR:HRMR#_08DHFoO=R:R''];R
RRRRRRRRRRRRRR RWRRRR:MRHR0R#8F_DoRHO:'=R]
';RRRRRRRRRRRRRRRRW7q7)RR:HRMR#_08DHFoOC_POs0F5RRgRI8FMR0Fj;2R
RRRRRRRRRRRRRRRR1vqi:RRRRHMR8#0_oDFHPO_CFO0s45R68RRF0IMF2RjRR;
RRRRRRRRRRRRRWRR7qqaRH:RM#RR0D8_FOoH_OPC05FsRR46RI8FMR0FjR2
RRRRRRRRRRRRR;R2

RRRCR
M18RAq_)v.4jcnG4h
);
ONsECH0Os0kCAR1_v)q4cj.Gh4n))_qBF]RVAR1_v)q4cj.Gh4n)#RH
oLCH
MRCRM81)A_qjv4.4cGn_h)q])B;RRR-R--1)A_qjv4.4cGn
h)
-
---------------------------------------
S-1-RAq_)v.4jcnG4h-W
-------------------------------------D-
HNLssQ$R ;  
Ck#R Q  a317m_pt_QB4c4n3DND;#
kC RQ 1 3ap7_mBtQ_1zhQ th7D3NDk;
#QCR 3  #_08DHFoOs_NH30EN;DD
 z1R Q  k3MlHCsO0_#8p3qp
;
CHM001$RAq_)v.4jcnG4hHWR#R

RMoCCOsHR
5RRRRRRRRRRQRRh_QajRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QacRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ6a_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QaURR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQga_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QaBRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ7a_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_ :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RRRRRRRRRRRQahQ_R4j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R44:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R46:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R47:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4 :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
RRRRRRRRRRQQhaj_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha4_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha._.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhad_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhac_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha6_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhan_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha(_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaU_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhag_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaq_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaA_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaB_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha7_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha _.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaw_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R

RRRRRRRRRhRQQda_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"RR
RRRRRRRRR2RRRR;
RRRRRRRRRsbF0
5RRRRRRRRRRRRRRRRR)a7qqRR:FRk0#_08DHFoOC_POs0F56R4RFR8IFM0RRj2;R
RRRRRRRRRRRRRRBR)pRiR:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRBR)pRi :MRHR0R#8F_DoRHO:'=R]
';RRRRRRRRRRRRRRRR)R RRRR:HRMR#_08DHFoO=R:R''];R
RRRRRRRRRRRRRRqR)7R7):MRHR0R#8F_Do_HOP0COFRs5g8RRF0IMF2RjRR;
RRRRRRRRRRRRRWRRBhpiRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRRWRRB piRH:RM#RR0D8_FOoHRR:=';]'
RRRRRRRRRRRRRRRRRW R:RRRRHMR8#0_oDFH:OR=]R''R;
RRRRRRRRRRRRRWRRq)77RH:RM#RR0D8_FOoH_OPC05FsRRgR8MFI0jFR2
R;RRRRRRRRRRRRRRRRviq1RRR:HRMR#_08DHFoOC_POs0F56R4RFR8IFM0RRj2;R
RRRRRRRRRRRRRR7RWqRaq:MRHR0R#8F_Do_HOP0COFRs54R6R8MFI0jFR2R
RRRRRRRRRRRRRR
2;RRR
RM
C8AR1_v)q4cj.Gh4nW
;
NEsOHO0C0CksR_1A)4qvjG.c4Wnh_Bq)]VRFR_1A)4qvjG.c4WnhR
H#LHCoMCR
M18RAq_)v.4jcnG4hqW_);B]R-RR-1-RAq_)v.4jcnG4h
W

-
---------------------------------------
S-1-RAq_)v.4jcnG4hW)h
---------------------------------------
LDHs$NsR Q  k;
#QCR 3  1_a7pQmtB4_4nNc3D
D;kR#CQ   371a_tpmQzB_ht1Qh3 7N;DD
Ck#R Q  03#8F_Do_HON0sHED3NDz;
1Q R 3  MCkls_HO#308q;pp
M
C0$H0R_1A)4qvjG.c4)nhhHWR#R

RMoCCOsHR
5RRRRRRRRRRQRRh_QajRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QacRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ6a_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QaURR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQga_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QaBRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ7a_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_ :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RRRRRRRRRRRQahQ_R4j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R44:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R46:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R47:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4 :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
RRRRRRRRRRQQhaj_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha4_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha._.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhad_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhac_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha6_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhan_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha(_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaU_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhag_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaq_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaA_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaB_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha7_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha _.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaw_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R

RRRRRRRRRhRQQda_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"RR
RRRRRRRRR2RRRR;
RRRRRRRRRsbF0
5RRRRRRRRRRRRRRRRR)a7qqRR:FRk0#_08DHFoOC_POs0F56R4RFR8IFM0RRj2;R
RRRRRRRRRRRRRRBR)pRih:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRBR)pRi :MRHR0R#8F_DoRHO:'=R]
';RRRRRRRRRRRRRRRR)R RRRR:HRMR#_08DHFoO=R:R''];R
RRRRRRRRRRRRRRqR)7R7):MRHR0R#8F_Do_HOP0COFRs5g8RRF0IMF2RjRR;
RRRRRRRRRRRRRWRRBhpiRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRRWRRB piRH:RM#RR0D8_FOoHRR:=';]'
RRRRRRRRRRRRRRRRRW R:RRRRHMR8#0_oDFH:OR=]R''R;
RRRRRRRRRRRRRWRRq)77RH:RM#RR0D8_FOoH_OPC05FsRRgR8MFI0jFR2
R;RRRRRRRRRRRRRRRRviq1RRR:HRMR#_08DHFoOC_POs0F56R4RFR8IFM0RRj2;R
RRRRRRRRRRRRRR7RWqRaq:MRHR0R#8F_Do_HOP0COFRs54R6R8MFI0jFR2R
RRRRRRRRRRRRRR
2;RRR
RM
C8AR1_v)q4cj.Gh4n);hW
s
NO0EHCkO0s1CRAq_)v.4jcnG4hW)h_Bq)]VRFR_1A)4qvjG.c4)nhhHWR#C
LoRHM
8CMR_1A)4qvjG.c4)nhhqW_);B]R-RR-1-RAq_)v.4jcnG4hW)h
-

-------------------------------------S-
-R--1)A_qjv.cUUG
---------------------------------------
LDHs$NsR Q  k;
#QCR 3  1_a7pQmtB4_4nNc3D
D;kR#CQ   371a_tpmQzB_ht1Qh3 7N;DD
Ck#R Q  03#8F_Do_HON0sHED3NDz;
1Q R 3  MCkls_HO#308q;pp
M
C0$H0R_1A).qvjGcUU#RH
R
RoCCMsRHO5RR
RRRRRRRRRhRQQja_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QadRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQca_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQUa_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QaARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQBa_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QawRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
RRRRRRRRRQRRh_Qa4:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RRRRRRRRRRRQahQ_R.j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R..:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R. :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
RRRRRRRRRRQQhaj_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha4_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha._dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhad_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhac_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha6_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhan_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha(_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaU_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhag_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaq_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaA_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaB_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha7_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha _dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaw_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jjRR
RRRRRRRRRRRR2;R
RRRRRRRRRb0Fs5RR
RRRRRRRRRRRRR)RR7qqaRF:Rk#0R0D8_FOoH_OPC05FsRR(R8MFI0jFR2
R;RRRRRRRRRRRRRRRR)iBpRRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRR)iBp RR:HRMR#_08DHFoO=R:R''];R
RRRRRRRRRRRRRR R)RRRR:MRHR0R#8F_DoRHO:'=R]
';RRRRRRRRRRRRRRRR)7q7)RR:HRMR#_08DHFoOC_POs0F5jR4RFR8IFM0RRj2;R
RRRRRRRRRRRRRRBRWpRiR:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRBRWpRi :MRHR0R#8F_DoRHO:'=R]
';RRRRRRRRRRRRRRRRWR RRRR:HRMR#_08DHFoO=R:R''];R
RRRRRRRRRRRRRRqRW7R7):MRHR0R#8F_Do_HOP0COFRs54RjR8MFI0jFR2
R;RRRRRRRRRRRRRRRRWa7qqRR:HRMR#_08DHFoOC_POs0F5RR(RI8FMR0FjR2
RRRRRRRRRRRRR;R2

RRRCR
M18RAq_)vc.jU;GU
s
NO0EHCkO0s1CRAq_)vc.jU_GUq])BRRFV1)A_qjv.cUUGR
H#LHCoMCR
M18RAq_)vc.jU_GUq])B;RRR-R--1)A_qjv.cUUG



-------------------------------------
--S---R_1A).qvjGcUU
h)-------------------------------------
--DsHLNRs$Q   ;#
kC RQ 1 3ap7_mBtQ_n44cD3NDk;
#QCR 3  1_a7pQmtBh_z1hQt N73D
D;kR#CQ   38#0_oDFHNO_sEH03DND;1
z  RQ M 3kslCH#O_0q83p
p;
0CMHR0$1)A_qjv.cUUGhH)R#R

RMoCCOsHR
5RRRRRRRRRRQRRh_QajRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QacRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ6a_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QaURR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQga_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QaBRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ7a_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_ :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RRRRRRRRRRRQahQ_R4j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R44:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R46:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R47:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4 :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
RRRRRRRRRRQQhaj_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha4_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha._.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhad_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhac_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha6_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhan_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha(_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaU_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhag_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaq_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaA_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaB_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha7_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha _.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaw_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R

RRRRRRRRRhRQQda_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"RR
RRRRRRRRR2RRRR;
RRRRRRRRRsbF0
5RRRRRRRRRRRRRRRRR)a7qqRR:FRk0#_08DHFoOC_POs0F5RR(RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRp)Bi:hRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRp)Bi: RRRHMR8#0_oDFH:OR=]R''R;
RRRRRRRRRRRRR)RR RRRRH:RM#RR0D8_FOoHRR:=';]'
RRRRRRRRRRRRRRRR7)q7:)RRRHMR8#0_oDFHPO_CFO0s45Rj8RRF0IMF2RjRR;
RRRRRRRRRRRRRWRRBRpiRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRRWRRB piRH:RM#RR0D8_FOoHRR:=';]'
RRRRRRRRRRRRRRRRRW R:RRRRHMR8#0_oDFH:OR=]R''R;
RRRRRRRRRRRRRWRRq)77RH:RM#RR0D8_FOoH_OPC05FsRR4jRI8FMR0Fj;2R
RRRRRRRRRRRRRRRRqW7a:qRRRHMR8#0_oDFHPO_CFO0s(5RRFR8IFM0R
j2RRRRRRRRRRRRR2RR;R
R

RRCRM81)A_qjv.cUUGh
);
ONsECH0Os0kCAR1_v)q.UjcG)Uh_Bq)]VRFR_1A).qvjGcUURh)HL#
CMoHRM
C8AR1_v)q.UjcG)Uh_Bq)]R;RR---R_1A).qvjGcUU
h)
-

-------------------------------------S-
-R--1)A_qjv.cUUGh-W
-------------------------------------D-
HNLssQ$R ;  
Ck#R Q  a317m_pt_QB4c4n3DND;#
kC RQ 1 3ap7_mBtQ_1zhQ th7D3NDk;
#QCR 3  #_08DHFoOs_NH30EN;DD
 z1R Q  k3MlHCsO0_#8p3qp
;
CHM001$RAq_)vc.jUhGUW#RH
R
RoCCMsRHO5RR
RRRRRRRRRhRQQja_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QadRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQca_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQUa_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QaARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQBa_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QawRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
RRRRRRRRRQRRh_Qa4:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RRRRRRRRRRRQahQ_R.j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R..:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R. :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"RR

RRRRRRRRRhRQQda_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"RR
RRRRRRRRR2RRRR;
RRRRRRRRRsbF0
5RRRRRRRRRRRRRRRRR)a7qqRR:FRk0#_08DHFoOC_POs0F5RR(RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRp)Bi:RRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRp)Bi: RRRHMR8#0_oDFH:OR=]R''R;
RRRRRRRRRRRRR)RR RRRRH:RM#RR0D8_FOoHRR:=';]'
RRRRRRRRRRRRRRRR7)q7:)RRRHMR8#0_oDFHPO_CFO0s45Rj8RRF0IMF2RjRR;
RRRRRRRRRRRRRWRRBhpiRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRRWRRB piRH:RM#RR0D8_FOoHRR:=';]'
RRRRRRRRRRRRRRRRRW R:RRRRHMR8#0_oDFH:OR=]R''R;
RRRRRRRRRRRRRWRRq)77RH:RM#RR0D8_FOoH_OPC05FsRR4jRI8FMR0Fj;2R
RRRRRRRRRRRRRRRRqW7a:qRRRHMR8#0_oDFHPO_CFO0s(5RRFR8IFM0R
j2RRRRRRRRRRRRR2RR;R
R

RRCRM81)A_qjv.cUUGh
W;
ONsECH0Os0kCAR1_v)q.UjcGWUh_Bq)]VRFR_1A).qvjGcUURhWHL#
CMoHRM
C8AR1_v)q.UjcGWUh_Bq)]R;RR---R_1A).qvjGcUU
hW
-
---------------------------------------
S-1-RAq_)vc.jUhGU)
hW-------------------------------------
--DsHLNRs$Q   ;#
kC RQ 1 3ap7_mBtQ_n44cD3NDk;
#QCR 3  1_a7pQmtBh_z1hQt N73D
D;kR#CQ   38#0_oDFHNO_sEH03DND;1
z  RQ M 3kslCH#O_0q83p
p;
0CMHR0$1)A_qjv.cUUGhW)hR
H#
oRRCsMCH5ORRR
RRRRRRRRRRQQhaR_j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QanRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ(a_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QaqRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQAa_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQwa_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;
R
RRRRRRRRRQRRh_Qa4:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjR";
R
RRRRRRRRRRQQhaj_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha4_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha._.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhad_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhac_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha6_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhan_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha(_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaU_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhag_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaq_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaA_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaB_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha7_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha _.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaw_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;
R
RRRRRRRRRQRRh_Qad:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
"RRRRRRRRRRRRR2
R;RRRRRRRRRFRbsR05
RRRRRRRRRRRRRRRRq)7a:qRR0FkR8#0_oDFHPO_CFO0s(5RRFR8IFM0RRj2;R
RRRRRRRRRRRRRRBR)pRih:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRBR)pRi :MRHR0R#8F_DoRHO:'=R]
';RRRRRRRRRRRRRRRR)R RRRR:HRMR#_08DHFoO=R:R''];R
RRRRRRRRRRRRRRqR)7R7):MRHR0R#8F_Do_HOP0COFRs54RjR8MFI0jFR2
R;RRRRRRRRRRRRRRRRWiBphRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRRWiBp RR:HRMR#_08DHFoO=R:R''];R
RRRRRRRRRRRRRR RWRRRR:MRHR0R#8F_DoRHO:'=R]
';RRRRRRRRRRRRRRRRW7q7)RR:HRMR#_08DHFoOC_POs0F5jR4RFR8IFM0RRj2;R
RRRRRRRRRRRRRR7RWqRaq:MRHR0R#8F_Do_HOP0COFRs5(8RRF0IMF2Rj
RRRRRRRRRRRRRRR2R;
RR
R
8CMR_1A).qvjGcUUhh)W
;
NEsOHO0C0CksR_1A).qvjGcUUhh)W)_qBF]RVAR1_v)q.UjcG)UhhHWR#C
LoRHM
8CMR_1A).qvjGcUUhh)W)_qBR];R-R--AR1_v)q.UjcG)Uhh
W

---------------------------------------
-S--AR1_v)qcnjgG-c
-------------------------------------D-
HNLssQ$R ;  
Ck#R Q  a317m_pt_QB4c4n3DND;#
kC RQ 1 3ap7_mBtQ_1zhQ th7D3NDk;
#QCR 3  #_08DHFoOs_NH30EN;DD
 z1R Q  k3MlHCsO0_#8p3qp
;
CHM001$RAq_)vgcjnRGcH
#
RCRoMHCsORR5
RRRRRRRRRRRQahQ_:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQna_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QagRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQqa_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ a_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"RR

RRRRRRRRRhRQQ4a_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;R
RRRRRRRRRRRQahQ_R.j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R..:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R. :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"RR

RRRRRRRRRhRQQda_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"RR
RRRRRRRRR2RRRR;
RRRRRRRRRsbF0
5RRRRRRRRRRRRRRRRR)a7qqRR:FRk0#_08DHFoOC_POs0F5RRdRI8FMR0Fj;2R
RRRRRRRRRRRRRRRRp)Bi:RRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRp)Bi: RRRHMR8#0_oDFH:OR=]R''R;
RRRRRRRRRRRRR)RR RRRRH:RM#RR0D8_FOoHRR:=';]'
RRRRRRRRRRRRRRRR7)q7:)RRRHMR8#0_oDFHPO_CFO0s45R48RRF0IMF2RjRR;
RRRRRRRRRRRRRWRRBRpiRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRRWRRB piRH:RM#RR0D8_FOoHRR:=';]'
RRRRRRRRRRRRRRRRRW R:RRRRHMR8#0_oDFH:OR=]R''R;
RRRRRRRRRRRRRWRRq)77RH:RM#RR0D8_FOoH_OPC05FsRR44RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRqW7a:qRRRHMR8#0_oDFHPO_CFO0sd5RRFR8IFM0R
j2RRRRRRRRRRRRR2RR;R
R

RRCRM81)A_qjvcgcnG;N

sHOE00COkRsC1)A_qjvcgcnG_Bq)]VRFR_1A)cqvjGgnc#RH
oLCH
MRCRM81)A_qjvcgcnG_Bq)]R;RR---R_1A)cqvjGgnc



---------------------------------------
-S--AR1_v)qcnjgG)ch
---------------------------------------
LDHs$NsR Q  k;
#QCR 3  1_a7pQmtB4_4nNc3D
D;kR#CQ   371a_tpmQzB_ht1Qh3 7N;DD
Ck#R Q  03#8F_Do_HON0sHED3NDz;
1Q R 3  MCkls_HO#308q;pp
M
C0$H0R_1A)cqvjGgncRh)H
#
RCRoMHCsORR5
RRRRRRRRRRRQahQ_:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQna_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QagRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQqa_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ a_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"RR

RRRRRRRRRhRQQ4a_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;R
RRRRRRRRRRRQahQ_R.j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R..:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R. :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"RR

RRRRRRRRRhRQQda_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"RR
RRRRRRRRR2RRRR;
RRRRRRRRRsbF0
5RRRRRRRRRRRRRRRRR)a7qqRR:FRk0#_08DHFoOC_POs0F5RRdRI8FMR0Fj;2R
RRRRRRRRRRRRRRRRp)Bi:hRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRp)Bi: RRRHMR8#0_oDFH:OR=]R''R;
RRRRRRRRRRRRR)RR RRRRH:RM#RR0D8_FOoHRR:=';]'
RRRRRRRRRRRRRRRR7)q7:)RRRHMR8#0_oDFHPO_CFO0s45R48RRF0IMF2RjRR;
RRRRRRRRRRRRRWRRBRpiRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRRWRRB piRH:RM#RR0D8_FOoHRR:=';]'
RRRRRRRRRRRRRRRRRW R:RRRRHMR8#0_oDFH:OR=]R''R;
RRRRRRRRRRRRRWRRq)77RH:RM#RR0D8_FOoH_OPC05FsRR44RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRqW7a:qRRRHMR8#0_oDFHPO_CFO0sd5RRFR8IFM0R
j2RRRRRRRRRRRRR2RR;R
R

RRCRM81)A_qjvcgcnGh
);
ONsECH0Os0kCAR1_v)qcnjgG)ch_Bq)]VRFR_1A)cqvjGgncRh)HL#
CMoHRM
C8AR1_v)qcnjgG)ch_Bq)]R;RR---R_1A)cqvjGgnc
h)
-
---------------------------------------
S-1-RAq_)vgcjnhGcW-
--------------------------------------H
DLssN$ RQ 
 ;kR#CQ   371a_tpmQ4B_43ncN;DD
Ck#R Q  a317m_pt_QBzQh1t7h 3DND;#
kC RQ # 30D8_FOoH_HNs0NE3D
D;zR1 Q   3lMkCOsH_8#03pqp;C

M00H$AR1_v)qcnjgGWchR
H#
oRRCsMCH5ORRR
RRRRRRRRRRQQhaR_j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QanRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ(a_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QaqRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQAa_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQwa_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;
R
RRRRRRRRRQRRh_Qa4:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjR";
R
RRRRRRRRRRQQhaj_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha4_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha._.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhad_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhac_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha6_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhan_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha(_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaU_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhag_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaq_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaA_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaB_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha7_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha _.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaw_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;
R
RRRRRRRRRQRRh_Qad:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
"RRRRRRRRRRRRR2
R;RRRRRRRRRFRbsR05
RRRRRRRRRRRRRRRRq)7a:qRR0FkR8#0_oDFHPO_CFO0sd5RRFR8IFM0RRj2;R
RRRRRRRRRRRRRRBR)pRiR:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRBR)pRi :MRHR0R#8F_DoRHO:'=R]
';RRRRRRRRRRRRRRRR)R RRRR:HRMR#_08DHFoO=R:R''];R
RRRRRRRRRRRRRRqR)7R7):MRHR0R#8F_Do_HOP0COFRs54R4R8MFI0jFR2
R;RRRRRRRRRRRRRRRRWiBphRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRRWiBp RR:HRMR#_08DHFoO=R:R''];R
RRRRRRRRRRRRRR RWRRRR:MRHR0R#8F_DoRHO:'=R]
';RRRRRRRRRRRRRRRRW7q7)RR:HRMR#_08DHFoOC_POs0F54R4RFR8IFM0RRj2;R
RRRRRRRRRRRRRR7RWqRaq:MRHR0R#8F_Do_HOP0COFRs5d8RRF0IMF2Rj
RRRRRRRRRRRRRRR2R;
RR
R
8CMR_1A)cqvjGgnc;hW
s
NO0EHCkO0s1CRAq_)vgcjnhGcW)_qBF]RVAR1_v)qcnjgGWchR
H#LHCoMCR
M18RAq_)vgcjnhGcW)_qBR];R-R--AR1_v)qcnjgGWch
-

-------------------------------------S-
-R--1)A_qjvcgcnGhW)h
---------------------------------------
LDHs$NsR Q  k;
#QCR 3  1_a7pQmtB4_4nNc3D
D;kR#CQ   371a_tpmQzB_ht1Qh3 7N;DD
Ck#R Q  03#8F_Do_HON0sHED3NDz;
1Q R 3  MCkls_HO#308q;pp
M
C0$H0R_1A)cqvjGgnchh)W#RH
R
RoCCMsRHO5RR
RRRRRRRRRhRQQja_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QadRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQca_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQUa_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QaARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQBa_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QawRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;R
RRRRRRRRRRRQahQ_R4j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R44:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R46:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R47:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4 :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"RR

RRRRRRRRRhRQQ.a_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;R
RRRRRRRRRRRQahQ_Rdj:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_Rd4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_Rd.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_Rdd:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_Rdc:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_Rd6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_Rdn:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_Rd(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_RdU:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_Rdg:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_Rdq:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_RdA:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_RdB:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_Rd7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_Rd :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_Rdw:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjRj"
RRRRRRRRRRRR;2R
RRRRRRRRbRRF5s0RR
RRRRRRRRRRRRRR7R)qRaq:kRF00R#8F_Do_HOP0COFRs5d8RRF0IMF2RjRR;
RRRRRRRRRRRRR)RRBhpiRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRR)RRB piRH:RM#RR0D8_FOoHRR:=';]'
RRRRRRRRRRRRRRRRR) R:RRRRHMR8#0_oDFH:OR=]R''R;
RRRRRRRRRRRRR)RRq)77RH:RM#RR0D8_FOoH_OPC05FsRR44RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRpWBi:hRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRpWBi: RRRHMR8#0_oDFH:OR=]R''R;
RRRRRRRRRRRRRWRR RRRRH:RM#RR0D8_FOoHRR:=';]'
RRRRRRRRRRRRRRRR7Wq7:)RRRHMR8#0_oDFHPO_CFO0s45R48RRF0IMF2RjRR;
RRRRRRRRRRRRRWRR7qqaRH:RM#RR0D8_FOoH_OPC05FsRRdR8MFI0jFR2R
RRRRRRRRRRRRRR
2;RRR
RM
C8AR1_v)qcnjgG)chh
W;
ONsECH0Os0kCAR1_v)qcnjgG)chhqW_)RB]F1VRAq_)vgcjnhGc)RhWHL#
CMoHRM
C8AR1_v)qcnjgG)chhqW_);B]R-RR-1-RAq_)vgcjnhGc)
hW
-
---------------------------------------
S-1-RAq_)vgU4.
G.-------------------------------------
--DsHLNRs$Q   ;#
kC RQ 1 3ap7_mBtQ_n44cD3NDk;
#QCR 3  1_a7pQmtBh_z1hQt N73D
D;kR#CQ   38#0_oDFHNO_sEH03DND;1
z  RQ M 3kslCH#O_0q83p
p;
0CMHR0$1)A_q4vUg..GR
H#
oRRCsMCH5ORRR
RRRRRRRRRRQQhaR_j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QanRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ(a_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QaqRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQAa_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQwa_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;
R
RRRRRRRRRQRRh_Qa4:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjR";
R
RRRRRRRRRRQQhaj_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha4_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha._.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhad_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhac_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha6_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhan_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha(_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaU_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhag_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaq_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaA_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaB_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha7_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha _.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaw_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;
R
RRRRRRRRRQRRh_Qad:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
"RRRRRRRRRRRRR2
R;RRRRRRRRRFRbsR05
RRRRRRRRRRRRRRRRq)7a:qRR0FkR8#0_oDFHPO_CFO0s45RRFR8IFM0RRj2;R
RRRRRRRRRRRRRRBR)pRiR:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRBR)pRi :MRHR0R#8F_DoRHO:'=R]
';RRRRRRRRRRRRRRRR)R RRRR:HRMR#_08DHFoO=R:R''];R
RRRRRRRRRRRRRRqR)7R7):MRHR0R#8F_Do_HOP0COFRs54R.R8MFI0jFR2
R;RRRRRRRRRRRRRRRRWiBpRRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRRWiBp RR:HRMR#_08DHFoO=R:R''];R
RRRRRRRRRRRRRR RWRRRR:MRHR0R#8F_DoRHO:'=R]
';RRRRRRRRRRRRRRRRW7q7)RR:HRMR#_08DHFoOC_POs0F5.R4RFR8IFM0RRj2;R
RRRRRRRRRRRRRR7RWqRaq:MRHR0R#8F_Do_HOP0COFRs548RRF0IMF2Rj
RRRRRRRRRRRRRRR2R;
RR
R
8CMR_1A)Uqv4Gg..
;
NEsOHO0C0CksR_1A)Uqv4Gg..)_qBF]RVAR1_v)qU.4gGH.R#C
LoRHM
8CMR_1A)Uqv4Gg..)_qBR];R-R--AR1_v)qU.4gG
.

---------------------------------------
-S--AR1_v)qU.4gG).h
---------------------------------------
LDHs$NsR Q  k;
#QCR 3  1_a7pQmtB4_4nNc3D
D;kR#CQ   371a_tpmQzB_ht1Qh3 7N;DD
Ck#R Q  03#8F_Do_HON0sHED3NDz;
1Q R 3  MCkls_HO#308q;pp
M
C0$H0R_1A)Uqv4Gg..Rh)H
#
RCRoMHCsORR5
RRRRRRRRRRRQahQ_:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQna_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QagRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQqa_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ a_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"RR

RRRRRRRRRhRQQ4a_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;R
RRRRRRRRRRRQahQ_R.j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R..:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R. :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"RR

RRRRRRRRRhRQQda_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"RR
RRRRRRRRR2RRRR;
RRRRRRRRRsbF0
5RRRRRRRRRRRRRRRRR)a7qqRR:FRk0#_08DHFoOC_POs0F5RR4RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRp)Bi:hRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRp)Bi: RRRHMR8#0_oDFH:OR=]R''R;
RRRRRRRRRRRRR)RR RRRRH:RM#RR0D8_FOoHRR:=';]'
RRRRRRRRRRRRRRRR7)q7:)RRRHMR8#0_oDFHPO_CFO0s45R.8RRF0IMF2RjRR;
RRRRRRRRRRRRRWRRBRpiRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRRWRRB piRH:RM#RR0D8_FOoHRR:=';]'
RRRRRRRRRRRRRRRRRW R:RRRRHMR8#0_oDFH:OR=]R''R;
RRRRRRRRRRRRRWRRq)77RH:RM#RR0D8_FOoH_OPC05FsRR4.RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRqW7a:qRRRHMR8#0_oDFHPO_CFO0s45RRFR8IFM0R
j2RRRRRRRRRRRRR2RR;R
R

RRCRM81)A_q4vUg..Gh
);
ONsECH0Os0kCAR1_v)qU.4gG).h_Bq)]VRFR_1A)Uqv4Gg..Rh)HL#
CMoHRM
C8AR1_v)qU.4gG).h_Bq)]R;RR---R_1A)Uqv4Gg..
h)
-
---------------------------------------
S-1-RAq_)vgU4.hG.W-
--------------------------------------H
DLssN$ RQ 
 ;kR#CQ   371a_tpmQ4B_43ncN;DD
Ck#R Q  a317m_pt_QBzQh1t7h 3DND;#
kC RQ # 30D8_FOoH_HNs0NE3D
D;zR1 Q   3lMkCOsH_8#03pqp;C

M00H$AR1_v)qU.4gGW.hR
H#
oRRCsMCH5ORRR
RRRRRRRRRRQQhaR_j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QanRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ(a_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QaqRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQAa_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQwa_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;
R
RRRRRRRRRQRRh_Qa4:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjR";
R
RRRRRRRRRRQQhaj_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha4_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha._.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhad_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhac_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha6_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhan_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha(_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaU_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhag_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaq_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaA_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaB_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha7_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha _.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaw_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;
R
RRRRRRRRRQRRh_Qad:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
"RRRRRRRRRRRRR2
R;RRRRRRRRRFRbsR05
RRRRRRRRRRRRRRRRq)7a:qRR0FkR8#0_oDFHPO_CFO0s45RRFR8IFM0RRj2;R
RRRRRRRRRRRRRRBR)pRiR:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRBR)pRi :MRHR0R#8F_DoRHO:'=R]
';RRRRRRRRRRRRRRRR)R RRRR:HRMR#_08DHFoO=R:R''];R
RRRRRRRRRRRRRRqR)7R7):MRHR0R#8F_Do_HOP0COFRs54R.R8MFI0jFR2
R;RRRRRRRRRRRRRRRRWiBphRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRRWiBp RR:HRMR#_08DHFoO=R:R''];R
RRRRRRRRRRRRRR RWRRRR:MRHR0R#8F_DoRHO:'=R]
';RRRRRRRRRRRRRRRRW7q7)RR:HRMR#_08DHFoOC_POs0F5.R4RFR8IFM0RRj2;R
RRRRRRRRRRRRRR7RWqRaq:MRHR0R#8F_Do_HOP0COFRs548RRF0IMF2Rj
RRRRRRRRRRRRRRR2R;
RR
R
8CMR_1A)Uqv4Gg..;hW
s
NO0EHCkO0s1CRAq_)vgU4.hG.W)_qBF]RVAR1_v)qU.4gGW.hR
H#LHCoMCR
M18RAq_)vgU4.hG.W)_qBR];R-R--AR1_v)qU.4gGW.h
-

-------------------------------------S-
-R--1)A_q4vUg..GhW)h
---------------------------------------
LDHs$NsR Q  k;
#QCR 3  1_a7pQmtB4_4nNc3D
D;kR#CQ   371a_tpmQzB_ht1Qh3 7N;DD
Ck#R Q  03#8F_Do_HON0sHED3NDz;
1Q R 3  MCkls_HO#308q;pp
M
C0$H0R_1A)Uqv4Gg..hh)W#RH
R
RoCCMsRHO5RR
RRRRRRRRRhRQQja_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QadRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQca_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQUa_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QaARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQBa_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QawRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;R
RRRRRRRRRRRQahQ_R4j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R44:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R46:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R47:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4 :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"RR

RRRRRRRRRhRQQ.a_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;R
RRRRRRRRRRRQahQ_Rdj:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_Rd4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_Rd.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_Rdd:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_Rdc:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_Rd6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_Rdn:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_Rd(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_RdU:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_Rdg:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_Rdq:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_RdA:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_RdB:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_Rd7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_Rd :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_Rdw:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjRj"
RRRRRRRRRRRR;2R
RRRRRRRRbRRF5s0RR
RRRRRRRRRRRRRR7R)qRaq:kRF00R#8F_Do_HOP0COFRs548RRF0IMF2RjRR;
RRRRRRRRRRRRR)RRBhpiRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRR)RRB piRH:RM#RR0D8_FOoHRR:=';]'
RRRRRRRRRRRRRRRRR) R:RRRRHMR8#0_oDFH:OR=]R''R;
RRRRRRRRRRRRR)RRq)77RH:RM#RR0D8_FOoH_OPC05FsRR4.RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRpWBi:hRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRpWBi: RRRHMR8#0_oDFH:OR=]R''R;
RRRRRRRRRRRRRWRR RRRRH:RM#RR0D8_FOoHRR:=';]'
RRRRRRRRRRRRRRRR7Wq7:)RRRHMR8#0_oDFHPO_CFO0s45R.8RRF0IMF2RjRR;
RRRRRRRRRRRRRWRR7qqaRH:RM#RR0D8_FOoH_OPC05FsRR4R8MFI0jFR2R
RRRRRRRRRRRRRR
2;RRR
RM
C8AR1_v)qU.4gG).hh
W;
ONsECH0Os0kCAR1_v)qU.4gG).hhqW_)RB]F1VRAq_)vgU4.hG.)RhWHL#
CMoHRM
C8AR1_v)qU.4gG).hhqW_);B]R-RR-1-RAq_)vgU4.hG.)
hW
LDHs$NsR Q  k;
#QCR 3  1_a7pQmtB4_4nNc3D
D;kR#CQ   371a_tpmQzB_ht1Qh3 7N;DD
Ck#R Q  03#8F_Do_HON0sHED3NDz;
1Q R 3  MCkls_HO#308q;pp
M
C0$H0R_1A)cqvj_v]4RniH
#
RCRoMHCsORR5
RSSR)RWQ_a v m7RH:RMo0CC:sR=;RjRR
RSRRRRRRR)7 q_7vm :RRR0HMCsoCRR:=j
;R
RRRRRRRRRRRQahQ_:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQna_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QagRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQqa_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ a_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"RR

RRRRRRRRRhRQQ4a_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;R
RRRRRRRRRRRQahQ_R.j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R..:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R. :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"RR

RRRRRRRRRhRQQda_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"RR
RRRRRRRRR2RRR
;
RRRRRRRRRFRbsR05
RRRRRRRRRRRRRRRRq)7a:qRR0FkR8#0_oDFHPO_CFO0s45R68RRF0IMF2RjRR;
RRRRRRRRRRRRR)RRBRpiRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRR)RRB piRH:RM#RR0D8_FOoHRR:=';]'
RRRRRRRRRRRRRRRRR) R:RRRRHMR8#0_oDFH:OR=]R''R;
RRRRRRRRRRRRR)RRq)77RH:RM#RR0D8_FOoH_OPC05FsRRgR8MFI0jFR2
R;RRRRRRRRRRRRRRRRWiBpRRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRRWiBp RR:HRMR#_08DHFoO=R:R''];R
RRRRRRRRRRRRRR RWRRRR:MRHR0R#8F_DoRHO:'=R]
';RRRRRRRRRRRRRRRRW7q7)RR:HRMR#_08DHFoOC_POs0F5RRgRI8FMR0Fj;2R
RRRRRRRRRRRRRRRR1vqi:RRRRHMR8#0_oDFHPO_CFO0s45R68RRF0IMF2RjRR;
RRRRRRRRRRRRRWRR7qqaRH:RM#RR0D8_FOoH_OPC05FsRR46RI8FMR0FjR2
RRRRRRRRRRRRR;R2

RRRCR
M18RAq_)vvcj]n_4i
;
NEsOHO0C0CksR_1A)cqvj_v]4_niq])BRRFV1)A_qjvcv4]_nHiR#C
LoRHM
8CMR_1A)cqvj_v]4_niq])B;RRR-R--1)A_qjvcv4]_n
i

---------------------------------------
-S--AR1_v)qc]jv_i4nh-)
-------------------------------------D-
HNLssQ$R ;  
Ck#R Q  a317m_pt_QB4c4n3DND;#
kC RQ 1 3ap7_mBtQ_1zhQ th7D3NDk;
#QCR 3  #_08DHFoOs_NH30EN;DD
 z1R Q  k3MlHCsO0_#8p3qp
;
CHM001$RAq_)vvcj]n_4iRh)H
#
RCRoMHCsORR5
RSSR)RWQ_a v m7RH:RMo0CC:sR=;RjRR
RSRRRRRRR)7 q_7vm :RRR0HMCsoCRR:=j
;R
RRRRRRRRRRRQahQ_:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQna_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QagRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQqa_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ a_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"RR

RRRRRRRRRhRQQ4a_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;R
RRRRRRRRRRRQahQ_R.j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R..:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R. :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"RR

RRRRRRRRRhRQQda_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"RR
RRRRRRRRR2RRRR;
RRRRRRRRRsbF0
5RRRRRRRRRRRRRRRRR)a7qqRR:FRk0#_08DHFoOC_POs0F56R4RFR8IFM0RRj2;R
RRRRRRRRRRRRRRBR)pRih:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRBR)pRi :MRHR0R#8F_DoRHO:'=R]
';RRRRRRRRRRRRRRRR)R RRRR:HRMR#_08DHFoO=R:R''];R
RRRRRRRRRRRRRRqR)7R7):MRHR0R#8F_Do_HOP0COFRs5g8RRF0IMF2RjRR;
RRRRRRRRRRRRRWRRBRpiRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRRWRRB piRH:RM#RR0D8_FOoHRR:=';]'
RRRRRRRRRRRRRRRRRW R:RRRRHMR8#0_oDFH:OR=]R''R;
RRRRRRRRRRRRRWRRq)77RH:RM#RR0D8_FOoH_OPC05FsRRgR8MFI0jFR2
R;RRRRRRRRRRRRRRRRviq1RRR:HRMR#_08DHFoOC_POs0F56R4RFR8IFM0RRj2;R
RRRRRRRRRRRRRR7RWqRaq:MRHR0R#8F_Do_HOP0COFRs54R6R8MFI0jFR2R
RRRRRRRRRRRRRR
2;RRR
RM
C8AR1_v)qc]jv_i4nh
);
ONsECH0Os0kCAR1_v)qc]jv_i4nhq)_)RB]F1VRAq_)vvcj]n_4iRh)HL#
CMoHRM
C8AR1_v)qc]jv_i4nhq)_);B]R-RR-1-RAq_)vvcj]n_4i
h)
-
---------------------------------------
S-1-RAq_)vvcj]n_4i
hW-------------------------------------
--DsHLNRs$Q   ;#
kC RQ 1 3ap7_mBtQ_n44cD3NDk;
#QCR 3  1_a7pQmtBh_z1hQt N73D
D;kR#CQ   38#0_oDFHNO_sEH03DND;1
z  RQ M 3kslCH#O_0q83p
p;
0CMHR0$1)A_qjvcv4]_nWihR
H#
oRRCsMCH5ORRS
SRWRR) Qa_7vm RR:HCM0oRCs:j=R;RR
RRSRRRRRRq) 7m_v7R R:MRH0CCos=R:RRj;
R
RRRRRRRRRRQQhaR_j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QanRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ(a_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QaqRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQAa_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQwa_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;
R
RRRRRRRRRQRRh_Qa4:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjR";
R
RRRRRRRRRRQQhaj_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha4_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha._.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhad_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhac_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha6_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhan_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha(_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaU_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhag_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaq_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaA_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaB_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha7_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha _.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaw_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;
R
RRRRRRRRRQRRh_Qad:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
"RRRRRRRRRRRRR2
R;RRRRRRRRRFRbsR05
RRRRRRRRRRRRRRRRq)7a:qRR0FkR8#0_oDFHPO_CFO0s45R68RRF0IMF2RjRR;
RRRRRRRRRRRRR)RRBRpiRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRR)RRB piRH:RM#RR0D8_FOoHRR:=';]'
RRRRRRRRRRRRRRRRR) R:RRRRHMR8#0_oDFH:OR=]R''R;
RRRRRRRRRRRRR)RRq)77RH:RM#RR0D8_FOoH_OPC05FsRRgR8MFI0jFR2
R;RRRRRRRRRRRRRRRRWiBphRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRRWiBp RR:HRMR#_08DHFoO=R:R''];R
RRRRRRRRRRRRRR RWRRRR:MRHR0R#8F_DoRHO:'=R]
';RRRRRRRRRRRRRRRRW7q7)RR:HRMR#_08DHFoOC_POs0F5RRgRI8FMR0Fj;2R
RRRRRRRRRRRRRRRR1vqi:RRRRHMR8#0_oDFHPO_CFO0s45R68RRF0IMF2RjRR;
RRRRRRRRRRRRRWRR7qqaRH:RM#RR0D8_FOoH_OPC05FsRR46RI8FMR0FjR2
RRRRRRRRRRRRR;R2

RRRCR
M18RAq_)vvcj]n_4i;hW
s
NO0EHCkO0s1CRAq_)vvcj]n_4i_hWq])BRRFV1)A_qjvcv4]_nWihR
H#LHCoMCR
M18RAq_)vvcj]n_4i_hWq])B;RRR-R--1)A_qjvcv4]_nWih



-------------------------------------
--S---R_1A)cqvj_v]4hni)
hW-------------------------------------
--DsHLNRs$Q   ;#
kC RQ 1 3ap7_mBtQ_n44cD3NDk;
#QCR 3  1_a7pQmtBh_z1hQt N73D
D;kR#CQ   38#0_oDFHNO_sEH03DND;1
z  RQ M 3kslCH#O_0q83p
p;
0CMHR0$1)A_qjvcv4]_n)ihhHWR#R

RMoCCOsHR
5RSRSRRQW)av _mR7 :MRH0CCos=R:RRj;
SRRRRRRR)RR _q7v m7RRR:HCM0oRCs:j=R;
R
RRRRRRRRRQRRh_QajRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QacRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ6a_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QaURR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQga_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QaBRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ7a_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_ :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjR";
R
RRRRRRRRRRQQhaj_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha4_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha._4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhad_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhac_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha6_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhan_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha(_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaU_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhag_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaq_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaA_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaB_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha7_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha _4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaw_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;
R
RRRRRRRRRQRRh_Qa.:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa.:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa.:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa.:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa.:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa.:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa.:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa.:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa.:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa.:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa.:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa.:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa.:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa.:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa.: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa.:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjR";
R
RRRRRRRRRRQQhaj_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha4_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha._dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhad_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhac_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha6_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhan_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha(_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaU_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhag_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaq_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaA_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaB_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha7_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha _dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaw_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jjRR
RRRRRRRRRRRR2;R
RRRRRRRRRb0Fs5RR
RRRRRRRRRRRRR)RR7qqaRF:Rk#0R0D8_FOoH_OPC05FsRR46RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRp)Bi:hRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRp)Bi: RRRHMR8#0_oDFH:OR=]R''R;
RRRRRRRRRRRRR)RR RRRRH:RM#RR0D8_FOoHRR:=';]'
RRRRRRRRRRRRRRRR7)q7:)RRRHMR8#0_oDFHPO_CFO0sg5RRFR8IFM0RRj2;R
RRRRRRRRRRRRRRBRWpRih:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRBRWpRi :MRHR0R#8F_DoRHO:'=R]
';RRRRRRRRRRRRRRRRWR RRRR:HRMR#_08DHFoO=R:R''];R
RRRRRRRRRRRRRRqRW7R7):MRHR0R#8F_Do_HOP0COFRs5g8RRF0IMF2RjRR;
RRRRRRRRRRRRRvRRqR1iRH:RM#RR0D8_FOoH_OPC05FsRR46RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRqW7a:qRRRHMR8#0_oDFHPO_CFO0s45R68RRF0IMF2Rj
RRRRRRRRRRRRRRR2R;
RR
R
8CMR_1A)cqvj_v]4hni);hW
s
NO0EHCkO0s1CRAq_)vvcj]n_4ihh)W)_qBF]RVAR1_v)qc]jv_i4nhW)hR
H#LHCoMCR
M18RAq_)vvcj]n_4ihh)W)_qBR];R-R--AR1_v)qc]jv_i4nhW)h




