------------------------------------------------------------------------
@E
---a-RERH#VCHDR#ENRR0FL#CREbHbCC8RM$Osb80C!
!!-a-RERH#VCHDRF#EkRD8MCCPsCRLRH#Eb8bCRRHMs8CNNCLDRsVFl!!!

---a-RERH#P#CsHRFMF0VREvCRq_a]BumvpR Xb	NONRoCH-#
-bR1CVOHH0ORF$R1MHbDVN$RMH8R#FRM0#RkNCLDRsVFRl#Hk0DNH
FM-B-RFsb$H0oER25ORg4gc1,R$DMbH0OH$Q,RMRO3qRDDsEHo0s#RCs#CP
C8---
-ERaC>R=RCFbsFN0s#RHRCk#8FR0RC#bO$HVRLNRk0HDRRHMHDlbCMlC0HN0F
MR-V-RFNsRRb0$CsRFRMVkOF0HM-3
--
-RCaER8FsCFsRVkRVMHO0FRM#NRM88DCON0sNH#FMRRH#MRF0HM8C0NHODFR0RC0E
R--FosHHDMNRsPC#MHFRsVFRO#Ck0sH$CRsNM#F#-3
--
-RCf]Ns8C:/R/#b$MDHHO0O$/F.lbjJ4U./b4ObFlHsDC#E/P8PD/El8/N_0EObFlD3CGPyE84
Rf---
-FRwskRwsC0EsCR8#HOsbF0HMCR80DNH#b,RD#CNCFRDFN	R0FROlMlC0L#RCIDF:-
------------------------------------------------------------------------
--
-RbBF$osHE40RgRgnLQ$R 3  RDqDRosHER0#sCC#s8PC3-
-
R--a#EHRk#FsROCVCHDRRH#NCMR#M#C0DHNRsbN0VRFR Q  0R18jR4(.n3-g4gnQ,R R  1M0N88NsR-
-R7e]pNRv0lECNO0HNuDRNNO	o3C#RHaE#FR#kCsORDVHCNRl$FRM0CRLRbOFH,C8RD#F8F,Rs-R
-MRHO8DkCI8RHR0E#0FVICNsRN0E0#RHRD#F8HRI0kEF0sRIHC00MCRbs#lH#MHFRFVslER0C RQ - 
-0R1NNM8sR8#7NCbsC0lMR03a#EHRk#FsROCVCHDR$lNRRLCk8#CRR0FHDlbCMlC0ER0H##R08NMNRs8
R--NRM8lRN$L8CRHs#0H0LkCH8RMFROlDbHCV8RFRslHNMRMl$RNCMMsFR#RMDFo#RNRC0ER-
-RlOFbCHD8FRVs8lRFRC#MRF0NFDDIHR8s0CORO8CFHlbDHN0FFMRVER0CsRFHMoHN#DRFOksCHRVD
C3-a-RERH##sFkOVCRHRDClRN$LOCRFCbH8FRVsMRH8HHP8DkNRCk#R0LCIMCCRODHCCM#8#RkC3s#R-
-RHaE#FR#kCsORDVHC#RHRFbsPCH88MRFRRNMqQ1R1NRL#3H#RCaER Q  HR8#NODHRl#qRhY
R--W)q)qYhaRu X)1 1RRm)QpvuQR 7QphBzh7QthRqYqRW)h)qamYRw Rv)qB]hAaqQapQY-R
-hRq7QRwa1h 1mRw)1Rz mRw)RRquaq)QpBzqu)Rzm)u1R 3aRECks#CRRFV0REC#sFkO
CR-V-RHRDC#DENDMRH8MClHRV$NRM8E8FDR Q  NREsClD#V#RsRFlNRM$8NNloRC#FDsRHHNLD$H0R-
-RHNs#oHMR0FkRRFV0RECkR#C0sECC3FV

---a-RHC0D:RRRRRRR1M0N88NsR7e]pNRv0lECNO0HNuDRNNO	oRC#5 Q  0R18jR4(.n3-g4gn-,
-RRRRRRRRRRRRvRRq_a]Bumvp2 X

---p-RHNLssR$:RRRRa#EHRObN	CNoRN#EDLDRCFROlDbHCH8RMR0FNHRDLssN$-
-RRRRRRRRRRRRR$R#lDLFHDONDM$RN8lCR Q  -3
--
-RP7CCbDFC:s#R RQ 7 RqR1Bep]7R0vNENCl0NHODNRuOo	NCW#RFHs	MtoRsbFk

---u-RkFsb#RC:RRRRa#EHRObN	CNoRV8CH#MCR#NR08NMNRs8VRFs8HC#osMC#FR0RCk#R
HM-R-RRRRRRRRRRRRR8OC#sHHLMeoR]R7plCF8D0#RERN0lCN	RCk#RRFVOlFlFBMRmpvu -X
-RRRRRRRRRRRRORRF0M#N#M0R8NMRlOFlRFMBumvpR XlEN0C0lNHDONRMVkOF0HMN#RM-8
-RRRRRRRRRRRRFRRbNCs0#Fs3-
-
R--pHHl0HN0FRM:RCaERDPNkRC#oCCMsCN08$RLRC0ERMVkOF0HMH#RMER0Hb#RNNO	olCRN-$
-RRRRRRRRRRRRPRRNRs$VlsFRNbD0sVFlFR0RNbD0sVFlN,RM08REbCRsHCO#MHFRRFVskC#D
0#-R-RRRRRRRRRRRRRHF#RMRD$oskNNCM0C08RFCRLRC0ERMlHHllkRJsCkCHs8$RLR Q  0R18jR4(
n--R-RRRRRRRRRRRRR4dgg3-
-
R--hCF0#-:
-RRRRRRRRRRRRhRRFCR8OsDNNF0HMF#RsCR8VHHM0MHF#ER#NRDDLHCRMkOD8RC8HRM,F-s
-RRRRRRRRRRRRCRRGkOD8RC8VlsF,ER0Hb#RNNO	o
C3-R-RRRRRRRRRRRRRaREC"ObN	CNoRO8CDNNs0MHF"CR8VCHM#ER0C$R0b,C#RL#k0C$b#N,RM-8
-RRRRRRRRRRRR8RRCNODsHN0FRM#FvVRq_a]Bumvp3 X
R--RRRRRRRRRRRRRCaERN#0Ms8N8NRl0lECNO0HN8DRCMVHHF0HMMRN8FROMMPC0MHFNlDRCHNMM-o
-RRRRRRRRRRRRFRRVER0CNRl0lECNO0HNVDRk0MOH#FMRN0E0sRNCNRbsF0RVER0H##R08NMN
s8-R-RRRRRRRRRRRRRssCbCM#C0ER0CFRVsDlNRl#CNHM0OF#RVER0ClRHblDCCNM00MHFRRFV0
EC-R-RRRRRRRRRRRRRv]qa_vBmuXp RObN	CNoRO8CDNNs0MHF3aRREbCRkFsb#FCRVER0C-
-RRRRRRRRRRRRRqRvaB]_mpvu bXRNNO	oLCRFR8$H0#RFsRbF8PHCRRNo8kHCMDHCFRVs-
-RRRRRRRRRRRRRlRHblDCCNM00MHF#FR0RsPCHRV$0HECslRHblDCCNM00MHFRRFVv]qa_vBmuXp 3-
-RRRRRRRRRRRRRFRaF8DRCDPCFsbC#NRl$EROFCF#RR0FHDlbCMlC0ER0CNRbOo	NCFRL8H$RM-
-RRRRRRRRRRRRRER0CFRl#C0RVOVHH0CMRMlNMRCsNHPNDDNLCFR0RC0El-3
--
-R------------------------------------------------------------------------------
-CResF#HMRRRR4:R3-6
-NR70RCRRRRRR.:RckRKD4$Rg
gn---R----------------------------------------------------------------------------
#
kCmRW)vi3q_a])p q3DND;N
bOo	NCqRvaB]_mpvu HXR#R
RRFROMN#0MB0RF)b$H0oEhHF0ORC:1Qa)hRt
RRRRRR:="bBF$osHE40RgRgnQ   3DRqDHRso#E0R#sCCCsP8;3"
R
RR-R-
RRRRR--aC$bRV7CH0MHH#FM
RRRR
--RRRR0C$bRvBmuXp R
H#RRRRRRRRsFCOsR8
RRRRRRRRRRRRR)RR ):R ;qpRRRRRRRR-)-RCRNDb0Ns
RRRRRRRRRRRRRRRR:QvRq) pR;RRRRRR-R-RNQloNHMsb$RN
s0RRRRRRRRCRM8sFCOs
8;
RRRRL#k0C$bR1umQeaQ  _)qHpR# R)qspRNCMoRjj3RR0F)p q't]Q]
;
RRRR#0kL$RbCuh)QBqQupq_epRz H)#R RqpsoNMCvR-q_a]u0QRFqRvau]_Q
;
RRRR0C$bRvBmuXp _pumqH)R#R
RRRRRRCRsO8Fs
RRRRRRRRRRRRRRRRtvq:mRu1QQae) _ ;qpRRRR-v-RNHoM0Ck8
RRRRRRRRRRRRRRRRtq):)RuQQhBu_qpezqp R;R-q-RMCoDRRHMsHN8N;M#Rq-vau]_Q#RHRDHDCDoN
RRRRRRRR8CMROsCF;s8
R
RR-R-
RRRRR--B#FM00NMRV7CH0MHH#FM
RRRR
--RRRRO#FM00NMRqRvaB]_A q1_R4:BumvpR X:B=Rmpvu 5X'4,3jRjj32R;
RORRF0M#NRM0Ravq]A_Bq_1 KB:Rmpvu :XR=mRBv upXj'53Rj,423j;R
RRFROMN#0MR0Rv]qa_ BZ)Rm:BumvpR X:B=Rmpvu 5X'j,3jRjj32
;

RRRR
--RRRR-m-RPDCsFCN88JRCkHND0N$RMH8RMkCJN0DH$bRFC0sNFRs#VRFsBumvp_ Xuqmp)R
RR-R-RJ5CkHND0N$RMH8RMkCJN0DH$bRFC0sNFRs#VRFsBumvpR XNRsCb8sCCMVHC
82RRRR-
-
RRRRVOkM0MHFR="/"RR5pH:RMmRBv upXm_up;q)R:R)RRHMBumvp_ Xuqmp)RR2skC0sAMRm mpq
h;RRRRRRRR-u-RkFsb#
C:RRRRRRRR-R-RRRRRR)RRCs0kMa#R)Rz HpVRRRH#MRF0CNJkDFR0RN)RMs8RCs0kMw#Rq p1
RRRRRRRRR--RRRRRRRRFC0Es#IHCR
RRRRRR-R-RC1bODHNRDPNk:C#
RRRRRRRRR--RRRRRRRRBumvp_ Xuqmp)j'53Rj,X/2R=mRBv upXm_up'q)5jj3,2RYR0sCk#sM
RRRRRRRRR--RRRRRRRRw1qp CRso8NsD#C#RRFV0RECPkNDCVRFRNXRMY8R3R
RRRRRR-R-Rl7FN:HM
RRRRRRRRR--RRRRRRRRpMRHRvBmuXp _pumqN)RMp8R3tq)RR/=-avq]Q_u
RRRRRRRRR--RRRRRRRR)MRHRvBmuXp _pumqN)RM)8R3tq)RR/=-avq]Q_u
RRRRRRRRR-- FsssFROM08HH#FM:R
RRRRRR-R-RRRRRRRRRs sFHsRV3RpqR)t=vR-q_a]uRQ
RRRRR-RR-RRRRRRRRsR sRFsH)VR3tq)R-=Rv]qa_
uQRRRRRRRR-)-RNCMo:R
RRRRRR-R-RRRRRRRRR="/",5p)H2R#HRC0sECRza) sRFRpwq1R 
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRRRRhCFM
R
RRkRVMHO0F"MR=5"RRRp:HBMRmpvu uX_m)pq;)RR:MRHRvBmuXp _pumq2)RR0sCkRsMApmm ;qh
RRRRRRRRR--ubksF:#C
RRRRRRRRR--RRRRRRRR)kC0sRM#a )zRRHVp#RHRkCJN0DRFRR)NRM8skC0sRM#w1qp 0RFEICsH
#CRRRRRRRR-1-RbHCONPDRNCDk#R:
RRRRR-RR-RRRRRRRRmRBv upXm_up'q)5jj3,2RXRB=Rmpvu uX_m)pq'35jjY,R2CRs0Mks#)RazR 
RRRRR-RR-RRRRRRRRCRso8NsD#C#RRFV0RECPkNDCVRFRNXRMY8R3R
RRRRRR-R-Rl7FN:HM
RRRRRRRRR--RRRRRRRRpMRHRvBmuXp _pumqN)RMp8R3tq)RR/=-avq]Q_u
RRRRRRRRR--RRRRRRRR)MRHRvBmuXp _pumqN)RM)8R3tq)RR/=-avq]Q_u
RRRRRRRRR-- FsssFROM08HH#FM:R
RRRRRR-R-RRRRRRRRRs sFHsRV3RpqR)t=vR-q_a]uRQ
RRRRR-RR-RRRRRRRRsR sRFsH)VR3tq)R-=Rv]qa_
uQRRRRRRRR-)-RNCMo:R
RRRRRR-R-RRRRRRRRR""=5)p,2#RHR0CHERCsa )zRRFsw1qp R
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRRhRRF
MC
RRRR
--RRRR-w-Rk0MOHRFM7DCON0sNH#FM
RRRR
--RRRRVOkM0MHFRat _Qu)huBQqep_q pz5RX:H)MR Rqp2CRs0MksRQu)huBQqep_q pz;R
RRRRRR-R-RsukbCF#:R
RRRRRR-R-RRRRRRRRR0)Ck#sMRHbsMbOHNPDRNCDkRRFVNDMoC;RXRHXRMNRs8MHN#R
RRRRRR-R-RC1bODHNRDPNk:C#
RRRRRRRRR--RRRRRRRRhCFM
RRRRRRRRR--7NFlH
M:RRRRRRRR-R-RRRRRRXRRRRHM)p q
RRRRRRRRR-- FsssFROM08HH#FM:R
RRRRRR-R-RRRRRRRRRMhFCR
RRRRRR-R-RM)No
C:RRRRRRRR-R-RRRRRR-RRv]qa_RuQ< Rta)_uQQhBu_qpezqp 25XRR<=v]qa_
uQRRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRRMhFCR

RVRRk0MOHRFMBpvuX:5XRRHM)p q;YRR:MRHRq) pR:=jR3j2CRs0MksRvBmuXp ;R
RRRRRR-R-RsukbCF#:R
RRRRRR-R-RRRRRRRRR0)Ck#sMRvBmuXp RlMkLRCsXRR+HRY
RRRRR-RR-bR1CNOHDNRPD#kC:R
RRRRRR-R-RRRRRRRRRMhFCR
RRRRRR-R-Rl7FN:HM
RRRRRRRRR--RRRRRRRRXMRHRq) pR
RRRRRR-R-RRRRRRRRRHYRM R)qRp
RRRRR-RR-sR sRFsO8FMHF0HM
#:RRRRRRRR-R-RRRRRRhRRF
MCRRRRRRRR-)-RNCMo:R
RRRRRR-R-RRRRRRRRRuBvpXX5,RY2Hl#RNC0ElHN0ODND$MRkLMFk8
C8RRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRRMhFCR

RVRRk0MOHRFMuqmp)m_a_vBmuXp 5RZ:HBMRmpvu uX_m)pqRs2RCs0kMmRBv upXR;
RRRRR-RR-kRus#bFCR:
RRRRR-RR-RRRRRRRRCR)0Mks#mRBv upXNRPDRkCFZVR
RRRRRRRRR--1ObCHRNDPkNDC
#:RRRRRRRR-R-RRRRRRhRRF
MCRRRRRRRR-7-RFHlNMR:
RRRRR-RR-RRRRRRRRRRZHBMRmpvu uX_m)pqR8NMRqZ3)/tR=vR-q_a]uRQ
RRRRR-RR-sR sRFsO8FMHF0HM
#:RRRRRRRR-R-RRRRRR RRsssFRRHVZ)3qtRR=-avq]Q_u
RRRRRRRRR--)oNMCR:
RRRRR-RR-RRRRRRRRmRup_q)aBm_mpvu ZX52#RHR0lNENCl0NHODRD$kFMLkCM88R
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRRhRRF
MC
RRRRMVkOF0HMmRBv upXm_a_pumqZ)5:MRHRvBmuXp Rs2RCs0kMmRBv upXm_up;q)
RRRRRRRRR--ubksF:#C
RRRRRRRRR--RRRRRRRR)kC0sRM#bMsHONHbDNRPDRkCBumvp_ Xuqmp)VRFRRZ
RRRRR-RR-bR1CNOHDNRPD#kC:R
RRRRRR-R-RRRRRRRRRvBmuXp __amuqmp)q5vaB]_Zm )2RR=Bumvp_ Xuqmp)j'53Rj,j23j
RRRRRRRRR--RRRRRRRRBumvp_ Xaum_m)pq5RZ2=mRBv upXm_up'q)51qA5QZ3v
2,RRRRRRRR-R-RRRRRRRRRRRRRRRRRRRRRRRRRRRRR1hQt5QZ3vv2*q_a]umQ_e_ ).H2RV3RZ)= RRjj3
RRRRRRRRR--7NFlH
M:RRRRRRRR-R-RRRRRRZRRRRHMBumvp
 XRRRRRRRR- -RsssFRMOF8HH0F:M#
RRRRRRRRR--RRRRRRRRhCFM
RRRRRRRRR--)oNMCR:
RRRRR-RR-RRRRRRRRCRs#0kD3tvqRR>=j
3jRRRRRRRR-R-RRRRRR-RRv]qa_RuQ<CRs#0kD3tq)RR<=v]qa_
uQRRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRRMhFCR

RVRRk0MOHRFM"1qA":5ZRRHMBumvp_ Xuqmp)RR2skC0suMRma1QQ_e )p q;R
RRRRRR-R-RsukbCF#:R
RRRRRR-R-RRRRRRRRR0)Ck#sMR#NLF0DkCNRPDRkC5olNMkH08RC2FZVR
RRRRRRRRR--1ObCHRNDPkNDC
#:RRRRRRRR-R-RRRRRRhRRF
MCRRRRRRRR-7-RFHlNMR:
RRRRR-RR-RRRRRRRRRRZHBMRmpvu uX_m)pqR8NMRqZ3)/tR=vR-q_a]uRQ
RRRRR-RR-sR sRFsO8FMHF0HM
#:RRRRRRRR-R-RRRRRR RRsssFRRHVZ)3qtRR=-avq]Q_u
RRRRRRRRR--)oNMCR:
RRRRR-RR-RRRRRRRRARq125ZRR>=j
3jRRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRR1qA5RZ2=3RZv
qt
RRRRMVkOF0HMqR"A51"ZH:RMmRBv upXRR2skC0suMRma1QQ_e )p q;R
RRRRRR-R-RsukbCF#:R
RRRRRR-R-RRRRRRRRR0)Ck#sMR#NLF0DkCNRPDRkC5olNMkH08RC2FZVR
RRRRRRRRR--1ObCHRNDPkNDC
#:RRRRRRRR-R-RRRRRRhRRF
MCRRRRRRRR-7-RFHlNMR:
RRRRR-RR-RRRRRRRRRRZHBMRmpvu RX
RRRRR-RR-sR sRFsO8FMHF0HM
#:RRRRRRRR-R-RRRRRRhRRF
MCRRRRRRRR-)-RNCMo:R
RRRRRR-R-RRRRRRRRR1qA5RZ2Hl#RNC0ElHN0ODND$MRkLMFk8
C8RRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRR1qA5RZ2=TR1)Za53*) Z 3)RZ+R3*QvZv3Q2R

RVRRk0MOHRFMq5)tZH:RMmRBv upXm_upRq)2CRs0MksRQu)huBQqep_q pz;R
RRRRRR-R-RsukbCF#:R
RRRRRR-R-RRRRRRRRR0)Ck#sMRoNskMlC0NR5MCoD2MRHR8sNH#NMRRFV0RECbMsHONHbDR
RRRRRR-R-RRRRRRRRRDPNkFCRV
RZRRRRRRRR-1-RbHCONPDRNCDk#R:
RRRRR-RR-RRRRRRRRFRhMRC
RRRRR-RR-FR7lMNH:R
RRRRRR-R-RRRRRRRRRHZRMmRBv upXm_upRq)NRM8Z)3qt=R/Rq-vau]_QR
RRRRRR-R-Rs sFOsRFHM80MHF#R:
RRRRR-RR-RRRRRRRRsR sRFsHZVR3tq)R-=Rv]qa_
uQRRRRRRRR-)-RNCMo:R
RRRRRR-R-RRRRRRRRRq-vau]_QRR<q5)tZ<2R=qRvau]_QR
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRRqRR)Zt52RR=Z)3qt


RRRRVOkM0MHFRtq)5RZ:HBMRmpvu 2XRR0sCkRsMuh)QBqQupq_ep;z 
RRRRRRRRR--ubksF:#C
RRRRRRRRR--RRRRRRRR)kC0sRM#Nksol0CMRM5No2DCRRHMsHN8NRM#F0VREbCRsOHMHDbN
RRRRRRRRR--RRRRRRRRPkNDCVRFRRZ
RRRRR-RR-bR1CNOHDNRPD#kC:R
RRRRRR-R-RRRRRRRRRtq)5RZ2=3RjjVRHR)Z3 =R>Rjj3R8NMRQZ3vRR=j
3jRRRRRRRR-R-RRRRRRqRR)Zt52RR=1hQt5QZ3vv2*q_a]umQ_e_ ).VRHR)Z3 RR=j
3jRRRRRRRR-R-RRRRRRqRR)Zt52RR=v]qa_RuQHZVR3R) <3RjjRRRRRRRR8NMRQZ3vRR=j
3jRRRRRRRR-7-RFHlNMR:
RRRRR-RR-RRRRRRRRRRZHBMRmpvu RX
RRRRR-RR-sR sRFsO8FMHF0HM
#:RRRRRRRR-R-RRRRRRhRRF
MCRRRRRRRR-)-RNCMo:R
RRRRRR-R-RRRRRRRRRq-vau]_QRR<q5)tZ<2R=qRvau]_QR
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRRqRR)Zt52RR=qa)BqZh53,QvR)Z3 
2
RRRRVOkM0MHFR""-R:5ZRRHMBumvp_ Xuqmp)RR2skC0sBMRmpvu uX_m)pq;R
RRRRRR-R-RsukbCF#:R
RRRRRR-R-RRRRRRRRR0)Ck#sMRHbsMbOHNPDRNCDkRRFVksMN$HRlMRk#FZVR
RRRRRRRRR--1ObCHRNDPkNDC
#:RRRRRRRR-R-RRRRRR"RR-Z"52RR=Bumvp_ Xuqmp)Z'53tvq,qRvau]_QH2RV3RZqR)t=3RjjR
RRRRRR-R-Rl7FN:HM
RRRRRRRRR--RRRRRRRRZMRHRvBmuXp _pumqN)RMZ8R3tq)RR/=-avq]Q_u
RRRRRRRRR-- FsssFROM08HH#FM:R
RRRRRR-R-RRRRRRRRRs sFHsRV3RZqR)t=vR-q_a]uRQ
RRRRR-RR-NR)M:oC
RRRRRRRRR--RRRRRRRRskC#Dv03q>tR=3RjjR
RRRRRR-R-RRRRRRRRRq-vau]_QRR<skC#Dq03)<tR=qRvau]_QR
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRR)RRCs0kMB#Rmpvu uX_m)pq'35Zv,qtRqZ3)-tRRt1Qh35Zq2)t*avq]Q_u2VRH
RRRRRRRRR--RRRRRRRRRRRRRZRR3tq)RR/=j
3j
RRRRMVkOF0HM-R""ZR5:MRHRvBmuXp Rs2RCs0kMmRBv upXR;
RRRRR-RR-kRus#bFCR:
RRRRR-RR-RRRRRRRRCR)0Mks#MRkNRs$lkHM#VRFRRZ
RRRRR-RR-bR1CNOHDNRPD#kC:R
RRRRRR-R-RRRRRRRRRMhFCR
RRRRRR-R-Rl7FN:HM
RRRRRRRRR--RRRRRRRRZMRHRvBmuXp 
RRRRRRRRR-- FsssFROM08HH#FM:R
RRRRRR-R-RRRRRRRRRMhFCR
RRRRRR-R-RM)No
C:RRRRRRRR-R-RRRRRR"RR-Z"52#RHR0lNENCl0NHODRD$kFMLkCM88R
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRR)RRCs0kM-#RG[R-$FRVs=RZR+GRR
[$
RRRRMVkOF0HMmRBh5KRZH:RMmRBv upXm_up2q)R0sCkRsMBumvp_ Xuqmp)R;
RRRRR-RR-kRus#bFCR:
RRRRR-RR-RRRRRRRRCR)0Mks#sRbHHMObRNDPkNDCVRFRlOFbGDCRMOF[Nko0FCRV
RZRRRRRRRR-1-RbHCONPDRNCDk#R:
RRRRR-RR-RRRRRRRRmRBhZK52RR=Bumvp_ Xuqmp)Z'53tvq,qRvau]_QH2RV3RZqR)t=qRvau]_QR
RRRRRR-R-Rl7FN:HM
RRRRRRRRR--RRRRRRRRZMRHRvBmuXp _pumqN)RMZ8R3tq)RR/=-avq]Q_u
RRRRRRRRR-- FsssFROM08HH#FM:R
RRRRRR-R-RRRRRRRRRs sFHsRV3RZqR)t=vR-q_a]uRQ
RRRRR-RR-NR)M:oC
RRRRRRRRR--RRRRRRRRskC#Dv03q>tR=3RjjR
RRRRRR-R-RRRRRRRRRq-vau]_QRR<skC#Dq03)<tR=qRvau]_QR
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRR)RRCs0kMB#Rmpvu uX_m)pq'35Zv,qtR3-Zq2)tRRHVZ)3qt=R/Ravq]Q_u
R
RRkRVMHO0FBMRmRhK5RZ:HBMRmpvu RX2skC0sBMRmpvu 
X;RRRRRRRR-u-RkFsb#
C:RRRRRRRR-R-RRRRRR)RRCs0kMO#RFDlbCOGRFkM[oCN0RRFVZR
RRRRRR-R-RC1bODHNRDPNk:C#
RRRRRRRRR--RRRRRRRRhCFM
RRRRRRRRR--7NFlH
M:RRRRRRRR-R-RRRRRRZRRRRHMBumvp
 XRRRRRRRR- -RsssFRMOF8HH0F:M#
RRRRRRRRR--RRRRRRRRhCFM
RRRRRRRRR--)oNMCR:
RRRRR-RR-RRRRRRRRmRBhZK52#RHR0lNENCl0NHODRD$kFMLkCM88R
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRR)RRCs0kMG#RR$-[RsVFRRZ=GRR+[
$
RRRRVOkM0MHFR)1Ta:5ZRRHMBumvp_ Xuqmp)RR2skC0sBMRmpvu uX_m)pq;R
RRRRRR-R-RsukbCF#:R
RRRRRR-R-RRRRRRRRR0)Ck#sMRk#JNRsCs0FFRRFVZHRI0bERF0#HHRPCsDCNRsbN0R
RRRRRR-R-RRRRRRRRR,FsRRHV0RECsDCNRsbN0#RHRsxCF0,REFCRMICRHR0EMMFMC0oNH
PCRRRRRRRR-R-RRRRRRHRRlHNoM$NsRsbN0R
RRRRRR-R-RC1bODHNRDPNk:C#
RRRRRRRRR--RRRRRRRR1aT)5RZ2=mRBv upXm_up'q)5jj3,3RjjH2RV3RZvRqt=3RjjR
RRRRRR-R-Rl7FN:HM
RRRRRRRRR--RRRRRRRRZMRHRvBmuXp _pumqN)RMZ8R3tq)RR/=-avq]Q_u
RRRRRRRRR-- FsssFROM08HH#FM:R
RRRRRR-R-RRRRRRRRRs sFHsRV3RZqR)t=vR-q_a]uRQ
RRRRR-RR-NR)M:oC
RRRRRRRRR--RRRRRRRRskC#Dv03q>tR=3RjjR
RRRRRR-R-RRRRRRRRRq-vau]_QRR<skC#Dq03)<tR=qRvau]_QR
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRRhRRF
MC
RRRRMVkOF0HMTR1)Za5:MRHRvBmuXp Rs2RCs0kMmRBv upXR;
RRRRR-RR-kRus#bFCR:
RRRRR-RR-RRRRRRRRCR)0Mks#JR#kCNsRFsF0VRFRIZRHR0EbHF#0CHPRNsCDNRbsR0
RRRRR-RR-RRRRRRRRsRF,VRHRC0ERNsCDNRbsH0R#CRxsRF,0RECFRMCIEH0RMMFMNCo0CHP
RRRRRRRRR--RRRRRRRRHolNHsMN$NRbsR0
RRRRR-RR-bR1CNOHDNRPD#kC:R
RRRRRR-R-RRRRRRRRR)1Taq5vaB]_Zm )2RR=v]qa_ BZ)Rm
RRRRR-RR-FR7lMNH:R
RRRRRR-R-RRRRRRRRRHZRMmRBv upXR
RRRRRR-R-Rs sFOsRFHM80MHF#R:
RRRRR-RR-RRRRRRRRFRhMRC
RRRRR-RR-NR)M:oC
RRRRRRRRR--RRRRRRRR1aT)5RZ2Hl#RNC0ElHN0ODND$MRkLMFk8
C8RRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRRMhFCR

RVRRk0MOHRFM 5XuZH:RMmRBv upXm_upRq)2CRs0MksRvBmuXp _pumq
);RRRRRRRR-u-RkFsb#
C:RRRRRRRR-R-RRRRRR)RRCs0kMb#RsOHMHDbNRDPNkFCRVGRCbCFMMN0HDVRFRRZ
RRRRR-RR-bR1CNOHDNRPD#kC:R
RRRRRR-R-RRRRRRRRRu X5RZ2=mRBv upXm_up'q)5j43,3RjjH2RV3RZvRqt=jj3R8NM
RRRRRRRRR--RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRZRR3tq)Rj=R3Rj
RRRRR-RR-RRRRRRRRXR u25ZRB=Rmpvu uX_m)pq'354jv,Rq_a]uRQ2HZVR3tvqRv=Rq_a]uNQRMR8
RRRRR-RR-RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR1qA5qZ3)Rt2=qRvau]_Qe_m .)_
RRRRRRRRR--RRRRRRRR 5XuZ=2RRvBmuXp _pumq5)'4,3jRavq]Q_u_ me)2_.R
HVRRRRRRRR-R-RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR3RZvRqt=qRvau]_Qe_m .)_R8NM
RRRRRRRRR--RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRZRR3tq)Rv=Rq_a]umQ_e_ ).R
RRRRRR-R-RRRRRRRRRu X5RZ2=mRBv upXm_up'q)5j43,vR-q_a]umQ_e_ ).H2RVR
RRRRRR-R-RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRZq3vtRR=v]qa__uQm)e _N.RMR8
RRRRR-RR-RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRqZ3)=tRRq-vau]_Qe_m .)_
RRRRRRRRR--7NFlH
M:RRRRRRRR-R-RRRRRRZRRRRHMBumvp_ Xuqmp)MRN83RZqR)t/-=Rv]qa_
uQRRRRRRRR- -RsssFRMOF8HH0F:M#
RRRRRRRRR--RRRRRRRR FsssVRHRqZ3)=tRRq-vau]_QR
RRRRRR-R-RM)No
C:RRRRRRRR-R-RRRRRRsRRCD#k0q3vt=R>Rjj3
RRRRRRRRR--RRRRRRRR-avq]Q_uRs<RCD#k0)3qt=R<Ravq]Q_u
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRRFRhM
C
RRRRVOkM0MHFRu X5RZ:HBMRmpvu 2XRR0sCkRsMBumvp; X
RRRRRRRRR--ubksF:#C
RRRRRRRRR--RRRRRRRR)kC0sRM#CFGbM0CMHRNDFZVR
RRRRRRRRR--1ObCHRNDPkNDC
#:RRRRRRRR-R-RRRRRR RRXvu5q_a]B)Z m=2RRavq]A_Bq_1 4R
RRRRRR-R-RRRRRRRRRu X5RZ2=vR-q_a]B1Aq R_4HZVR3R) =3RjjMRN8ARq135ZQRv2=qRvau]_QR
RRRRRR-R-RRRRRRRRRu X5RZ2=QR1tZh532Qv*avq]A_Bq_1 KVRHR)Z3 RR=jR3jN
M8RRRRRRRR-R-RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRq5A1Zv3Q2RR=Ravq]Q_u_ me)
_.RRRRRRRR-7-RFHlNMR:
RRRRR-RR-RRRRRRRRRRZHBMRmpvu RX
RRRRR-RR-sR sRFsO8FMHF0HM
#:RRRRRRRR-R-RRRRRRhRRF
MCRRRRRRRR-)-RNCMo:R
RRRRRR-R-RRRRRRRRRu X5RZ2Hl#RNC0ElHN0ODND$MRkLMFk8
C8RRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRRMhFC



RRRRMVkOF0HMmRptZ.5:MRHRvBmuXp Rs2RCs0kMmRBv upXR;
RRRRR-RR-kRus#bFCR:
RRRRR-RR-RRRRRRRRCR)0Mks#FRDoHNs0RElLCN#RF.RV
RZRRRRRRRR-1-RbHCONPDRNCDk#R:
RRRRR-RR-RRRRRRRRmRptv.5q_a]B1Aq 2_4Rv=Rq_a]B)Z mR
RRRRRR-R-RRRRRRRRRtpm.25ZRv=Rq_a]B1Aq R_4HZVRRB=Rmpvu 5X'.,3jRjj32R
RRRRRR-R-Rl7FN:HM
RRRRRRRRR--RRRRRRRRZMRHRvBmuXp R8NMR1qA5RZ2/j=R3Rj
RRRRR-RR-sR sRFsO8FMHF0HM
#:RRRRRRRR-R-RRRRRR RRsssFRRHVq5A1Z=2RRjj3
RRRRRRRRR--)oNMCR:
RRRRR-RR-RRRRRRRRmRptZ.52#RHR0lNENCl0NHODRD$kFMLkCM88R
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRRhRRF
MC
RRRRMVkOF0HMmRpt:5ZRRHMBumvpR X2CRs0MksRvBmuXp ;R
RRRRRR-R-RsukbCF#:R
RRRRRR-R-RRRRRRRRR0)Ck#sMR0MNkDsNRoDFN0sHEFlRV
RZRRRRRRRR-1-RbHCONPDRNCDk#R:
RRRRR-RR-RRRRRRRRmRptq5vaB]_A q1_R42=qRvaB]_Zm )
RRRRRRRRR--RRRRRRRRp5mt-avq]A_Bq_1 4=2RRvBmuXp '35jjv,Rq_a]u
Q2RRRRRRRR-R-RRRRRRpRRmvt5q_a]B1Aq 2_KRB=Rmpvu 5X'j,3jRavq]Q_u_ me)2_.
RRRRRRRRR--RRRRRRRRp5mt-avq]A_Bq_1 K=2RRvBmuXp '35jj-,Rv]qa__uQm)e _
.2RRRRRRRR-R-RRRRRRpRRmZt52RR=v]qa_qBA14 _RRHVZRR=Bumvp' X5avq],_ Rjj32R
RRRRRR-R-Rl7FN:HM
RRRRRRRRR--RRRRRRRRZMRHRvBmuXp R8NMR1qA5RZ2/j=R3Rj
RRRRR-RR-sR sRFsO8FMHF0HM
#:RRRRRRRR-R-RRRRRR RRsssFRRHVq5A1Z=2RRjj3
RRRRRRRRR--)oNMCR:
RRRRR-RR-RRRRRRRRmRpt25ZRRH#lEN0C0lNHDONDk$RMkLFM88C
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRRFRhM
C
RRRRVOkM0MHFRtpm4Zj5:MRHRvBmuXp Rs2RCs0kMmRBv upXR;
RRRRR-RR-kRus#bFCR:
RRRRR-RR-RRRRRRRRCR)0Mks#FRDoHNs0RElLCN#RR4jFZVR
RRRRRRRRR--1ObCHRNDPkNDC
#:RRRRRRRR-R-RRRRRRpRRmjt45avq]A_Bq_1 4=2RRavq]Z_B 
)mRRRRRRRR-R-RRRRRRpRRmjt45RZ2=qRvaB]_A q1_H4RVRRZ=mRBv upX4'5j,3jRjj32R
RRRRRR-R-Rl7FN:HM
RRRRRRRRR--RRRRRRRRZMRHRvBmuXp R8NMR1qA5RZ2/j=R3Rj
RRRRR-RR-sR sRFsO8FMHF0HM
#:RRRRRRRR-R-RRRRRR RRsssFRRHVq5A1Z=2RRjj3
RRRRRRRRR--)oNMCR:
RRRRR-RR-RRRRRRRRmRpt54jZH2R#NRl0lECNO0HN$DDRLkMF8kMCR8
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRRRRhCFM
R
RRkRVMHO0FpMRm5t.ZH:RMmRBv upXm_upRq)2CRs0MksRvBmuXp _pumq
);RRRRRRRR-u-RkFsb#
C:RRRRRRRR-R-RRRRRR)RRCs0kMb#RsOHMHDbNRDPNkFCRVFRDoHNs0RElLCN#RF.RV
RZRRRRRRRR-1-RbHCONPDRNCDk#R:
RRRRR-RR-RRRRRRRRmRptZ.52RR=Bumvp_ Xuqmp)j'53Rj,j23jRRHVZq3vtRR=4R3jN
M8RRRRRRRR-R-RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRZ)3qtRR=j
3jRRRRRRRR-R-RRRRRRpRRm5t.Z=2RRvBmuXp _pumq5)'4,3jRjj32VRHRvZ3q=tRRj.3R8NM
RRRRRRRRR--RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRZ)3qtRR=j
3jRRRRRRRR-7-RFHlNMR:
RRRRR-RR-RRRRRRRRRRZHBMRmpvu uX_m)pqR8NMRqZ3)/tR=vR-q_a]uRQ
RRRRR-RR-RRRRRRRR3RZvRqt/j=R3Rj
RRRRR-RR-sR sRFsO8FMHF0HM
#:RRRRRRRR-R-RRRRRR RRsssFRRHVZ)3qtRR=-avq]Q_u
RRRRRRRRR--RRRRRRRR FsssVRHRvZ3q=tRRjj3
RRRRRRRRR--)oNMCR:
RRRRR-RR-RRRRRRRRCRs#0kD3tvqRR>=j
3jRRRRRRRR-R-RRRRRR-RRv]qa_RuQ<CRs#0kD3tq)RR<=v]qa_
uQRRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRhCFM
R
RRkRVMHO0FpMRmZt5:MRHRvBmuXp _pumq2)RR0sCkRsMBumvp_ Xuqmp)R;
RRRRR-RR-kRus#bFCR:
RRRRR-RR-RRRRRRRRCR)0Mks#sRbHHMObRNDPkNDCVRFR0MNkDsNRoDFN0sHEFlRV
RZRRRRRRRR-1-RbHCONPDRNCDk#R:
RRRRR-RR-RRRRRRRRmRpt25ZRB=Rmpvu uX_m)pq'35jjj,R3Rj2HZVR3tvqR4=R3NjRMR8
RRRRR-RR-RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR3RZqR)t=3RjjR
RRRRRR-R-RRRRRRRRRtpm5RZ2=mRBv upXm_up'q)5avq]Q_u,qRvau]_Qe_m .)_2VRH
RRRRRRRRR--RRRRRRRRRRRRRRRRRRRRRRRRRRRRRvZ3q=tRRj43R8NMRqZ3)=tRRavq]Q_u
RRRRRRRRR--RRRRRRRRp5mtZ=2RRvBmuXp _pumq5)'v]qa__uQm)e _R.,v]qa__uQm)e _R.2HRV
RRRRR-RR-RRRRRRRRRRRRRRRRRRRRRRRRRRRRZRR3tvqR4=R3NjRMR8RZ)3qtRR=v]qa__uQm)e _R.
RRRRR-RR-RRRRRRRRmRpt25ZRB=Rmpvu uX_m)pq'q5vau]_Qe_m .)_,vR-q_a]umQ_e_ ).H2RVR
RRRRRR-R-RRRRRRRRRRRRRRRRRRRRRRRRRRRRR3RZvRqt=3R4jMRN8ZRR3tq)R-=Rv]qa__uQm)e _R.
RRRRR-RR-RRRRRRRRmRpt25ZRB=Rmpvu uX_m)pq'354jj,R3Rj2HZVR3tvqRv=Rq_a] MRN8R
RRRRRR-R-RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRqZ3)=tRRjj3
RRRRRRRRR--7NFlH
M:RRRRRRRR-R-RRRRRRZRRRRHMBumvp_ Xuqmp)MRN83RZqR)t/-=Rv]qa_
uQRRRRRRRR-R-RRRRRRZRR3tvqRR/=j
3jRRRRRRRR- -RsssFRMOF8HH0F:M#
RRRRRRRRR--RRRRRRRR FsssVRHRqZ3)=tRRq-vau]_QR
RRRRRR-R-RRRRRRRRRs sFHsRV3RZvRqt=3RjjR
RRRRRR-R-RM)No
C:RRRRRRRR-R-RRRRRRsRRCD#k0q3vt=R>Rjj3
RRRRRRRRR--RRRRRRRR-avq]Q_uRs<RCD#k0)3qt=R<Ravq]Q_u
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRRFRhM
C
RRRRVOkM0MHFRtpm4Zj5:MRHRvBmuXp _pumq2)RR0sCkRsMBumvp_ Xuqmp)R;
RRRRR-RR-kRus#bFCR:
RRRRR-RR-RRRRRRRRCR)0Mks#sRbHHMObRNDPkNDCVRFRoDFN0sHELlRNR#C4FjRV
RZRRRRRRRR-1-RbHCONPDRNCDk#R:
RRRRR-RR-RRRRRRRRmRpt54jZ=2RRvBmuXp _pumq5)'j,3jRjj32VRHRvZ3q=tRRj43R8NM
RRRRRRRRR--RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR3RZqR)t=3RjjR
RRRRRR-R-RRRRRRRRRtpm4Zj52RR=Bumvp_ Xuqmp)4'53Rj,j23jRRHVZq3vtRR=4jj3R8NM
RRRRRRRRR--RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR3RZqR)t=3RjjR
RRRRRR-R-Rl7FN:HM
RRRRRRRRR--RRRRRRRRZMRHRvBmuXp _pumqN)RMZ8R3tq)RR/=-avq]Q_u
RRRRRRRRR--RRRRRRRRZq3vt=R/Rjj3
RRRRRRRRR-- FsssFROM08HH#FM:R
RRRRRR-R-RRRRRRRRRs sFHsRV3RZqR)t=vR-q_a]uRQ
RRRRR-RR-RRRRRRRRsR sRFsHZVR3tvqRj=R3Rj
RRRRR-RR-NR)M:oC
RRRRRRRRR--RRRRRRRRskC#Dv03q>tR=3RjjR
RRRRRR-R-RRRRRRRRRq-vau]_QRR<skC#Dq03)<tR=qRvau]_QR
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRRhRRF
MC
RRRRMVkOF0HMmRpt:5ZRRHMBumvp; XR1Aq H:RM R)qRp2skC0sBMRmpvu 
X;RRRRRRRR-u-RkFsb#
C:RRRRRRRR-R-RRRRRR)RRCs0kMD#RFsoNHl0ER#LNCqRA1F RV
RZRRRRRRRR-1-RbHCONPDRNCDk#R:
RRRRR-RR-RRRRRRRRmRptq5vaB]_A q1_R4,A q12RR=v]qa_ BZ)Rm
RRRRR-RR-RRRRRRRRmRpt,5ZA q12RR=v]qa_qBA14 _RRHVZRR=Bumvp' X51Aq j,R3
j2RRRRRRRR-7-RFHlNMR:
RRRRR-RR-RRRRRRRRRRZHBMRmpvu NXRMq8RAZ152=R/Rjj3
RRRRRRRRR--RRRRRRRRA q1Rj>R3Rj
RRRRR-RR-RRRRRRRRqRA1/ R=3R4jR
RRRRRR-R-Rs sFOsRFHM80MHF#R:
RRRRR-RR-RRRRRRRRsR sRFsHqVRAZ152RR=j
3jRRRRRRRR-R-RRRRRR RRsssFRRHVA q1RR<=j
3jRRRRRRRR-R-RRRRRR RRsssFRRHVA q1R4=R3Rj
RRRRR-RR-NR)M:oC
RRRRRRRRR--RRRRRRRRp5mtZq,A1R 2Hl#RNC0ElHN0ODND$MRkLMFk8
C8RRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRRMhFCR

RVRRk0MOHRFMp5mtZH:RMmRBv upXm_up;q)R1Aq H:RM R)q2pRR0sCkRsMBumvp_ Xuqmp)R;
RRRRR-RR-kRus#bFCR:
RRRRR-RR-RRRRRRRRCR)0Mks#sRbHHMObRNDPkNDCVRFRoDFN0sHELlRNR#CA q1RRFVZR
RRRRRR-R-RC1bODHNRDPNk:C#
RRRRRRRRR--RRRRRRRRp5mtZA,Rq21 RB=Rmpvu uX_m)pq'35jjj,R3Rj2HZVR3tvqR4=R3NjRMR8
RRRRR-RR-RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRqZ3)=tRRjj3
RRRRRRRRR--RRRRRRRRp5mtZA,Rq21 RB=Rmpvu uX_m)pq'354jj,R3Rj2HZVR3tvqRA=RqR1 N
M8RRRRRRRR-R-RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR3RZqR)t=3RjjR
RRRRRR-R-Rl7FN:HM
RRRRRRRRR--RRRRRRRRZMRHRvBmuXp _pumqN)RMZ8R3tq)RR/=-avq]Q_u
RRRRRRRRR--RRRRRRRRZq3vt=R/Rjj3
RRRRRRRRR--RRRRRRRRA q1Rj>R3Rj
RRRRR-RR-RRRRRRRRqRA1/ R=3R4jR
RRRRRR-R-Rs sFOsRFHM80MHF#R:
RRRRR-RR-RRRRRRRRsR sRFsHZVR3tq)R-=Rv]qa_
uQRRRRRRRR-R-RRRRRR RRsssFRRHVZq3vtRR=j
3jRRRRRRRR-R-RRRRRR RRsssFRRHVA q1RR<=j
3jRRRRRRRR-R-RRRRRR RRsssFRRHVA q1R4=R3Rj
RRRRR-RR-NR)M:oC
RRRRRRRRR--RRRRRRRRskC#Dv03q>tR=3RjjR
RRRRRR-R-RRRRRRRRRq-vau]_QRR<skC#Dq03)<tR=qRvau]_QR
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRRhRRF
MC
RRRRMVkOF0HMQR1hZR5RH:RMmRBv upXm_upRq)2CRs0MksRvBmuXp _pumq
);RRRRRRRR-u-RkFsb#
C:RRRRRRRR-R-RRRRRR)RRCs0kMb#RsOHMHDbNRDPNkFCRVHR#MFCRV
RZRRRRRRRR-1-RbHCONPDRNCDk#R:
RRRRR-RR-RRRRRRRRQR1h25ZRB=Rmpvu uX_m)pq'35jjj,R3Rj2HZVR3tvqRj=R3NjRMR8
RRRRR-RR-RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRqZ3)=tRRjj3
RRRRRRRRR--RRRRRRRR15QhZ=2RRvBmuXp _pumq5)'j,3jRjj32VRHRvZ3q=tRRavq]Q_uR8NM
RRRRRRRRR--RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRZRR3tq)Rj=R3Rj
RRRRR-RR-FR7lMNH:R
RRRRRR-R-RRRRRRRRRHZRMmRBv upXm_upRq)NRM8Z)3qt=R/Rq-vau]_QR
RRRRRR-R-Rs sFOsRFHM80MHF#R:
RRRRR-RR-RRRRRRRRsR sRFsHZVR3tq)R-=Rv]qa_
uQRRRRRRRR-)-RNCMo:R
RRRRRR-R-RRRRRRRRR#sCk3D0vRqt>j=R3Rj
RRRRR-RR-RRRRRRRRvR-q_a]u<QRR#sCk3D0qR)t<v=Rq_a]uRQ
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRRRRhCFM
R
RRkRVMHO0F1MRQ5hRZRR:HBMRmpvu 2XRR0sCkRsMBumvp; X
RRRRRRRRR--ubksF:#C
RRRRRRRRR--RRRRRRRR)kC0sRM##CHMRRFVZR
RRRRRR-R-RC1bODHNRDPNk:C#
RRRRRRRRR--RRRRRRRR15Qhv]qa_ BZ)Rm2=qRvaB]_Zm )
RRRRRRRRR--RRRRRRRR15QhZ=2RRavq]Z_B R)mHZVRRB=Rmpvu 5X'v]qa_,uQRjj32R
RRRRRR-R-Rl7FN:HM
RRRRRRRRR--RRRRRRRRZMRHRvBmuXp 
RRRRRRRRR-- FsssFROM08HH#FM:R
RRRRRR-R-RRRRRRRRRMhFCR
RRRRRR-R-RM)No
C:RRRRRRRR-R-RRRRRRqRRA115QZh52<2R=TR1)1a5QZh532) *h1Q5)Z3 +2R
RRRRRRRRR--RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR1]Qh5QZ3v12*Q5h]Zv3Q2R2
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRRRRhCFM
R
RRkRVMHO0FRMRBRm15:ZRRRHMBumvpR X2CRs0MksRvBmuXp ;R
RRRRRR-R-RsukbCF#:R
RRRRRR-R-RRRRRRRRR0)Ck#sMR#OFHRMCFZVR
RRRRRRRRR--1ObCHRNDPkNDC
#:RRRRRRRR-R-RRRRRRBRRmZ152RR=v]qa_ BZ)HmRVRRZ=mRBv upXv'5q_a]umQ_e_ ).j,R3
j2RRRRRRRR-R-RRRRRRBRRmZ152RR=v]qa_ BZ)HmRVRRZ=mRBv upX-'5v]qa__uQm)e _R.,j23j
RRRRRRRRR--7NFlH
M:RRRRRRRR-R-RRRRRRZRRRRHMBumvp
 XRRRRRRRR- -RsssFRMOF8HH0F:M#
RRRRRRRRR--RRRRRRRRhCFM
RRRRRRRRR--)oNMCR:
RRRRR-RR-RRRRRRRRARq1m5B125Z2=R<R)1Tam5B135Z)* 2B5m1Z 3)2
R+RRRRRRRR-R-RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR1RRQ5h]Zv3Q2Q*1hZ]532Qv2R
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRRhRRF
MC
R
RRkRVMHO0FRMRBRm15:ZRRRHMBumvp_ Xuqmp)RR2skC0sBMRmpvu uX_m)pq;R
RRRRRR-R-RsukbCF#:R
RRRRRR-R-RRRRRRRRR0)Ck#sMRHbsMbOHNPDRNCDkRRFVOHF#MFCRV
RZRRRRRRRR-1-RbHCONPDRNCDk#R:
RRRRR-RR-RRRRRRRRmRB125ZRB=Rmpvu uX_m)pq'35jjj,R3Rj2HZVR3tvqRv=Rq_a]umQ_e_ ).R
RRRRRR-R-RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRNRRMZ8R3tq)Rj=R3Rj
RRRRR-RR-RRRRRRRRmRB125ZRB=Rmpvu uX_m)pq'35jjj,R3Rj2HZVR3tvqRv=Rq_a]umQ_e_ ).R
RRRRRR-R-RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRNRRMZ8R3tq)Rv=Rq_a]uRQ
RRRRR-RR-FR7lMNH:R
RRRRRR-R-RRRRRRRRRHZRMmRBv upXm_upRq)NRM8Z)3qt=R/Rq-vau]_QR
RRRRRR-R-Rs sFOsRFHM80MHF#R:
RRRRR-RR-RRRRRRRRsR sRFsHZVR3tq)R-=Rv]qa_
uQRRRRRRRR-)-RNCMo:R
RRRRRR-R-RRRRRRRRR#sCk3D0vRqt>j=R3Rj
RRRRR-RR-RRRRRRRRvR-q_a]u<QRR#sCk3D0qR)t<v=Rq_a]uRQ
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRRRRhCFM
R
RRkRVMHO0F1MRQRh]5:ZRRRHMBumvpR X2CRs0MksRvBmuXp ;R
RRRRRR-R-RsukbCF#:R
RRRRRR-R-RRRRRRRRR0)Ck#sMRbE$CFsLDRHO#CHMRRFVZR
RRRRRR-R-RC1bODHNRDPNk:C#
RRRRRRRRR--RRRRRRRR1]Qh5avq]Z_B 2)mRv=Rq_a]B)Z mR
RRRRRR-R-RRRRRRRRRh1Q]25ZRv=Rq_a]B)Z mVRHR)Z3 RR=jR3jNRM8Zv3QRv=Rq_a]uRQ
RRRRR-RR-RRRRRRRRQR1hZ]52RR=v]qa_qBA1K _RRHVZ 3)Rj=R3NjRMR8
RRRRR-RR-RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRZv3QRv=Rq_a]umQ_e_ ).R
RRRRRR-R-RRRRRRRRRh1Q]25ZR-=Rv]qa_qBA1K _RRHVZ 3)Rj=R3NjRMR8
RRRRR-RR-RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRZv3QR-=Rv]qa__uQm)e _R.
RRRRR-RR-FR7lMNH:R
RRRRRR-R-RRRRRRRRRHZRMmRBv upXR
RRRRRR-R-Rs sFOsRFHM80MHF#R:
RRRRR-RR-RRRRRRRRFRhMRC
RRRRR-RR-NR)M:oC
RRRRRRRRR--RRRRRRRRq5A11]Qh52Z2RR<=1aT)5h1Q]35Z)* 21]Qh5)Z3 +2R
RRRRRRRRR--RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR15QhZv3Q2Q*1h35ZQ2v2
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRRFRhM
C
RRRRVOkM0MHFRh1Q]ZR5RH:RMmRBv upXm_upRq)2CRs0MksRvBmuXp _pumq
);RRRRRRRR-u-RkFsb#
C:RRRRRRRR-R-RRRRRR)RRCs0kMb#RsOHMHDbNRDPNkFCRV$REbLCsFODHRM#HCVRFRRZ
RRRRR-RR-bR1CNOHDNRPD#kC:R
RRRRRR-R-RRRRRRRRRh1Q]25ZRB=Rmpvu uX_m)pq'35jjj,R3Rj2HZVR3tvqRj=R3NjRMR8
RRRRR-RR-RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRqZ3)=tRRjj3
RRRRRRRRR--RRRRRRRR1]Qh5RZ2=mRBv upXm_up'q)5jj3,3RjjH2RV3RZvRqt=qRvau]_QMRN8R
RRRRRR-R-RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRZ)3qtRR=v]qa__uQm)e _R.
RRRRR-RR-RRRRRRRRQR1hZ]52RR=Bumvp_ Xuqmp)4'53Rj,v]qa__uQm)e _R.2HZVR3tvqRR=
RRRRR-RR-RRRRRRRRRRRRRRRRRRRRRRRRqRvau]_Qe_m .)_R8NMRqZ3)=tRRavq]Q_u_ me)
_.RRRRRRRR-R-RRRRRR1RRQ5h]Z=2RRvBmuXp _pumq5)'4,3jRq-vau]_Qe_m .)_2VRHRvZ3q=tR
RRRRRRRRR--RRRRRRRRRRRRRRRRRRRRRRRRv]qa__uQm)e _N.RMZ8R3tq)R-=Rv]qa__uQm)e _R.
RRRRR-RR-FR7lMNH:R
RRRRRR-R-RRRRRRRRRHZRMmRBv upXm_upRq)NRM8Z)3qt=R/Rq-vau]_QR
RRRRRR-R-Rs sFOsRFHM80MHF#R:
RRRRR-RR-RRRRRRRRsR sRFsHZVR3tq)R-=Rv]qa_
uQRRRRRRRR-)-RNCMo:R
RRRRRR-R-RRRRRRRRR#sCk3D0vRqt>j=R3Rj
RRRRR-RR-RRRRRRRRvR-q_a]u<QRR#sCk3D0qR)t<v=Rq_a]uRQ
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRRRRhCFM
R
RRkRVMHO0FBMRmR1]5:ZRRRHMBumvpR X2CRs0MksRvBmuXp ;R
RRRRRR-R-RsukbCF#:R
RRRRRR-R-RRRRRRRRR0)Ck#sMRbE$CFsLDRHOOHF#MFCRV
RZRRRRRRRR-1-RbHCONPDRNCDk#R:
RRRRR-RR-RRRRRRRRmRB1v]5q_a]B)Z m=2RRavq]A_Bq_1 4R
RRRRRR-R-RRRRRRRRR1Bm]25ZR-=Rv]qa_qBA14 _RRHVZ 3)Rj=R3NjRMZ8R3RQv=qRvau]_QR
RRRRRR-R-RRRRRRRRR1Bm]25ZRv=Rq_a]B)Z mVRHR)Z3 RR=jR3jNRM8Zv3QRv=Rq_a]umQ_e_ ).R
RRRRRR-R-RRRRRRRRR1Bm]25ZRv=Rq_a]B)Z mVRHR)Z3 RR=jR3jNRM8Zv3QR-=Rv]qa__uQm)e _R.
RRRRR-RR-FR7lMNH:R
RRRRRR-R-RRRRRRRRRHZRMmRBv upXR
RRRRRR-R-Rs sFOsRFHM80MHF#R:
RRRRR-RR-RRRRRRRRFRhMRC
RRRRR-RR-NR)M:oC
RRRRRRRRR--RRRRRRRRq5A1B]m152Z2RR<=1aT)5h1Q]35Z)* 21]Qh5)Z3 +2R
RRRRRRRRR--RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRB5m1Zv3Q2m*B135ZQ2v2
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRRFRhM
C

RRRRMVkOF0HMmRB15]RZRR:HBMRmpvu uX_m)pqRs2RCs0kMmRBv upXm_up;q)
RRRRRRRRR--ubksF:#C
RRRRRRRRR--RRRRRRRR)kC0sRM#bMsHONHbDNRPDRkCFEVR$sbCLHFDOFRO#CHMRRFVZR
RRRRRR-R-RC1bODHNRDPNk:C#
RRRRRRRRR--RRRRRRRRB]m15RZ2=mRBv upXm_up'q)5j43,3RjjH2RV3RZvRqt=3RjjMRN8R
RRRRRR-R-RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRZ)3qtRR=j
3jRRRRRRRR-R-RRRRRRBRRm51]Z=2RRvBmuXp _pumq5)'4,3jRavq]Q_u2VRHRvZ3q=tRRavq]Q_uR8NM
RRRRRRRRR--RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRZRR3tq)Rv=Rq_a]umQ_e_ ).R
RRRRRR-R-RRRRRRRRR1Bm]25ZRB=Rmpvu uX_m)pq'35jjj,R3Rj2HZVR3tvqRR=
RRRRR-RR-RRRRRRRRRRRRRRRRRRRRRRRRavq]Q_u_ me)R_.NRM8Z)3qtRR=v]qa__uQm)e _R.
RRRRR-RR-RRRRRRRRmRB1Z]52RR=Bumvp_ Xuqmp)j'53Rj,j23jRRHVZq3vt
R=RRRRRRRR-R-RRRRRRRRRRRRRRRRRRRRRRqRvau]_Qe_m .)_R8NMRqZ3)=tRRq-vau]_Qe_m .)_
RRRRRRRRR--7NFlH
M:RRRRRRRR-R-RRRRRRZRRRRHMBumvp_ Xuqmp)MRN83RZqR)t/-=Rv]qa_
uQRRRRRRRR- -RsssFRMOF8HH0F:M#
RRRRRRRRR--RRRRRRRR FsssVRHRqZ3)=tRRq-vau]_QR
RRRRRR-R-RM)No
C:RRRRRRRR-R-RRRRRRsRRCD#k0q3vt=R>Rjj3
RRRRRRRRR--RRRRRRRR-avq]Q_uRs<RCD#k0)3qt=R<Ravq]Q_u
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRRFRhM
C
RRRR-R-
R-RR-sRqHl0ECO0HRCmbsFN0sR#
R-RR-R

RVRRk0MOHRFM"R+"5:RpRRHMBumvp; XR:R)RRHMBumvpR X2CRs0MksRvBmuXp ;R
RRRRRR-R-RsukbCF#:R
RRRRRR-R-RRRRRRRRR0)Ck#sMRHNs0CEl0RHONH880MHFRRFVpMRN8
R)RRRRRRRR-1-RbHCONPDRNCDk#R:
RRRRR-RR-RRRRRRRRFRhMRC
RRRRR-RR-FR7lMNH:R
RRRRRR-R-RRRRRRRRRHpRMmRBv upXR
RRRRRR-R-RRRRRRRRRH)RMmRBv upXR
RRRRRR-R-Rs sFOsRFHM80MHF#R:
RRRRR-RR-RRRRRRRRFRhMRC
RRRRR-RR-NR)M:oC
RRRRRRRRR--RRRRRRRR"5+"ZH2R#NRl0lECNO0HN$DDRLkMF8kMCR8
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRRRRhCFM
R
RRkRVMHO0F"MR+5"RRRp:H)MR ;qpRRRRRR):HBMRmpvu 2XRR0sCkRsMBumvp; X
RRRRRRRRR--ubksF:#C
RRRRRRRRR--RRRRRRRR)kC0sRM#N0sHE0lCHNOR808HHRFMFpVRR8NMRR)
RRRRR-RR-bR1CNOHDNRPD#kC:R
RRRRRR-R-RRRRRRRRRMhFCR
RRRRRR-R-Rl7FN:HM
RRRRRRRRR--RRRRRRRRpMRHRq) pR
RRRRRR-R-RRRRRRRRRH)RMmRBv upXR
RRRRRR-R-Rs sFOsRFHM80MHF#R:
RRRRR-RR-RRRRRRRRFRhMRC
RRRRR-RR-NR)M:oC
RRRRRRRRR--RRRRRRRR"5+"ZH2R#NRl0lECNO0HN$DDRLkMF8kMCR8
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRRRRhCFM
R
RRkRVMHO0F"MR+5"RRRp:HBMRmpvu uX_m)pq;:R)RRHMBumvp_ Xuqmp)R2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRsRRCs0kMmRBv upXm_up;q)
RRRRRRRRR--ubksF:#C
RRRRRRRRR--RRRRRRRR)kC0sRM#N0sHE0lCHNOR808HHRFMFpVRR8NMRR)
RRRRR-RR-bR1CNOHDNRPD#kC:R
RRRRRR-R-RRRRRRRRRMhFCR
RRRRRR-R-Rl7FN:HM
RRRRRRRRR--RRRRRRRRpMRHRvBmuXp _pumqN)RMp8R3tq)RR/=-avq]Q_u
RRRRRRRRR--RRRRRRRR)MRHRvBmuXp _pumqN)RM)8R3tq)RR/=-avq]Q_u
RRRRRRRRR-- FsssFROM08HH#FM:R
RRRRRR-R-RRRRRRRRRs sFHsRV3RpqR)t=vR-q_a]uRQ
RRRRR-RR-RRRRRRRRsR sRFsH)VR3tq)R-=Rv]qa_
uQRRRRRRRR-)-RNCMo:R
RRRRRR-R-RRRRRRRRR#sCk3D0vRqt>j=R3Rj
RRRRR-RR-RRRRRRRRvR-q_a]u<QRR#sCk3D0qR)t<v=Rq_a]uRQ
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRRRRhCFM
R

RVRRk0MOHRFM"R+"5:RpRRHMBumvp; XR:R)RRHM)p qRR2RRCRs0MksRvBmuXp ;R
RRRRRR-R-RsukbCF#:R
RRRRRR-R-RRRRRRRRR0)Ck#sMRHNs0CEl0RHONH880MHFRRFVpMRN8
R)RRRRRRRR-1-RbHCONPDRNCDk#R:
RRRRR-RR-RRRRRRRRFRhMRC
RRRRR-RR-FR7lMNH:R
RRRRRR-R-RRRRRRRRRHpRMmRBv upXR
RRRRRR-R-RRRRRRRRRH)RM R)qRp
RRRRR-RR-sR sRFsO8FMHF0HM
#:RRRRRRRR-R-RRRRRRhRRF
MCRRRRRRRR-)-RNCMo:R
RRRRRR-R-RRRRRRRRR""+5RZ2Hl#RNC0ElHN0ODND$MRkLMFk8
C8RRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRRMhFCR

RVRRk0MOHRFM"R+"5:RpRRHMBumvp_ Xuqmp)R;R)H:RM R)qRp2skC0sBMRmpvu uX_m)pq;R
RRRRRR-R-RsukbCF#:R
RRRRRR-R-RRRRRRRRR0)Ck#sMRHNs0CEl0RHONH880MHFRRFVpMRN8
R)RRRRRRRR-1-RbHCONPDRNCDk#R:
RRRRR-RR-RRRRRRRRFRhMRC
RRRRR-RR-FR7lMNH:R
RRRRRR-R-RRRRRRRRRHpRMmRBv upXm_upRq)NRM8p)3qt=R/Rq-vau]_QR
RRRRRR-R-RRRRRRRRRH)RM R)qRp
RRRRR-RR-sR sRFsO8FMHF0HM
#:RRRRRRRR-R-RRRRRR RRsssFRRHVp)3qtRR=-avq]Q_u
RRRRRRRRR--)oNMCR:
RRRRR-RR-RRRRRRRRCRs#0kD3tvqRR>=j
3jRRRRRRRR-R-RRRRRR-RRv]qa_RuQ<CRs#0kD3tq)RR<=v]qa_
uQRRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRRMhFCR

RVRRk0MOHRFM"R+"5:RpRRHM)p q;)RR:MRHRvBmuXp _pumqR)2skC0sBMRmpvu uX_m)pq;R
RRRRRR-R-RsukbCF#:R
RRRRRR-R-RRRRRRRRR0)Ck#sMRHNs0CEl0RHONH880MHFRRFVpMRN8
R)RRRRRRRR-1-RbHCONPDRNCDk#R:
RRRRR-RR-RRRRRRRRFRhMRC
RRRRR-RR-FR7lMNH:R
RRRRRR-R-RRRRRRRRRHpRM R)qRp
RRRRR-RR-RRRRRRRRRR)HBMRmpvu uX_m)pqR8NMRq)3)/tR=vR-q_a]uRQ
RRRRR-RR-sR sRFsO8FMHF0HM
#:RRRRRRRR-R-RRRRRR RRsssFRRHV))3qtRR=-avq]Q_u
RRRRRRRRR--)oNMCR:
RRRRR-RR-RRRRRRRRCRs#0kD3tvqRR>=j
3jRRRRRRRR-R-RRRRRR-RRv]qa_RuQ<CRs#0kD3tq)RR<=v]qa_
uQRRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRRMhFCR

RVRRk0MOHRFM"R-"5:RpRRHM)p q;RRRR:R)RRHMBumvpR X2CRs0MksRvBmuXp ;R
RRRRRR-R-RsukbCF#:R
RRRRRR-R-RRRRRRRRR0)Ck#sMRHNs0CEl0RHO#0kLs0NOHRFMFpVRRMlHk)#R
RRRRRRRRR--1ObCHRNDPkNDC
#:RRRRRRRR-R-RRRRRRhRRF
MCRRRRRRRR-7-RFHlNMR:
RRRRR-RR-RRRRRRRRRRpH)MR 
qpRRRRRRRR-R-RRRRRR)RRRRHMBumvp
 XRRRRRRRR- -RsssFRMOF8HH0F:M#
RRRRRRRRR--RRRRRRRRhCFM
RRRRRRRRR--)oNMCR:
RRRRR-RR-RRRRRRRR-R""25ZRRH#lEN0C0lNHDONDk$RMkLFM88C
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRRFRhM
C
RRRRVOkM0MHFR""-Rp5R:MRHRvBmuXp ;)RR:MRHRvBmuXp Rs2RCs0kMmRBv upXR;
RRRRR-RR-kRus#bFCR:
RRRRR-RR-RRRRRRRRCR)0Mks#sRNHl0ECO0HRL#k0OsN0MHFRRFVpHRlMRk#)R
RRRRRR-R-RC1bODHNRDPNk:C#
RRRRRRRRR--RRRRRRRRhCFM
RRRRRRRRR--7NFlH
M:RRRRRRRR-R-RRRRRRpRRRRHMBumvp
 XRRRRRRRR-R-RRRRRR)RRRRHMBumvp
 XRRRRRRRR- -RsssFRMOF8HH0F:M#
RRRRRRRRR--RRRRRRRRhCFM
RRRRRRRRR--)oNMCR:
RRRRR-RR-RRRRRRRR-R""25ZRRH#lEN0C0lNHDONDk$RMkLFM88C
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRRFRhM
C
RRRRVOkM0MHFR""-Rp5R:MRHRvBmuXp ;)RR:MRHRq) pRR2RsRRCs0kMmRBv upXR;
RRRRR-RR-kRus#bFCR:
RRRRR-RR-RRRRRRRRCR)0Mks#sRNHl0ECO0HRL#k0OsN0MHFRRFVpHRlMRk#)R
RRRRRR-R-RC1bODHNRDPNk:C#
RRRRRRRRR--RRRRRRRRhCFM
RRRRRRRRR--7NFlH
M:RRRRRRRR-R-RRRRRRpRRRRHMBumvp
 XRRRRRRRR-R-RRRRRR)RRRRHM)p q
RRRRRRRRR-- FsssFROM08HH#FM:R
RRRRRR-R-RRRRRRRRRMhFCR
RRRRRR-R-RM)No
C:RRRRRRRR-R-RRRRRR"RR-Z"52#RHR0lNENCl0NHODRD$kFMLkCM88R
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRRhRRF
MC
RRRRMVkOF0HM-R""RR5pH:RM R)qRp;RR):HBMRmpvu uX_m)pq2CRs0MksRvBmuXp _pumq
);RRRRRRRR-u-RkFsb#
C:RRRRRRRR-R-RRRRRR)RRCs0kMN#RsEH0lHC0OkR#LN0sOF0HMVRFRlpRH#MkRR)
RRRRR-RR-bR1CNOHDNRPD#kC:R
RRRRRR-R-RRRRRRRRRMhFCR
RRRRRR-R-Rl7FN:HM
RRRRRRRRR--RRRRRRRRpMRHRq) pR
RRRRRR-R-RRRRRRRRRH)RMmRBv upXm_upRq)NRM8))3qt=R/Rq-vau]_QR
RRRRRR-R-Rs sFOsRFHM80MHF#R:
RRRRR-RR-RRRRRRRRsR sRFsH)VR3tq)R-=Rv]qa_
uQRRRRRRRR-)-RNCMo:R
RRRRRR-R-RRRRRRRRR#sCk3D0vRqt>j=R3Rj
RRRRR-RR-RRRRRRRRvR-q_a]u<QRR#sCk3D0qR)t<v=Rq_a]uRQ
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRRRRhCFM
R

RVRRk0MOHRFM"R-"5:RpRRHMBumvp_ Xuqmp));R:MRHRvBmuXp _pumq
)2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRskC0sBMRmpvu uX_m)pq;R
RRRRRR-R-RsukbCF#:R
RRRRRR-R-RRRRRRRRR0)Ck#sMRHNs0CEl0RHO#0kLs0NOHRFMFpVRRMlHk)#R
RRRRRRRRR--1ObCHRNDPkNDC
#:RRRRRRRR-R-RRRRRRhRRF
MCRRRRRRRR-7-RFHlNMR:
RRRRR-RR-RRRRRRRRRRpHBMRmpvu uX_m)pqR8NMRqp3)/tR=vR-q_a]uRQ
RRRRR-RR-RRRRRRRRRR)HBMRmpvu uX_m)pqR8NMRq)3)/tR=vR-q_a]uRQ
RRRRR-RR-sR sRFsO8FMHF0HM
#:RRRRRRRR-R-RRRRRR RRsssFRRHVp)3qtRR=-avq]Q_u
RRRRRRRRR--RRRRRRRR FsssVRHRq)3)=tRRq-vau]_QR
RRRRRR-R-RM)No
C:RRRRRRRR-R-RRRRRRsRRCD#k0q3vt=R>Rjj3
RRRRRRRRR--RRRRRRRR-avq]Q_uRs<RCD#k0)3qt=R<Ravq]Q_u
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRRFRhM
C
RRRRVOkM0MHFR""-Rp5R:MRHRvBmuXp _pumqR);RR):H)MR 2qpR0sCkRsMBumvp_ Xuqmp)R;
RRRRR-RR-kRus#bFCR:
RRRRR-RR-RRRRRRRRCR)0Mks#sRNHl0ECO0HRL#k0OsN0MHFRRFVpHRlMRk#)R
RRRRRR-R-RC1bODHNRDPNk:C#
RRRRRRRRR--RRRRRRRRhCFM
RRRRRRRRR--7NFlH
M:RRRRRRRR-R-RRRRRRpRRRRHMBumvp_ Xuqmp)MRN83RpqR)t/-=Rv]qa_
uQRRRRRRRR-R-RRRRRR)RRRRHM)p q
RRRRRRRRR-- FsssFROM08HH#FM:R
RRRRRR-R-RRRRRRRRRs sFHsRV3RpqR)t=vR-q_a]uRQ
RRRRR-RR-NR)M:oC
RRRRRRRRR--RRRRRRRRskC#Dv03q>tR=3RjjR
RRRRRR-R-RRRRRRRRRq-vau]_QRR<skC#Dq03)<tR=qRvau]_QR
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRRhRRF
MC
RRRRMVkOF0HM*R""RR5pH:RMmRBv upXR;R)H:RMmRBv upXRR2skC0sBMRmpvu 
X;RRRRRRRR-u-RkFsb#
C:RRRRRRRR-R-RRRRRR)RRCs0kMN#RsEH0lHC0OkRlDb0HDNHO0MHFRRFVpMRN8
R)RRRRRRRR-1-RbHCONPDRNCDk#R:
RRRRR-RR-RRRRRRRRFRhMRC
RRRRR-RR-FR7lMNH:R
RRRRRR-R-RRRRRRRRRHpRMmRBv upXR
RRRRRR-R-RRRRRRRRRH)RMmRBv upXR
RRRRRR-R-Rs sFOsRFHM80MHF#R:
RRRRR-RR-RRRRRRRRFRhMRC
RRRRR-RR-NR)M:oC
RRRRRRRRR--RRRRRRRR"5*"ZH2R#NRl0lECNO0HN$DDRLkMF8kMCR8
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRRRRhCFM
R
RRkRVMHO0F"MR*5"RRRp:HBMRmpvu RX;RR):H)MR Rqp2sRRCs0kMmRBv upXR;
RRRRR-RR-kRus#bFCR:
RRRRR-RR-RRRRRRRRCR)0Mks#sRNHl0ECO0HRDlk0DHbH0ONHRFMFpVRR8NMRR)
RRRRR-RR-bR1CNOHDNRPD#kC:R
RRRRRR-R-RRRRRRRRRMhFCR
RRRRRR-R-Rl7FN:HM
RRRRRRRRR--RRRRRRRRpMRHRvBmuXp 
RRRRRRRRR--RRRRRRRR)MRHRq) pR
RRRRRR-R-Rs sFOsRFHM80MHF#R:
RRRRR-RR-RRRRRRRRFRhM
C
RRRRRRRR-)-RNCMo:R
RRRRRR-R-RRRRRRRRR""*5RZ2Hl#RNC0ElHN0ODND$MRkLMFk8
C8RRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRRMhFCR

RVRRk0MOHRFM"R*"5:RpRRHM)p q;)RR:MRHRvBmuXp Rs2RCs0kMmRBv upXR;
RRRRR-RR-kRus#bFCR:
RRRRR-RR-RRRRRRRRCR)0Mks#sRNHl0ECO0HRDlk0DHbH0ONHRFMFpVRR8NMRR)
RRRRR-RR-bR1CNOHDNRPD#kC:R
RRRRRR-R-RRRRRRRRRMhFCR
RRRRRR-R-Rl7FN:HM
RRRRRRRRR--RRRRRRRRpMRHRq) pR
RRRRRR-R-RRRRRRRRRH)RMmRBv upXR
RRRRRR-R-Rs sFOsRFHM80MHF#R:
RRRRR-RR-RRRRRRRRFRhMRC
RRRRR-RR-NR)M:oC
RRRRRRRRR--RRRRRRRR"5*"ZH2R#NRl0lECNO0HN$DDRLkMF8kMCR8
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRRRRhCFM
R
RRkRVMHO0F"MR*5"RRRp:HBMRmpvu uX_m)pq;:R)RRHMBumvp_ Xuqmp)R2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRsRRCs0kMmRBv upXm_up;q)
RRRRRRRRR--ubksF:#C
RRRRRRRRR--RRRRRRRR)kC0sRM#N0sHE0lCHlORkHD0bODHNF0HMVRFRNpRM)8R
RRRRRRRRR--1ObCHRNDPkNDC
#:RRRRRRRR-R-RRRRRRhRRF
MCRRRRRRRR-7-RFHlNMR:
RRRRR-RR-RRRRRRRRRRpHBMRmpvu uX_m)pqR8NMRqp3)/tR=vR-q_a]uRQ
RRRRR-RR-RRRRRRRRRR)HBMRmpvu uX_m)pqR8NMRq)3)/tR=vR-q_a]uRQ
RRRRR-RR-sR sRFsO8FMHF0HM
#:RRRRRRRR-R-RRRRRR RRsssFRRHVp)3qtRR=-avq]Q_u
RRRRRRRRR--RRRRRRRR FsssVRHRq)3)=tRRq-vau]_QR
RRRRRR-R-RM)No
C:RRRRRRRR-R-RRRRRRsRRCD#k0q3vt=R>Rjj3
RRRRRRRRR--RRRRRRRR-avq]Q_uRs<RCD#k0)3qt=R<Ravq]Q_u
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRRFRhM
C
RRRRVOkM0MHFR""*Rp5R:MRHRq) pR;R)H:RMmRBv upXm_up2q)R0sCkRsMBumvp_ Xuqmp)R;
RRRRR-RR-kRus#bFCR:
RRRRR-RR-RRRRRRRRCR)0Mks#sRNHl0ECO0HRDlk0DHbH0ONHRFMFpVRR8NMRR)
RRRRR-RR-bR1CNOHDNRPD#kC:R
RRRRRR-R-RRRRRRRRRMhFCR
RRRRRR-R-Rl7FN:HM
RRRRRRRRR--RRRRRRRRpMRHRq) pR
RRRRRR-R-RRRRRRRRRH)RMmRBv upXm_upRq)NRM8))3qt=R/Rq-vau]_QR
RRRRRR-R-Rs sFOsRFHM80MHF#R:
RRRRR-RR-RRRRRRRRsR sRFsH)VR3tq)R-=Rv]qa_
uQRRRRRRRR-)-RNCMo:R
RRRRRR-R-RRRRRRRRR#sCk3D0vRqt>j=R3Rj
RRRRR-RR-RRRRRRRRvR-q_a]u<QRR#sCk3D0qR)t<v=Rq_a]uRQ
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRRRRhCFM
R
RRkRVMHO0F"MR*5"RRRp:HBMRmpvu uX_m)pq;)RR:MRHRq) ps2RCs0kMmRBv upXm_up;q)
RRRRRRRRR--ubksF:#C
RRRRRRRRR--RRRRRRRR)kC0sRM#N0sHE0lCHlORkHD0bODHNF0HMVRFRNpRM)8R
RRRRRRRRR--1ObCHRNDPkNDC
#:RRRRRRRR-R-RRRRRRhRRF
MCRRRRRRRR-7-RFHlNMR:
RRRRR-RR-RRRRRRRRRRpHBMRmpvu uX_m)pqR8NMRqp3)/tR=vR-q_a]uRQ
RRRRR-RR-RRRRRRRRRR)H)MR 
qpRRRRRRRR- -RsssFRMOF8HH0F:M#
RRRRRRRRR--RRRRRRRR FsssVRHRqp3)=tRRq-vau]_QR
RRRRRR-R-RM)No
C:RRRRRRRR-R-RRRRRRsRRCD#k0q3vt=R>Rjj3
RRRRRRRRR--RRRRRRRR-avq]Q_uRs<RCD#k0)3qt=R<Ravq]Q_u
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRRFRhM
C

RRRRMVkOF0HM/R""RR5pH:RM R)qRp;RR):HBMRmpvu 2XRR0sCkRsMBumvp; X
RRRRRRRRR--ubksF:#C
RRRRRRRRR--RRRRRRRR)kC0sRM#N0sHE0lCH8ORH#PHHRFMFpVRRRL$)R
RRRRRR-R-RC1bODHNRDPNk:C#
RRRRRRRRR--RRRRRRRRhCFM
RRRRRRRRR--7NFlH
M:RRRRRRRR-R-RRRRRRpRRRRHM)p q
RRRRRRRRR--RRRRRRRR)MRHRvBmuXp R8NMR/)R=qRvaB]_Zm )
RRRRRRRRR-- FsssFROM08HH#FM:R
RRRRRR-R-RRRRRRRRRs sFHsRVRR)=qRvaB]_Zm )
RRRRRRRRR--)oNMCR:
RRRRR-RR-RRRRRRRR/R""25ZRRH#lEN0C0lNHDONDk$RMkLFM88C
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRRFRhM
C
RRRRVOkM0MHFR""/Rp5R:MRHRvBmuXp ;)RR:MRHRvBmuXp Rs2RCs0kMmRBv upXR;
RRRRR-RR-kRus#bFCR:
RRRRR-RR-RRRRRRRRCR)0Mks#sRNHl0ECO0HRP8HHF#HMVRFRLpR$
R)RRRRRRRR-1-RbHCONPDRNCDk#R:
RRRRR-RR-RRRRRRRRFRhMRC
RRRRR-RR-FR7lMNH:R
RRRRRR-R-RRRRRRRRRHpRMmRBv upXR
RRRRRR-R-RRRRRRRRRH)RMmRBv upXMRN8RR)/v=Rq_a]B)Z mR
RRRRRR-R-Rs sFOsRFHM80MHF#R:
RRRRR-RR-RRRRRRRRsR sRFsH)VRRv=Rq_a]B)Z mR
RRRRRR-R-RM)No
C:RRRRRRRR-R-RRRRRR"RR/Z"52#RHR0lNENCl0NHODRD$kFMLkCM88R
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRRhRRF
MC
RRRRMVkOF0HM/R""RR5pH:RMmRBv upXR;R)H:RM R)q2pRRRRRskC0sBMRmpvu 
X;RRRRRRRR-u-RkFsb#
C:RRRRRRRR-R-RRRRRR)RRCs0kMN#RsEH0lHC0OHR8PHH#FFMRVRRpL)$R
RRRRRRRRR--1ObCHRNDPkNDC
#:RRRRRRRR-R-RRRRRRhRRF
MCRRRRRRRR-7-RFHlNMR:
RRRRR-RR-RRRRRRRRRRpHBMRmpvu RX
RRRRR-RR-RRRRRRRRRR)H)MR RqpNRM8)=R/Rjj3
RRRRRRRRR-- FsssFROM08HH#FM:R
RRRRRR-R-RRRRRRRRRs sFHsRVRR)=3RjjR
RRRRRR-R-RM)No
C:RRRRRRRR-R-RRRRRR"RR/Z"52#RHR0lNENCl0NHODRD$kFMLkCM88R
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRRhRRF
MC
RRRRMVkOF0HM/R""RR5pH:RMmRBv upXm_up;q)RR):HBMRmpvu uX_m)pq2R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRCRs0MksRvBmuXp _pumq
);RRRRRRRR-u-RkFsb#
C:RRRRRRRR-R-RRRRRR)RRCs0kMN#RsEH0lHC0OHR8PHH#FFMRVRRpL)$R
RRRRRRRRR--1ObCHRNDPkNDC
#:RRRRRRRR-R-RRRRRRhRRF
MCRRRRRRRR-7-RFHlNMR:
RRRRR-RR-RRRRRRRRRRpHBMRmpvu uX_m)pqR8NMRqp3)/tR=vR-q_a]uRQ
RRRRR-RR-RRRRRRRRRR)HBMRmpvu uX_m)pqR8NMRq)3)/tR=vR-q_a]uRQ
RRRRR-RR-RRRRRRRR3R)vRqt>3RjjR
RRRRRR-R-Rs sFOsRFHM80MHF#R:
RRRRR-RR-RRRRRRRRsR sRFsH)VR3tvqRR<=j
3jRRRRRRRR-R-RRRRRR RRsssFRRHVp)3qtRR=-avq]Q_u
RRRRRRRRR--RRRRRRRR FsssVRHRq)3)=tRRq-vau]_QR
RRRRRR-R-RM)No
C:RRRRRRRR-R-RRRRRRsRRCD#k0q3vt=R>Rjj3
RRRRRRRRR--RRRRRRRR-avq]Q_uRs<RCD#k0)3qt=R<Ravq]Q_u
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRRFRhM
C
RRRRVOkM0MHFR""/Rp5R:MRHRq) pR;R)H:RMmRBv upXm_up2q)R0sCkRsMBumvp_ Xuqmp)R;
RRRRR-RR-kRus#bFCR:
RRRRR-RR-RRRRRRRRCR)0Mks#sRNHl0ECO0HRP8HHF#HMVRFRLpR$
R)RRRRRRRR-1-RbHCONPDRNCDk#R:
RRRRR-RR-RRRRRRRRFRhMRC
RRRRR-RR-FR7lMNH:R
RRRRRR-R-RRRRRRRRRHpRM R)qRp
RRRRR-RR-RRRRRRRRRR)HBMRmpvu uX_m)pqR8NMRq)3)/tR=vR-q_a]uRQ
RRRRR-RR-RRRRRRRR3R)vRqt>3RjjR
RRRRRR-R-Rs sFOsRFHM80MHF#R:
RRRRR-RR-RRRRRRRRsR sRFsH)VR3tvqRR<=j
3jRRRRRRRR-R-RRRRRR RRsssFRRHV))3qtRR=-avq]Q_u
RRRRRRRRR--)oNMCR:
RRRRR-RR-RRRRRRRRCRs#0kD3tvqRR>=j
3jRRRRRRRR-R-RRRRRR-RRv]qa_RuQ<CRs#0kD3tq)RR<=v]qa_
uQRRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRRMhFCR

RVRRk0MOHRFM"R/"5:RpRRHMBumvp_ Xuqmp)R;R)H:RM R)qRp2skC0sBMRmpvu uX_m)pq;R
RRRRRR-R-RsukbCF#:R
RRRRRR-R-RRRRRRRRR0)Ck#sMRHNs0CEl0RHO8HHP#MHFRRFVp$RLRR)
RRRRR-RR-bR1CNOHDNRPD#kC:R
RRRRRR-R-RRRRRRRRRMhFCR
RRRRRR-R-Rl7FN:HM
RRRRRRRRR--RRRRRRRRpMRHRvBmuXp _pumqN)RMp8R3tq)RR/=-avq]Q_u
RRRRRRRRR--RRRRRRRR)=R/Rjj3
RRRRRRRRR-- FsssFROM08HH#FM:R
RRRRRR-R-RRRRRRRRRs sFHsRV3RpqR)t=vR-q_a]uRQ
RRRRR-RR-RRRRRRRRsR sRFsH)VRRj=R3Rj
RRRRR-RR-NR)M:oC
RRRRRRRRR--RRRRRRRRskC#Dv03q>tR=3RjjR
RRRRRR-R-RRRRRRRRRq-vau]_QRR<skC#Dq03)<tR=qRvau]_QR
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRRhRRF
MCCRM8Ravq]m_Bv upX-;
---------------------------------------------------------------------
-----
-FRBbH$soRE04nggRRL$Q   3DRqDHRso#E0R#sCCCsP8-3
--
-RHaE#FR#kCsORDVHC#RHRRNMHFMVs0lNHRPCb0NsRRFVQ   R810R(4jn-3.4ngg, RQ 1 R08NMNRs8
R--ep]7R0vNENCl0NHODNRuOo	NCR#3a#EHRk#FsROCVCHDR$lNR0MFRRLCOHFbCR8,#8FD,sRFR-
-ROHMDCk88HRI0#ERFIV0NRsC00ENRRH##8FDR0IHE0FkRHIs0M0CRsbCl#H#HRFMVlsFRC0ER Q  -
-RN10Ms8N87#RCsbN0MlC0a3RERH##sFkOVCRHRDClRN$LkCR#RC80HFRlCbDl0CMRH0E#0R#NNM8s
8R-N-RMl8RNL$RCHR8#H0sLCk08MRHRlOFbCHD8FRVsHlRMMRN$NRlMsMCRR#FDoFMRRN#0REC
R--ObFlH8DCRsVFlFR8CM#RFN0RDIDFRs8HCRO08FCOlDbHNF0HMVRFRC0ERHFsoNHMDFR#kCsORDVHC-3
-ERaH##RFOksCHRVDlCRNL$RCFROb8HCRsVFR8HMH8PHkRNDkR#CLIC0CRCMDCHOM8#CRCk#sR#3
R--a#EHRk#FsROCVCHDRRH#bPsFH88CRRFMNqMR11RQR#LNHR#3aRECQ   R#8HOHDNlq#Rh
YR-W-Rqq))hRaY )Xu R11mQ)RvQup Q7RhzBp7tQhRYqhR)Wq)aqhYwRmR)v Bh]qaQqApYQaR-
-R7qhRawQh1 1R)wmR z1R)wmRuqRqQ)aBqzp)zRu)1um a3REkCR#RCsF0VRE#CRFOksC-R
-HRVD#CREDNDR8HMCHlMVN$RME8RFRD8Q   RsENl#DC#sRVFNlRM8$RNolNCF#RsHRDNDLHHR0$
R--N#sHHRMoFRk0F0VREkCR#0CRECCsF
V3---
-HRa0:DCRRRRR1RR08NMNRs8ep]7R0vNENCl0NHODNRuOo	NC5#RQ   R810R(4jn-3.4ngg,-
-RRRRRRRRRRRRRqRvaB]_mpvu 
X2---
-HRpLssN$R:RRaRRERH#b	NONRoC#DENDCRLRlOFbCHD8MRH0NFRRLDHs$Ns
R--RRRRRRRRRRRRRl#$LHFDODND$NRMlRC8Q   3-
-
R--7CCPDCFbsR#:R Q  qR71eBR]R7pvEN0C0lNHDONROuN	CNo#FRWsM	HosRtF
kb---
-kRus#bFCR:RRaRRERH#b	NONRoCL$F8RRH#NFRMMsMFlHN0PHCRlCbDl0CMNF0HMVRFRC0ER-
-RRRRRRRRRRRRRkRVMHO0FDMNHR0$8HCVMRC8H0MREvCRq_a]BumvpR Xb	NONRoC8DCON0sNH3FM

---p-RH0lHNF0HMR:RaRECPkNDCo#RCsMCN80CRRL$0RECVOkM0MHF#MRHRH0E#NRbOo	NCNRl$-
-RRRRRRRRRRRRRNRPsV$RsRFlb0DNVlFsRR0Fb0DNVlFs,MRN8ER0CsRbC#OHHRFMFsVRCD#k0-#
-RRRRRRRRRRRRHRR#MRFDo$RkNNsMC0C8FR0RRLC0REClHHMlRklskCJH8sCRRL$Q   R810R(4jn-
-RRRRRRRRRRRRR4R-g3gd

---h-RF#0C:-
-RRRRRRRRRRRRRERaCbR"NNO	o8CRCNODsHN0FRM"8HCVMRC#0REC0C$b##,Rk$L0b,C#R8NM
R--RRRRRRRRRRRRRO8CDNNs0MHF#VRFRavq]m_Bv upX-3
-RRRRRRRRRRRRaRRE#CR08NMNRs8lEN0C0lNHDONRV8CH0MHHRFMNRM8OPFMCHM0FDMNRNlCMoHM
R--RRRRRRRRRRRRRRFV0REClEN0C0lNHDONRMVkOF0HM0#RERN0NRsCb0NsRRFV0#EHRN#0Ms8N8-
-RRRRRRRRRRRRRCRsb#sCCRM00RECVlFsN#DRCMlN0#HORRFV0RECHDlbCMlC0HN0FFMRVER0C-
-RRRRRRRRRRRRRqRvaB]_mpvu bXRNNO	o8CRCNODsHN0FRM3RCaERsbkbCF#RRFV0
EC-R-RRRRRRRRRRRRRv]qa_vBmuXp RObN	CNoR8LF$#RHRR0FOsDNHRV$#EkORl#CNHM0ON#RM-8
-RRRRRRRRRRRRbRRsHFP8NCRRHok8HCDMVCRFHsRlCbDl0CMNF0HM0#RFCRPs$HVRC0EH-s
-RRRRRRRRRRRRHRRlCbDl0CMNF0HMVRFRavq]m_Bv upXR3RaDFFRP8CCbDFCRs#lRN$OFEF#0CRF-
-RRRRRRRRRRRRRlRHblDCCRM00RECb	NONRoCL$F8RRHM0RECl0F#RVCVHCOHMl0RNCMMs-
-RRRRRRRRRRRRRPRNNNHDLRDC00FRE3Cl

-----R----------------------------------------------------------------------------
R--e#CsHRFMR:RRR643
R--7CN0RRRRR:RRRR.cK$kDRg4gn-
-R----------------------------------------------------------------------------
-
kR#CWim)3avq] _)qNp3D
D;
ObN	CNoR8LF$qRvaB]_mpvu HXR#R

R-RR-R
RR-R-Rk JN0DH$MRN8MRQCNJkD$H0RCmbsFN0sV#RFBsRmpvu uX_m)pq
RRRR
--RRRRVOkM0MHFR""=Rp5R:MRHRvBmuXp _pumqR);RR):HBMRmpvu uX_m)pqRs2RCs0kMmRAmqp hR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRHRR#R
RRRRRR-R-R#7CObsH0MHF:R
RRRRRR-R-RRRRRRRR1RCCVOkM0MHFRO8CDNNs0MHFRRHMQ   R810R(4jn-3.4ngg
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRRRN2)kC0sRM#w1qp MRFRsCsFRs
RLRRCMoH
RRRRRRRRR--BOEC	NRPDHH80F$RVMRHbRk0Nksol0CM#R
RRRRRRVRHRp5R3tq)R-=Rv]qa_RuQ2ER0CRM
RRRRRRRRRRRRRNRR#s#C0qRwp
1 RRRRRRRRRRRRRRRRRRRRRRRRRRRRsFCbs"0Rp)3qtRR=-avq]Q_uRRHM=,5p)
2"RRRRRRRRRRRRRRRRRRRRRRRRRRRR#CCPs$H0R) )m
);RRRRRRRRRRRRRRRRskC0swMRq p1;R
RRRRRRMRC8VRH;R

RRRRRHRRVRR5))3qtRR=-avq]Q_uR02RE
CMRRRRRRRRRRRRRRRRNC##sw0Rq p1
RRRRRRRRRRRRRRRRRRRRRRRRRRRRbsCFRs0"q)3)=tRRq-vau]_QMRHRp=5,")2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRP#CC0sH$)R );m)
RRRRRRRRRRRRRRRR0sCkRsMw1qp R;
RRRRRCRRMH8RV
;
RRRRRRRR-t-RC#0RbHCONPDRNCDk#R
RRRRRRVRHRp5R3tvqRj=R3NjRM)8R3tvqRj=R32jRRC0EMR
RRRRRRRRRRRRRRCRs0MksRza) R;
RRRRRCRRMH8RV
;
RRRRRRRR-t-RCP0RNCDkRsVFRMoCCDsNR#ONCR
RRRRRRVRHRp5R3tvqR)=R3tvqR8NMRqp3)=tRRq)3)2tRRC0EMR
RRRRRRRRRRRRRRCRs0MksRza) R;
RRRRRCRRMH8RV
;
RRRRRRRRskC0swMRq p1;R
RRMRC8=R""
;

RRRRMVkOF0HM/R"=5"RRRp:HBMRmpvu uX_m)pq;)RR:MRHRvBmuXp _pumq2)RR0sCkRsMApmm 
qhRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR
H#RRRRRRRR-7-RCs#OHHb0F
M:RRRRRRRR-R-RRRRRRCR1CkRVMHO0F8MRCNODsHN0FHMRM RQ 1 R048Rj3(n.g-4gRn
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRNRR2CR)0Mks#qRwpR1 FCMRsssF
RRRRoLCHRM
RRRRR-RR-ERBCRO	PHND8$H0RRFVHkMb0sRNoCklM
0#RRRRRRRRH5VRRqp3)=tRRq-vau]_QRR20MEC
RRRRRRRRRRRRRRRR#N#CRs0w1qp R
RRRRRRRRRRRRRRRRRRRRRRRRRRCRsb0FsR3"pqR)t=vR-q_a]uHQRM=R/5)p,2R"
RRRRRRRRRRRRRRRRRRRRRRRRR#RRCsPCHR0$ m)))R;
RRRRRRRRRRRRRsRRCs0kMqRwp;1 
RRRRRRRR8CMR;HV
R
RRRRRRVRHR)5R3tq)R-=Rv]qa_RuQ2ER0CRM
RRRRRRRRRRRRRNRR#s#C0qRwp
1 RRRRRRRRRRRRRRRRRRRRRRRRRRRRsFCbs"0R))3qtRR=-avq]Q_uRRHM/p=5,")2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRP#CC0sH$)R );m)
RRRRRRRRRRRRRRRR0sCkRsMw1qp R;
RRRRRCRRMH8RV
;
RRRRRRRR-t-RC#0RbHCONPDRNCDk#R
RRRRRRVRHRp5R3tvqRj=R3NjRM)8R3tvqRj=R32jRRC0EMR
RRRRRRRRRRRRRRCRs0MksRpwq1
 ;RRRRRRRRCRM8H
V;
RRRRRRRRR--tRC0PkNDCFRVsCRoMNCsDNRO#RC
RRRRRHRRVRR5pq3vtRR=)q3vtMRN83RpqR)t=3R)qR)t2ER0CRM
RRRRRRRRRRRRRsRRCs0kMqRwp;1 
RRRRRRRR8CMR;HV
R
RRRRRRCRs0MksRza) R;
RCRRM"8R/;="
R
RR-R-
RRRRR--mC0EskRwMHO0FRM#1s0N0CR]sRC
R-RR-R

RVRRk0MOHRFMt_ auh)QBqQupq_ep5z XH:RM R)q2pRR0sCkRsMuh)QBqQupq_epRz HR#
RRRRR-RR-CR7#HOsbF0HMR:
RRRRR-RR-RRRRRRRRC1CRMVkOF0HMCR8OsDNNF0HMMRHR Q  0R18jR4(.n3-g4gnR
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRRFRhMRC
RRRRRPRRNNsHLRDCau v: R)q
p;RRRRLHCoMR
RRRRRR-R-RCBEOH	RVDRNs8CN$RRNbMsHONHbDNRPD
kCRRRRRRRRH5VRR>XRRq-vau]_QMRN8RRX<v=Rq_a]u2QRRC0EMR
RRRRRRRRRRRRRRCRs0MksRQu)huBQqep_q pz'25X;R
RRRRRRMRC8VRH;R

RRRRR-RR-CRt0sRbHHMObRNDPkNDCR
RRRRRR Rav:uR=;RX
RRRRRRRRHIED5CRRva u=R<Rq-vau]_QRR2DbFF
RRRRRRRRRRRRRRRRva u=R:Rva uRR+v]qa_u._QR;
RRRRRCRRMD8RF;Fb
RRRRRRRRHIED5CRau vRv>Rq_a]u2QRRFDFbR
RRRRRRRRRRRRRR Rav:uR= Rav-uRRavq]__.u
Q;RRRRRRRRCRM8DbFF;R

RRRRRsRRCs0kM)RuQQhBu_qpezqp a'5 2vu;R
RRMRC8 Rta)_uQQhBu_qpezqp 
;
RRRRVOkM0MHFRuBvpXX5:MRHRq) pR;RYH:RM R)q:pR=3RjjRR2skC0sBMRmpvu HXR#R
RRRRRR-R-R#7CObsH0MHF:R
RRRRRR-R-RRRRRRRR1RCCVOkM0MHFRO8CDNNs0MHFRRHMQ   R810R(4jn-3.4ngg
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRRMhFCR
RRCRLo
HMRRRRRRRRskC0sBMRmpvu 5X'XY,R2R;
RCRRMB8RvXup;R

RVRRk0MOHRFMuqmp)m_a_vBmuXp 5RZ:HBMRmpvu uX_m)pqRs2RCs0kMmRBv upX#RH
RRRRRRRRR--7OC#s0HbH:FM
RRRRRRRRR--RRRRR1RRCVCRk0MOHRFM8DCON0sNHRFMHQMR R  1R084nj(34.-g
gnRRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRN)2RCs0kMv#Rq_a]B)Z mMRFRsCsFRs
RLRRCMoH
RRRRRRRRR--BOEC	NRPDHH80F$RVMRHbRk0Nksol0CM#R
RRRRRRVRHRZ5R3tq)R-=Rv]qa_RuQ2ER0CRM
RRRRRRRRRRRRRNRR#s#C0qRwp
1 RRRRRRRRRRRRRRRRRRRRRsRRCsbF0ZR"3tq)R-=Rv]qa_RuQHuMRm)pq__amBumvp5 XZ
2"RRRRRRRRRRRRRRRRRRRRR#RRCsPCHR0$ m)))R;
RRRRRRRRRRRRRsRRCs0kMqRvaB]_Zm );R
RRRRRRMRC8VRH;R

RRRRR-RR-CRt0NRPDRkCVRFsoCCMsRNDOCN#
RRRRRRRR0sCkRsMBumvp' X53RZv*qtB5m1Z)3qtR2,Zq3vtQ*1h35Zq2)tR
2;RRRRCRM8uqmp)m_a_vBmuXp ;



RRRRMVkOF0HMmRBv upXm_a_pumqZ)5:MRHRvBmuXp Rs2RCs0kMmRBv upXm_upRq)HR#
RRRRR-RR-CR7#HOsbF0HMR:
RRRRR-RR-RRRRRRRRC1CRMVkOF0HMCR8OsDNNF0HMMRHR Q  0R18jR4(.n3-g4gnR
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRRFRhMRC
RRRRRPRRNNsHLRDCau v: R)q
p;RRRRLHCoMR
RRRRRR-R-R0tCRDPNkVCRF#sRbHCONODRN##C
RRRRRRRRRHV53RZ)= RRjj3R02RE
CMRRRRRRRRRRRRH5VRRQZ3vRR=jR3j2ER0CRM
RRRRRRRRRRRRRsRRCs0kMmRBv upXm_up'q)5jj3,3Rjj
2;RRRRRRRRRRRRCHD#VRR5Zv3QRj>R32jRRC0EMR
RRRRRRRRRRRRRRCRs0MksRvBmuXp _pumq5)'Zv3Q,qRvau]_Qe_m .)_2R;
RRRRRRRRRCRRD
#CRRRRRRRRRRRRRRRRskC0sBMRmpvu uX_m)pq'Z5-3,QvRq-vau]_Qe_m .)_2R;
RRRRRRRRRCRRMH8RVR;
RRRRRCRRMH8RV
;
RRRRRRRRH5VRRQZ3vRR=jR3j2ER0CRM
RRRRRRRRRHRRVRR5Z 3)Rj=R32jRRC0EMR
RRRRRRRRRRRRRRCRs0MksRvBmuXp _pumq5)'j,3jRjj32R;
RRRRRRRRRCRRDV#HRZ5R3R) >3RjjRR20MEC
RRRRRRRRRRRRRRRR0sCkRsMBumvp_ Xuqmp)Z'53,) Rjj32R;
RRRRRRRRRCRRD
#CRRRRRRRRRRRRRRRRskC0sBMRmpvu uX_m)pq'Z5-3,) Ravq]Q_u2R;
RRRRRRRRRCRRMH8RVR;
RRRRRCRRMH8RV
;
RRRRRRRR-t-RCb0RsOHMHDbNRDPNkVCRFosRCsMCNODRN
#CRRRRRRRRau vRR:=qa)BqZh53,QvR)Z3 
2;
RRRRRRRR0sCkRsMBumvp_ Xuqmp)1'5T5)aZ 3)*)Z3 RR+Zv3Q*QZ3v
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRat _Qu)huBQqep_q pz5va u;22
RRRR8CMRvBmuXp __amuqmp)
;
RRRRVOkM0MHFRA"q1Z"5:MRHRvBmuXp Rs2RCs0kMmRu1QQae) _ RqpHR#
RRRRR-RR-CR7#HOsbF0HMR:
RRRRR-RR-RRRRRRRRC1CRMVkOF0HMCR8OsDNNF0HMMRHR Q  0R18jR4(.n3-g4gnR
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRR2RNR1qA5RZ2=TR1)Za53*) Z 3)RZ+R3*QvZv3Q2R

RLRRCMoH
RRRRRRRRR--tRC0PkNDCFRVsCRoMNCsDNRO#RC
RRRRRsRRCs0kMmRu1QQae) _ 'qp5)1Ta35Z)Z *3R) +3RZQZv*32Qv2R;
RCRRM"8Rq"A1;R

RVRRk0MOHRFM"1qA":5ZRRHMBumvp_ Xuqmp)RR2skC0suMRma1QQ_e )p qR
H#RRRRRRRR-7-RCs#OHHb0F
M:RRRRRRRR-R-RRRRRRCR1CkRVMHO0F8MRCNODsHN0FHMRM RQ 1 R048Rj3(n.g-4gRn
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRNRR2ARq125ZRZ=R3tvq
RRRRRRRRR--RRRRRLRR2CR)0Mks#3RjjMRFRsCsF
s
RRRRLHCoMR
RRRRRR-R-RCBEOP	RN8DHHR0$FHVRM0bkRoNskMlC0R#
RRRRRHRRVRR5Z)3qtRR=-avq]Q_uR02RE
CMRRRRRRRRRRRRRRRRR#RN#0CsRpwq1R 
RRRRRRRRRRRRRRRRRRRRRRRRRsRRCsbF0ZR"3tq)R-=Rv]qa_RuQHqMRAZ152R"
RRRRRRRRRRRRRRRRRRRRRRRRR#RRCsPCHR0$ m)))R;
RRRRRRRRRRRRRRRRR0sCkRsMj;3j
RRRRRRRR8CMR;HV
R
RRRRRR-R-R0tCRDPNkVCRFosRCsMCNODRN
#CRRRRRRRRskC0sZMR3tvq;R
RRMRC8qR"A;1"
R

RVRRk0MOHRFMq5)tZH:RMmRBv upXRR2skC0suMR)BQhQpuq_peqzH R#R
RRRRRR-R-R#7CObsH0MHF:R
RRRRRR-R-RRRRRRRR1RCCVOkM0MHFRO8CDNNs0MHFRRHMQ   R810R(4jn-3.4ngg
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRRRN2q5)tZ=2RRBq)a5qhZv3Q,3RZ)
 2
RRRRRRRRsPNHDNLCaRZ Rvu:mRBv upXm_up;q)
RRRRoLCHRM
RRRRR-RR-CRt0NRPDRkCVRFsoCCMsRNDOCN#
RRRRRRRR Zav:uR=mRBv upXm_a_pumqZ)52R;
RRRRRsRRCs0kMaRZ 3vuq;)t
RRRR8CMRtq);R

RVRRk0MOHRFMq5)tZH:RMmRBv upXm_upRq)2CRs0MksRQu)huBQqep_q pzR
H#RRRRRRRR-7-RCs#OHHb0F
M:RRRRRRRR-R-RRRRRRCR1CkRVMHO0F8MRCNODsHN0FHMRM RQ 1 R048Rj3(n.g-4gRn
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRNRR2)Rqt25ZRZ=R3tq)
RRRRRRRRR--RRRRRLRR2CR)0Mks#3RjjMRFRsCsF
s
RRRRLHCoMR
RRRRRR-R-RCBEOP	RN8DHHR0$FHVRM0bkRoNskMlC0R#
RRRRRHRRVRR5Z)3qtRR=-avq]Q_uR02RE
CMRRRRRRRRRRRRRRRRR#RN#0CsRpwq1R 
RRRRRRRRRRRRRRRRRRRRRRRRRsRRCsbF0ZR"3tq)R-=Rv]qa_RuQHqMR)Zt52R"
RRRRRRRRRRRRRRRRRRRRRRRRR#RRCsPCHR0$ m)))R;
RRRRRRRRRRRRRRRRR0sCkRsMj;3j
RRRRRRRR8CMR;HV
R
RRRRRR-R-R0tCRDPNkVCRFosRCsMCNODRN
#CRRRRRRRRskC0sZMR3tq);R
RRMRC8)Rqt
;
RRRRVOkM0MHFR""-R:5ZRRHMBumvpR X2CRs0MksRvBmuXp R
H#RRRRRRRR-7-RCs#OHHb0F
M:RRRRRRRR-R-RRRRRRCR1CkRVMHO0F8MRCNODsHN0FHMRM RQ 1 R048Rj3(n.g-4gRn
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRNRR2CR)0Mks#GR-R$-[RsVFR=ZRR+GRR
[$RRRRLHCoMR
RRRRRR-R-R0tCRDPNkVCRFosRCsMCNODRN
#CRRRRRRRRskC0sBMRmpvu 5X'-)Z3 -,RZv3Q2R;
RCRRM"8R-
";
RRRRMVkOF0HM-R""ZR5:MRHRvBmuXp _pumq2)RR0sCkRsMBumvp_ Xuqmp)#RH
RRRRRRRRR--7OC#s0HbH:FM
RRRRRRRRR--RRRRR1RRCVCRk0MOHRFM8DCON0sNHRFMHQMR R  1R084nj(34.-g
gnRRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRN)2RCs0kM5#RZq3vtZ,R3tq)Rv+Rq_a]u
Q2RRRRRRRR-R-RRRRRR2RLR0)Ck#sMRFZRMsRCs
FsRRRRRRRRPHNsNCLDRva u):R ;qp
RRRRoLCHRM
RRRRR-RR-ERBCRO	PHND8$H0RRFVHkMb0sRNoCklM
0#RRRRRRRRH5VRRqZ3)=tRRq-vau]_QRR20MEC
RRRRRRRRRRRRRRRRNRR#s#C0qRwp
1 RRRRRRRRRRRRRRRRRRRRRRRRRRRRsFCbs"0RZ)3qtRR=-avq]Q_uRRHM-25Z"R
RRRRRRRRRRRRRRRRRRRRRRRRRRCR#PHCs0 $R)))m;R
RRRRRRRRRRRRRRRRRskC0sZMR;R
RRRRRRMRC8VRH;R

RRRRR-RR-CRt0sRbHHMObRNDPkNDCFRVsCRoMNCsDNRO#RC
RRRRRaRR Rvu:)=R 'qp5qZ3)Rt2+qRvau]_Q
;
RRRRRRRRskC0sBMRmpvu uX_m)pq'35Zv,qtRat _Qu)huBQqep_q pz5va u;22
RRRR8CMR""-;R

RVRRk0MOHRFMBKmhR:5ZRRHMBumvp2 XR0sCkRsMBumvpR XHR#
RRRRR-RR-CR7#HOsbF0HMR:
RRRRR-RR-RRRRRRRRC1CRMVkOF0HMCR8OsDNNF0HMMRHR Q  0R18jR4(.n3-g4gnR
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRR2RNR0)Ck#sMR-GRRR[$VRFsZRR=GRR+[R$
RLRRCMoH
RRRRRRRRR--tRC0PkNDCFRVsCRoMNCsDNRO#RC
RRRRRsRRCs0kMmRBv upXZ'53,) R3-ZQ;v2
RRRR8CMRhBmK
;
RRRRVOkM0MHFRhBmKZR5:MRHRvBmuXp _pumqR)2skC0sBMRmpvu uX_m)pqR
H#RRRRRRRR-7-RCs#OHHb0F
M:RRRRRRRR-R-RRRRRRCR1CkRVMHO0F8MRCNODsHN0FHMRM RQ 1 R048Rj3(n.g-4gRn
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRNRR2CR)0Mks#mRBv upXFROMo[kNR0C5vZ3qRt,-qZ3)
t2RRRRRRRR-R-RRRRRR2RLR0)Ck#sMRFZRMsRCs
FsRRRRRRRR-R-
RRRRRPRRNNsHLRDCau v:)RuQQhBu_qpezqp R;
RLRRCMoH
RRRRRRRRR--BOEC	NRPDHH80F$RVMRHbRk0Nksol0CM#R
RRRRRRVRHRZ5R3tq)R-=Rv]qa_RuQ2ER0CRM
RRRRRRRRRRRRRRRRR#N#CRs0w1qp R
RRRRRRRRRRRRRRRRRRRRRRRRRRCRsb0FsR3"ZqR)t=vR-q_a]uHQRMmRBhZK52R"
RRRRRRRRRRRRRRRRRRRRRRRRR#RRCsPCHR0$ m)))R;
RRRRRRRRRRRRRRRRR0sCkRsMZR;
RRRRRCRRMH8RV
;
RRRRRRRR-t-RCb0RsOHMHDbNRDPNkVCRFosRCsMCNODRN
#CRRRRRRRRH5VRRqZ3)=tRRavq]Q_uRRFsZ)3qtRR=jR3j2ER0CRM
RRRRRRRRRRRRRaRR Rvu:Z=R3tq);R
RRRRRRDRC#RC
RRRRRRRRRRRRRaRR Rvu:-=RZ)3qtR;
RRRRRCRRMH8RV
;
RRRRRRRRR0sCkRsMBumvp_ Xuqmp)Z'53tvq, Rav;u2
RRRR8CMRhBmK
;
RRRRVOkM0MHFR)1Ta:5ZRRHMBumvpR X2CRs0MksRvBmuXp R
H#RRRRRRRR-7-RCs#OHHb0F
M:RRRRRRRR-R-RRRRRRCR1CkRVMHO0F8MRCNODsHN0FHMRM RQ 1 R048Rj3(n.g-4gRn
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRhRRF
MCRRRRRRRRPHNsNCLDR Zav:uRRvBmuXp _pumq
);RRRRRRRRPHNsNCLDRzZmaRR:Bumvp; X
RRRRRRRRsPNHDNLCvRaq:tRRq) pR;
RRRRRPRRNNsHLRDCatq)R):R ;qp
RRRRoLCHRM
RRRRR-RR-CRt0NRPDRkCVRFs#ObCHRNDOCN##R
RRRRRRVRHRZ5RRv=Rq_a]B)Z mRR20MEC
RRRRRRRRRRRRRRRR0sCkRsMv]qa_ BZ)
m;RRRRRRRRCRM8H
V;
RRRRRRRRR--tRC0PkNDCFRVsCRoMNCsDNRO#RC
RRRRRZRRau vRR:=Bumvp_ Xaum_m)pq5;Z2
RRRRRRRRqavt=R:R)1Taa5Z 3vuv2qt;R
RRRRRRqRa):tR=3Rj6a*Z 3vuq;)t
R
RRRRRRVRHRB5Rma15q2)tRj>R32jRRC0EMR
RRRRRRRRRRRRRRmRZz)a3 =R:Rqavtm*B1q5a);t2
RRRRRRRRRRRRRRRRzZmav3QRR:=atvq*h1Q5)aqt
2;RRRRRRRRRRRRRRRRskC0sZMRm;za
RRRRRRRR8CMR;HV
R
RRRRRRVRHRB5Rma15q2)tRj<R32jRRC0EMR
RRRRRRRRRRRRRRmRZz)a3 =R:Rqavtm*B1q5a)+tRRavq]Q_u2R;
RRRRRRRRRRRRRZRRm3zaQ:vR=vRaq1t*Qah5qR)t+qRvau]_Q
2;RRRRRRRRRRRRRRRRskC0sZMRm;za
RRRRRRRR8CMR;HV
R
RRRRRRVRHR15RQah5q2)tRj>R32jRRC0EMR
RRRRRRRRRRRRRRmRZz)a3 =R:Rjj3;R
RRRRRRRRRRRRRRmRZzQa3v=R:RqavtQ*1hq5a);t2
RRRRRRRRRRRRRRRR0sCkRsMZamz;R
RRRRRRMRC8VRH;R

RRRRRZRRm3za): R=3RjjR;
RRRRRZRRm3zaQ:vR=vRaq1t*Qah5qR)t+qRvau]_Q
2;RRRRRRRRskC0sZMRm;za
RRRR8CMR)1Ta
;
RRRRVOkM0MHFR)1Ta:5ZRRHMBumvp_ Xuqmp)RR2skC0sBMRmpvu uX_m)pqR
H#RRRRRRRR-7-RCs#OHHb0F
M:RRRRRRRR-R-RRRRRRCR1CkRVMHO0F8MRCNODsHN0FHMRM RQ 1 R048Rj3(n.g-4gRn
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRNRR2CR)0Mks#RRZFCMRsssF
R
RRRRRRNRPsLHNDZCRmRza:mRBv upXm_up;q)
RRRRRRRRsPNHDNLCvRaq:tRRq) pR;
RRRRRPRRNNsHLRDCatq)R):R ;qp
RRRRoLCHRM
RRRRR-RR-ERBCRO	PHND8$H0RRFVHkMb0sRNoCklM
0#RRRRRRRRH5VRRqZ3)=tRRq-vau]_QRR20MEC
RRRRRRRRRRRRRRRRNRR#s#C0qRwp
1 RRRRRRRRRRRRRRRRRRRRRRRRRRRRsFCbs"0RZ)3qtRR=-avq]Q_uRRHM1aT)5"Z2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRP#CC0sH$)R );m)
RRRRRRRRRRRRRRRRsRRCs0kM;RZ
RRRRRRRR8CMR;HV
R
RRRRRR-R-R0tCRDPNkVCRF#sRbHCONODRN##C
RRRRRRRRRHV53RZvRqt=3RjjMRN83RZqR)t=3RjjRR20MEC
RRRRRRRRRRRRRRRR0sCkRsMZR;
RRRRRCRRMH8RV
;
RRRRRRRR-t-RCb0RsOHMHDbNRDPNkVCRFosRCsMCNODRN
#CRRRRRRRRatvqRR:=1aT)5vZ3q;t2
RRRRRRRR)aqt=R:R6j3*qZ3)
t;
RRRRRRRRzZmaq3vt=R:R1umQeaQ  _)q5p'atvq2
;
RRRRRRRRH5VRR1Bm5)aqt<2RRjj3R02RE
CMRRRRRRRRRRRRRRRRatq)RR:=atq)Rv+Rq_a]u
Q;RRRRRRRRCRM8H
V;
RRRRRRRRRHV5BR5ma15q2)tRj=R3Rj2NRM85h1Q5)aqt<2RRjj32RR20MEC
RRRRRRRRRRRRRRRR)aqt=R:R)aqtRR+v]qa_;uQ
RRRRRRRR8CMR;HV
R
RRRRRRmRZzqa3):tR= Rta)_uQQhBu_qpezqp q5a);t2
RRRRRRRR0sCkRsMZamz;R
RRMRC8TR1)
a;
RRRRMVkOF0HMXR u:5ZRRHMBumvpR X2CRs0MksRvBmuXp R
H#RRRRRRRR-7-RCs#OHHb0F
M:RRRRRRRR-R-RRRRRRCR1CkRVMHO0F8MRCNODsHN0FHMRM RQ 1 R048Rj3(n.g-4gRn
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRhRRF
MC
RRRRRRRRsPNHDNLC RavRu:)p q;R
RRCRLo
HMRRRRRRRR-t-RCP0RNCDkRsVFRC#bODHNR#ONCR#
RRRRRHRRVRR5ZRR=v]qa_ BZ)2mRRC0EMR
RRRRRRRRRRRRRRCRs0MksRavq]A_Bq_1 4R;
RRRRRCRRMH8RV
;
RRRRRRRRH5VRR)Z3 RR=jR3j2ER0CRM
RRRRRRRRRRRRRHRRVRR5Zv3QRv=Rq_a]uFQRs3RZQ=vRRq-vau]_QRR20MEC
RRRRRRRRRRRRRRRRRRRRRRRR0sCkRsMBumvp' X53-4jj,R3;j2
RRRRRRRRRRRRRRRR8CMR;HV
R
RRRRRRRRRRRRRRVRHRZ5R3RQv=qRvau]_Qe_m .)_R02RE
CMRRRRRRRRRRRRRRRRRRRRRRRRskC0svMRq_a]B1Aq ;_K
RRRRRRRRRRRRRRRR8CMR;HV
R
RRRRRRRRRRRRRRVRHRZ5R3RQv=vR-q_a]umQ_e_ ).RR20MEC
RRRRRRRRRRRRRRRRRRRRRRRR0sCkRsMBumvp' X5jj3,4R-3;j2
RRRRRRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMR;HV
R
RRRRRR-R-R0tCRDPNkVCRFosRCsMCNODRN
#CRRRRRRRRau vRR:= 5XuZ 3)2R;
RRRRRsRRCs0kMmRBv upXa'5 *vuB5m1Zv3Q2a,R *vu15QhZv3Q2
2;RRRRCRM8 ;Xu
R
RRkRVMHO0F MRXZu5:MRHRvBmuXp _pumq2)RR0sCkRsMBumvp_ Xuqmp)#RH
RRRRRRRRR--7OC#s0HbH:FM
RRRRRRRRR--RRRRR1RRCVCRk0MOHRFM8DCON0sNHRFMHQMR R  1R084nj(34.-g
gnRRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRN)2RCs0kMZ#RRRFMCFsssR

RRRRRPRRNNsHLRDCZva uRR:Bumvp; X
RRRRRRRRsPNHDNLCCR0lRb:)p q;R
RRRRRRNRPsLHNDZCRmRza:mRBv upXm_up;q)
RRRRoLCHRM
RRRRR-RR-ERBCRO	PHND8$H0RRFVHkMb0sRNoCklM
0#RRRRRRRRH5VRRqZ3)=tRRq-vau]_QRR20MEC
RRRRRRRRRRRRRRRRNRR#s#C0qRwp
1 RRRRRRRRRRRRRRRRRRRRRRRRRRRRsFCbs"0RZ)3qtRR=-avq]Q_uRRHM 5XuZ
2"RRRRRRRRRRRRRRRRRRRRRRRRRRRR#CCPs$H0R) )m
);RRRRRRRRRRRRRRRRRCRs0MksR
Z;RRRRRRRRCRM8H
V;
RRRRRRRRR--tRC0PkNDCFRVsbR#CNOHDNRO#
C#RRRRRRRRH5VRRvZ3q=tRRjj3R8NMRqZ3)=tRRjj3R02RE
CMRRRRRRRRRRRRRRRRskC0sBMRmpvu uX_m)pq'354jj,R3;j2
RRRRRRRR8CMR;HV
R
RRRRRRVRHRZ5R3tvqRv=Rq_a]uNQRM58RZ)3qtRR=v]qa__uQm)e _F.RsR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRZRR3tq)R-=Rv]qa__uQm)e _2.R2ER0CRM
RRRRRRRRRRRRRsRRCs0kMmRBv upXm_up'q)5j43,qRvau]_Q
2;RRRRRRRRCRM8H
V;
RRRRRRRRRHV53RZvRqt=qRvau]_Qe_m .)_R02RE
CMRRRRRRRRRRRRRRRRH5VRRqZ3)=tRRavq]Q_u_ me)R_.2ER0CRM
RRRRRRRRRRRRRRRRRRRRRsRRCs0kMmRBv upXm_up'q)5j43,qRvau]_Qe_m .)_2R;
RRRRRRRRRRRRRCRRMH8RV
;
RRRRRRRRRRRRRRRRH5VRRqZ3)=tRRq-vau]_Qe_m .)_R02RE
CMRRRRRRRRRRRRRRRRRRRRRRRRskC0sBMRmpvu uX_m)pq'354j-,Rv]qa__uQm)e _;.2
RRRRRRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMR;HV
R
RRRRRR-R-R0tCRHbsMbOHNPDRNCDkRsVFRMoCCDsNR#ONCR
RRRRRRaRZ Rvu:u=Rm)pq__amBumvp5 XZ
2;RRRRRRRRZamz3tvqRR:=uQm1a Qe_q) p '5XZu5au v32) 2R;
RRRRRZRRm3zaqR)t:t=R ua_)BQhQpuq_peqzZ 5au v32Qv;R

RRRRRsRRCs0kMmRZz
a;RRRRCRM8 ;Xu
R
RRkRVMHO0FpMRmZt5:MRHRvBmuXp Rs2RCs0kMmRBv upX#RH
RRRRRRRRR--7OC#s0HbH:FM
RRRRRRRRR--RRRRR1RRCVCRk0MOHRFM8DCON0sNHRFMHQMR R  1R084nj(34.-g
gnRRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRN)2RCs0kMB#Rmpvu 5X')p q'Wpm,3RjjF2RMsRCs
Fs
RRRRRRRRsPNHDNLCaRZ Rvu:mRBv upXm_up;q)
RRRRRRRRsPNHDNLC Rav:uRRq) pR;
RLRRCMoH
RRRRRRRRR--BOEC	NRPDHH80F$RVMRHbRk0Nksol0CM#R
RRRRRRVRHRZ5R3R) =3RjjNRRMZ8R3RQv=3RjjRR20MEC
RRRRRRRRRRRRRRRR#N#CRs0w1qp R
RRRRRRRRRRRRRRRRRRRRRRCRsb0FsR3"Z)= RRjj3R8NMRQZ3vRR=jR3jHpMRmZt52R"
RRRRRRRRRRRRRRRRRRRRR#RRCsPCHR0$ m)))R;
RRRRRRRRRRRRRsRRCs0kMmRBv upX)'5 'qpp,mWRjj32R;
RRRRRCRRMH8RV
;
RRRRRRRR-t-RCP0RNCDkRsVFRC#bODHNR#ONCR#
RRRRRHRRVRR5Zv3QRj=R32jRRC0EMR
RRRRRRRRRRRRRRVRHRZ5R3R) =4R-32jRRC0EMR
RRRRRRRRRRRRRRRRRRRRRRCRs0MksRvBmuXp '35jjv,Rq_a]u;Q2
RRRRRRRRRRRRRRRR8CMR;HV
RRRRRRRRRRRRRRRRRHV53RZ)= RRavq]R_ 2ER0CRM
RRRRRRRRRRRRRRRRRRRRRsRRCs0kMqRvaB]_A q1_
4;RRRRRRRRRRRRRRRRCRM8H
V;RRRRRRRRRRRRRRRRH5VRR)Z3 RR=4R3j2ER0CRM
RRRRRRRRRRRRRRRRRRRRRsRRCs0kMqRvaB]_Zm );R
RRRRRRRRRRRRRRMRC8VRH;R
RRRRRRMRC8VRH;R

RRRRRHRRVRR5Z 3)Rj=R32jRRC0EMR
RRRRRRRRRRRRRRVRHR35ZQ=vRRj432ER0CRM
RRRRRRRRRRRRRRRRRRRRRsRRCs0kMmRBv upXj'53Rj,v]qa__uQm)e _;.2
RRRRRRRRRRRRRRRR8CMR;HV
RRRRRRRRRRRRRRRRRHV5QZ3vRR=-j432ER0CRM
RRRRRRRRRRRRRRRRRRRRRsRRCs0kMmRBv upXj'53Rj,-avq]Q_u_ me)2_.;R
RRRRRRRRRRRRRRMRC8VRH;R
RRRRRRMRC8VRH;R

RRRRR-RR-CRt0NRPDRkCVRFsoCCMsRNDOCN#
RRRRRRRR Zav:uR=mRBv upXm_a_pumqZ)52R;
RRRRRaRR Rvu:p=RmZt5au v3tvq2R;
RRRRRsRRCs0kMmRBv upXa'5 ,vuR Zavqu3);t2
RRRR8CMRtpm;R

RVRRk0MOHRFMp.mt5RZ:HBMRmpvu 2XRR0sCkRsMBumvpR XHR#
RRRRR-RR-CR7#HOsbF0HMR:
RRRRR-RR-RRRRRRRRC1CRMVkOF0HMCR8OsDNNF0HMMRHR Q  0R18jR4(.n3-g4gnR
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRR2RNR0)Ck#sMRvBmuXp ' 5)qpp'mRW,j23jRRFMCFsssR

RRRRRPRRNNsHLRDCZva uRR:Bumvp_ Xuqmp)R;
RRRRRPRRNNsHLRDCau vR):R ;qp
RRRRoLCH
M
RRRRRRRR-B-RE	CORDPNH08H$VRFRbHMkN0RslokC#M0
RRRRRRRRRHV53RZ)= RRjj3RMRN83RZQ=vRRjj3R02RE
CMRRRRRRRRRRRRRRRRNC##sw0Rq p1
RRRRRRRRRRRRRRRRRRRRRRRRbsCFRs0")Z3 RR=jR3jNRM8Zv3QRj=R3HjRMmRptZ.52R"
RRRRRRRRRRRRRRRRRRRRR#RRCsPCHR0$ m)))R;
RRRRRRRRRRRRRsRRCs0kMmRBv upX)'5 'qpp,mWRjj32R;
RRRRRCRRMH8RV
;
RRRRRRRR-t-RCP0RNCDkRsVFRC#bODHNR#ONCR#
RRRRRHRRVRR5Zv3QRj=R32jRRC0EMR
RRRRRRRRRRRRRRVRHRZ5R3R) =3R.jRR20MEC
RRRRRRRRRRRRRRRRRRRRRRRR0sCkRsMv]qa_qBA14 _;R
RRRRRRRRRRRRRRMRC8VRH;R
RRRRRRRRRRRRRRVRHRZ5R3R) =3R4jRR20MEC
RRRRRRRRRRRRRRRRRRRRRRRR0sCkRsMv]qa_ BZ)
m;RRRRRRRRRRRRRRRRCRM8H
V;RRRRRRRRCRM8H
V;
RRRRRRRRR--tRC0PkNDCFRVsCRoMNCsDNRO#RC
RRRRRZRRau vRR:=Bumvp_ Xaum_m)pq5;Z2
RRRRRRRRva u=R:Ravq]m_ptm._w*_ p5mtZva uq3vt
2;RRRRRRRRskC0sBMRmpvu 5X'au v,qRvap]_m_t.m w_* Zavqu3);t2
RRRR8CMRtpm.
;
RRRRVOkM0MHFRtpm4Zj5:MRHRvBmuXp Rs2RCs0kMmRBv upX#RH
RRRRRRRRR--7OC#s0HbH:FM
RRRRRRRRR--RRRRR1RRCVCRk0MOHRFM8DCON0sNHRFMHQMR R  1R084nj(34.-g
gnRRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRN)2RCs0kMB#Rmpvu 5X')p q'Wpm,3RjjF2RMsRCs
Fs
RRRRRRRRsPNHDNLCaRZ Rvu:mRBv upXm_up;q)
RRRRRRRRsPNHDNLC Rav:uRRq) pR;
RLRRCMoH
RRRRRRRRR--BOEC	NRPDHH80F$RVMRHbRk0Nksol0CM#R
RRRRRRVRHRZ5R3R) =3RjjNRRMZ8R3RQv=3RjjRR20MEC
RRRRRRRRRRRRRRRR#N#CRs0w1qp R
RRRRRRRRRRRRRRRRRRRRRRCRsb0FsR3"Z)= RRjj3R8NMRQZ3vRR=jR3jHpMRmjt45"Z2
RRRRRRRRRRRRRRRRRRRRRRRRP#CC0sH$)R );m)
RRRRRRRRRRRRRRRR0sCkRsMBumvp' X5q) pm'pWj,R3;j2
RRRRRRRR8CMR;HV
R
RRRRRR-R-R0tCRDPNkVCRF#sRbHCONODRN##C
RRRRRRRRRHV53RZQ=vRRjj3R02RE
CMRRRRRRRRRRRRRRRRH5VRR)Z3 RR=4jj3R02RE
CMRRRRRRRRRRRRRRRRRRRRRRRRskC0svMRq_a]B1Aq ;_4
RRRRRRRRRRRRRRRR8CMR;HV
RRRRRRRRRRRRRRRRRHV53RZ)= RRj43R02RE
CMRRRRRRRRRRRRRRRRRRRRRRRRskC0svMRq_a]B)Z mR;
RRRRRRRRRRRRRCRRMH8RVR;
RRRRRCRRMH8RV
;
RRRRRRRR-t-RCP0RNCDkRsVFRMoCCDsNR#ONCR
RRRRRRaRZ Rvu:B=Rmpvu aX_mm_up5q)Z
2;RRRRRRRRau vRR:=v]qa_tpm4mj_w*_ p5mtZva uq3vt
2;RRRRRRRRskC0sBMRmpvu 5X'au v,qRvap]_mjt4__mw a*Z 3vuq2)t;R
RRMRC8mRpt;4j
R

RVRRk0MOHRFMp5mtZH:RMmRBv upXm_upRq)2CRs0MksRvBmuXp _pumqH)R#R
RRRRRR-R-R#7CObsH0MHF:R
RRRRRR-R-RRRRRRRR1RCCVOkM0MHFRO8CDNNs0MHFRRHMQ   R810R(4jn-3.4ngg
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRRRN2)kC0sRM#Bumvp_ Xuqmp) 5)q]p'Q,t]Ravq]Q_u2MRFRsCsF
s
RRRRRRRRPHNsNCLDR Zav:uRRvBmuXp ;R
RRRRRRNRPsLHNDZCRmRza:mRBv upXm_up;q)
RRRRoLCHRM
RRRRR-RR-ERBCRO	PHND8$H0RRFVHkMb0sRNoCklM
0#RRRRRRRRH5VRRvZ3q<tR=3RjjRR20MEC
RRRRRRRRRRRRRRRR#N#CRs0w1qp R
RRRRRRRRRRRRRRRRRRRRRRCRsb0FsR3"ZvRqt<j=R3HjRMmRpt25Z"R
RRRRRRRRRRRRRRRRRRRRRRCR#PHCs0 $R)))m;R
RRRRRRRRRRRRRRCRs0MksRvBmuXp _pumq5)')p q't]Q]v,Rq_a]u;Q2
RRRRRRRR8CMR;HV
R
RRRRRRVRHRZ5R3tq)R-=Rv]qa_RuQ2ER0CRM
RRRRRRRRRRRRRRRRR#N#CRs0w1qp R
RRRRRRRRRRRRRRRRRRRRRRRRRRCRsb0FsR3"ZqR)t=vR-q_a]uHQRMmRpt25Z"R
RRRRRRRRRRRRRRRRRRRRRRRRRRCR#PHCs0 $R)))m;R
RRRRRRRRRRRRRRCRs0MksRvBmuXp _pumq5)')p q't]Q]v,Rq_a]u;Q2
RRRRRRRR8CMR;HV
R
RRRRRR-R-RlBFbCk0RDPNkVCRF#sRbHCONODRN##C
RRRRRRRRRHV5vZ3q=tRRj43R02RE
CMRRRRRRRRRRRRRRRRH5VRRqZ3)=tRRjj3R02RE
CMRRRRRRRRRRRRRRRRRRRRRRRRskC0sBMRmpvu uX_m)pq'35jjj,R3;j2
RRRRRRRRRRRRRRRR8CMR;HV
R
RRRRRRRRRRRRRRVRHRZ5R3tq)Rv=Rq_a]u2QRRC0EMR
RRRRRRRRRRRRRRRRRRRRRRCRs0MksRvBmuXp _pumq5)'v]qa_,uQRavq]Q_u_ me)2_.;R
RRRRRRRRRRRRRRMRC8VRH;R

RRRRRRRRRRRRRHRRVRR5Z)3qtRR=v]qa__uQm)e _2.RRC0EMR
RRRRRRRRRRRRRRRRRRRRRRCRs0MksRvBmuXp _pumq5)'v]qa__uQm)e _R.,v]qa__uQm)e _;.2
RRRRRRRRRRRRRRRR8CMR;HV
R
RRRRRRRRRRRRRRVRHRZ5R3tq)R-=Rv]qa__uQm)e _2.RRC0EMR
RRRRRRRRRRRRRRRRRRRRRRCRs0MksRvBmuXp _pumq5)'v]qa__uQm)e _R.,-avq]Q_u_ me)2_.;R
RRRRRRRRRRRRRRMRC8VRH;R
RRRRRRMRC8VRH;R

RRRRRHRRVRR5Zq3vtRR=v]qa_N RMZ8R3tq)Rj=R32jRRC0EMR
RRRRRRRRRRRRRRCRs0MksRvBmuXp _pumq5)'4,3jRjj32R;
RRRRRCRRMH8RV
;
RRRRRRRR-B-RFklb0PCRNCDkRsVFRMoCCDsNR#ONCR
RRRRRRaRZ 3vu): R=mRpt35Zv2qt;R
RRRRRRaRZ 3vuQ:vR=3RZq;)t
RRRRRRRRzZma=R:RvBmuXp __amuqmp)a5Z 2vu;R
RRRRRRCRs0MksRzZmaR;
RCRRMp8Rm
t;
R

RVRRk0MOHRFMp.mt5RZ:HBMRmpvu uX_m)pqRs2RCs0kMmRBv upXm_upRq)HR#
RRRRR-RR-CR7#HOsbF0HMR:
RRRRR-RR-RRRRRRRRC1CRMVkOF0HMCR8OsDNNF0HMMRHR Q  0R18jR4(.n3-g4gnR
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRR2RNR0)Ck#sMRvBmuXp _pumq))5 'qp]]Qt,qRvau]_QF2RMsRCs
Fs
RRRRRRRRsPNHDNLCaRZ Rvu:mRBv upXR;
RRRRRPRRNNsHLRDCZamzRB:Rmpvu uX_m)pq;R
RRCRLo
HMRRRRRRRR-B-RE	CORDPNH08H$VRFRbHMkN0RslokC#M0
RRRRRRRRRHV53RZvRqt<j=R32jRRC0EMR
RRRRRRRRRRRRRR#RN#0CsRpwq1R 
RRRRRRRRRRRRRRRRRRRRRsRRCsbF0ZR"3tvqRR<=jR3jHpMRm5t.Z
2"RRRRRRRRRRRRRRRRRRRRRRRR#CCPs$H0R) )m
);RRRRRRRRRRRRRRRRskC0sBMRmpvu uX_m)pq' 5)q]p'Q,t]Ravq]Q_u2R;
RRRRRCRRMH8RV
;
RRRRRRRRH5VRRqZ3)=tRRq-vau]_QRR20MEC
RRRRRRRRRRRRRRRRNRR#s#C0qRwp
1 RRRRRRRRRRRRRRRRRRRRRRRRRRRRsFCbs"0RZ)3qtRR=-avq]Q_uRRHMp.mt5"Z2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRP#CC0sH$)R );m)
RRRRRRRRRRRRRRRR0sCkRsMBumvp_ Xuqmp))'5 'qp]]Qt,qRvau]_Q
2;RRRRRRRRCRM8H
V;
RRRRRRRRR--BbFlkR0CPkNDCFRVsbR#CNOHDNRO#
C#RRRRRRRRH5VRZq3vtRR=4R3jNRM8Z)3qtRR=jR3j2ER0CRM
RRRRRRRRRRRRRsRRCs0kMmRBv upXm_up'q)5jj3,3Rjj
2;RRRRRRRRCRM8H
V;
RRRRRRRRRHV53RZvRqt=3R.jMRN83RZqR)t=3RjjRR20MEC
RRRRRRRRRRRRRRRR0sCkRsMBumvp_ Xuqmp)4'53Rj,j23j;R
RRRRRRMRC8VRH;R

RRRRR-RR-FRBl0bkCNRPDRkCVRFsoCCMsRNDOCN#
RRRRRRRR Zav)u3 =R:Ravq]m_ptm._w*_ p5mtZq3vt
2;RRRRRRRRZva uv3QRR:=v]qa_tpm.w_m_Z *3tq);R
RRRRRRmRZz:aR=mRBv upXm_a_pumqZ)5au v2R;
RRRRRsRRCs0kMmRZz
a;RRRRCRM8p.mt;R

RVRRk0MOHRFMp4mtj:5ZRRHMBumvp_ Xuqmp)RR2skC0sBMRmpvu uX_m)pqR
H#RRRRRRRR-7-RCs#OHHb0F
M:RRRRRRRR-R-RRRRRRCR1CkRVMHO0F8MRCNODsHN0FHMRM RQ 1 R048Rj3(n.g-4gRn
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRNRR2CR)0Mks#mRBv upXm_up5q))p q't]Q]v,Rq_a]uRQ2FCMRsssF
RRRRRRRRsPNHDNLCaRZ Rvu:mRBv upXR;
RRRRRPRRNNsHLRDCZamzRB:Rmpvu uX_m)pq;R
RRCRLo
HMRRRRRRRR-B-RE	CORDPNH08H$VRFRbHMkN0RslokC#M0
RRRRRRRRRHV53RZvRqt<j=R32jRRC0EMR
RRRRRRRRRRRRRR#RN#0CsRpwq1R 
RRRRRRRRRRRRRRRRRRRRRsRRCsbF0ZR"3tvqRR<=jR3jHpMRmjt45"Z2
RRRRRRRRRRRRRRRRRRRRRRRRP#CC0sH$)R );m)
RRRRRRRRRRRRRRRR0sCkRsMBumvp_ Xuqmp))'5 'qp]]Qt,qRvau]_Q
2;RRRRRRRRCRM8H
V;
R
RRRRRRVRHRZ5R3tq)R-=Rv]qa_RuQ2ER0CRM
RRRRRRRRRRRRRRRRR#N#CRs0w1qp R
RRRRRRRRRRRRRRRRRRRRRRRRRRbsCFRs0"qZ3)=tRRq-vau]_QMRHRtpm4Zj52R"
RRRRRRRRRRRRRRRRRRRRRRRRRCR#PHCs0 $R)))m;R
RRRRRRRRRRRRRRCRs0MksRvBmuXp _pumq5)')p q't]Q]v,Rq_a]u;Q2
RRRRRRRR8CMR;HV
R
RRRRRR-R-RlBFbCk0RDPNkVCRF#sRbHCONODRN##C
RRRRRRRRRHV5vZ3q=tRRj43R8NMRqZ3)=tRRjj3R02RE
CMRRRRRRRRRRRRRRRRskC0sBMRmpvu uX_m)pq'35jjj,R3;j2
RRRRRRRR8CMR;HV
R
RRRRRRVRHRZ5R3tvqR4=RjR3jNRM8Z)3qtRR=jR3j2ER0CRM
RRRRRRRRRRRRRsRRCs0kMmRBv upXm_up'q)5j43,3Rjj
2;RRRRRRRRCRM8H
V;
RRRRRRRRR--BbFlkR0CPkNDCFRVsCRoMNCsDNRO#RC
RRRRRZRRau v3R) :v=Rq_a]p4mtjw_m_p *mZt53tvq2R;
RRRRRZRRau v3RQv:v=Rq_a]p4mtjw_m_Z *3tq);R
RRRRRRmRZz:aR=mRBv upXm_a_pumqZ)5au v2R;
RRRRRsRRCs0kMmRZz
a;RRRRCRM8p4mtj
;
RRRRVOkM0MHFRtpm5RZ:HBMRmpvu RX;A q1:MRHRq) pRR2skC0sBMRmpvu HXR#R
RRRRRR-R-R#7CObsH0MHF:R
RRRRRR-R-RRRRRRRR1RCCVOkM0MHFRO8CDNNs0MHFRRHMQ   R810R(4jn-3.4ngg
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRRRN2)kC0sRM#Bumvp' X5q) pm'pWj,R3Rj2FCMRsssF
R
RRRRRRNRPsLHNDZCRau vRB:Rmpvu uX_m)pq;R
RRRRRRNRPsLHNDaCR )vu RR:)p q;R
RRRRRRNRPsLHNDaCR QvuvRR:)p q;R
RRCRLo
HMRRRRRRRR-B-RE	CORDPNH08H$VRFRbHMkN0RslokC#M0
RRRRRRRRRHV53RZ)= RRjj3RMRN83RZQ=vRRjj3R02RE
CMRRRRRRRRRRRRRRRRNC##sw0Rq p1
RRRRRRRRRRRRRRRRRRRRRRRRbsCFRs0")Z3 RR=jR3jNRM8Zv3QRj=R3HjRMmRpt,5ZA q12R"
RRRRRRRRRRRRRRRRRRRRR#RRCsPCHR0$ m)))R;
RRRRRRRRRRRRRsRRCs0kMmRBv upX)'5 'qpp,mWRjj32R;
RRRRRCRRMH8RV
;
RRRRRRRRH5VRR1Aq =R<Rjj3RRFsA q1R4=R32jRRC0EMR
RRRRRRRRRRRRRR#RN#0CsRpwq1R 
RRRRRRRRRRRRRRRRRRRRRsRRCsbF0AR"qR1 <j=R3FjRsqRA1= RRj43RRHMp5mtZq,A1" 2
RRRRRRRRRRRRRRRRRRRRRRRRP#CC0sH$)R );m)
RRRRRRRRRRRRRRRR0sCkRsMBumvp' X5q) pm'pWj,R3;j2
RRRRRRRR8CMR;HV
R
RRRRRR-R-R0tCRDPNkVCRF#sRbHCONODRN##C
RRRRRRRRRHV53RZQ=vRRjj3R02RE
CMRRRRRRRRRRRRRRRRH5VRR)Z3 RR=A q1R02RE
CMRRRRRRRRRRRRRRRRRRRRRRRRskC0svMRq_a]B1Aq ;_4
RRRRRRRRRRRRRRRR8CMR;HV
RRRRRRRRRRRRRRRRRHV53RZ)= RRj43R02RE
CMRRRRRRRRRRRRRRRRRRRRRRRRskC0svMRq_a]B)Z mR;
RRRRRRRRRRRRRCRRMH8RVR;
RRRRRCRRMH8RV
;
RRRRRRRR-t-RCP0RNCDkRsVFRMoCCDsNR#ONCR
RRRRRRaRZ Rvu:B=Rmpvu aX_mm_up5q)Z
2;RRRRRRRRau v): R=mRpta5Z 3vuv,qtR1Aq 
2;RRRRRRRRau vQ:vR=aRZ 3vuq/)tp5mtA q12R;
RRRRRsRRCs0kMmRBv upXa'5 )vu a,R Qvuv
2;RRRRCRM8p;mt
R
RRkRVMHO0FpMRmZt5:MRHRvBmuXp _pumqR);A q1:MRHRq) pRR2skC0sBMRmpvu uX_m)pqR
H#RRRRRRRR-7-RCs#OHHb0F
M:RRRRRRRR-R-RRRRRRCR1CkRVMHO0F8MRCNODsHN0FHMRM RQ 1 R048Rj3(n.g-4gRn
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRNRR2CR)0Mks#mRBv upXm_up5q))p q't]Q]v,Rq_a]uRQ2FCMRsssF
R
RRRRRRNRPsLHNDZCRau vRB:Rmpvu 
X;RRRRRRRRPHNsNCLDRzZmaRR:Bumvp_ Xuqmp)R;
RLRRCMoH
RRRRRRRRR--BOEC	NRPDHH80F$RVMRHbRk0Nksol0CM#R
RRRRRRVRHRZ5R3tvqRR<=jR3j2ER0CRM
RRRRRRRRRRRRRNRR#s#C0qRwp
1 RRRRRRRRRRRRRRRRRRRRRRRRsFCbs"0RZq3vt=R<Rjj3RRHMp5mtZq,A1" 2
RRRRRRRRRRRRRRRRRRRRRRRRP#CC0sH$)R );m)
RRRRRRRRRRRRRRRR0sCkRsMBumvp_ Xuqmp))'5 'qp]]Qt,qRvau]_Q
2;RRRRRRRRCRM8H
V;
RRRRRRRRRHV5qRA1< R=3RjjsRFR1Aq RR=4R3j2ER0CRM
RRRRRRRRRRRRRNRR#s#C0qRwp
1 RRRRRRRRRRRRRRRRRRRRRRRRsFCbs"0RA q1RR<=jR3jFAsRqR1 =3R4jMRHRtpm5AZ,q21 "R
RRRRRRRRRRRRRRRRRRRRRRCR#PHCs0 $R)))m;R
RRRRRRRRRRRRRRCRs0MksRvBmuXp _pumq5)')p q't]Q]v,Rq_a]u;Q2
RRRRRRRR8CMR;HV
R
RRRRRRVRHRZ5R3tq)R-=Rv]qa_RuQ2ER0CRM
RRRRRRRRRRRRRNRR#s#C0qRwp
1 RRRRRRRRRRRRRRRRRRRRRRRRRsRRCsbF0ZR"3tq)R-=Rv]qa_RuQHpMRmZt5,1Aq 
2"RRRRRRRRRRRRRRRRRRRRRRRRR#RRCsPCHR0$ m)))R;
RRRRRRRRRRRRRsRRCs0kMmRBv upXm_up'q)5q) pQ']tR],v]qa_2uQ;R
RRRRRRMRC8VRH;R

RRRRR-RR-FRBl0bkCNRPDRkCVRFs#ObCHRNDOCN##R
RRRRRRVRHR35ZvRqt=3R4jMRN83RZqR)t=3RjjRR20MEC
RRRRRRRRRRRRRRRR0sCkRsMBumvp_ Xuqmp)j'53Rj,j23j;R
RRRRRRMRC8VRH;R

RRRRRHRRVRR5Zq3vtRR=A q1R8NMRqZ3)=tRRjj3R02RE
CMRRRRRRRRRRRRRRRRskC0sBMRmpvu uX_m)pq'354jj,R3;j2
RRRRRRRR8CMR;HV
R
RRRRRR-R-RlBFbCk0RDPNkVCRFosRCsMCNODRN
#CRRRRRRRRZva u 3)RR:=p5mtZq3vtA,Rq21 ;R
RRRRRRaRZ 3vuQ:vR=3RZq/)tp5mtA q12R;
RRRRRZRRmRza:B=Rmpvu aX_mm_up5q)Zva u
2;RRRRRRRRskC0sZMRm;za
RRRR8CMRtpm;


RRRRVOkM0MHFRh1Q5RZ:HBMRmpvu 2XRR0sCkRsMBumvpR XHR#
RRRRR-RR-CR7#HOsbF0HMR:
RRRRR-RR-RRRRRRRRC1CRMVkOF0HMCR8OsDNNF0HMMRHR Q  0R18jR4(.n3-g4gnR
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRRFRhMRC
RLRRCMoH
RRRRRRRRR--tRC0PkNDCFRVsbR#CNOHDNRO#
C#RRRRRRRRH5VRRQZ3vRR=jR3j2ER0CRM
RRRRRRRRRRRRRHRRVRR5Z 3)Rj=R3FjRs3RZ)= RRavq]Q_u2ER0CRM
RRRRRRRRRRRRRRRRRRRRRsRRCs0kMqRvaB]_Zm );R
RRRRRRRRRRRRRRMRC8VRH;R
RRRRRRMRC8VRH;R

RRRRR-RR-CRt0NRPDRkCVRFsoCCMsRNDOCN#
RRRRRRRR0sCkRsMBumvp' X5h1Q5)Z3 B2*m51]Zv3Q2B,RmZ1532) *h1Q]35ZQ2v2;R
RRMRC8QR1h
;
RRRRVOkM0MHFRh1Q5RZ:HBMRmpvu uX_m)pqRs2RCs0kMmRBv upXm_upRq)HR#
RRRRR-RR-CR7#HOsbF0HMR:
RRRRR-RR-RRRRRRRRC1CRMVkOF0HMCR8OsDNNF0HMMRHR Q  0R18jR4(.n3-g4gnR
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRR2RNR0)Ck#sMRvBmuXp _pumqj)53Rj,j23jRRFMCFsssR

RRRRRPRRNNsHLRDCZR4,Z:.RRvBmuXp ;R
RRRRRRNRPsLHNDZCRmRza:mRBv upXm_up;q)
RRRRoLCHRM
RRRRR-RR-ERBCRO	PHND8$H0RRFVHkMb0sRNoCklM
0#RRRRRRRRH5VRRqZ3)=tRRq-vau]_QRR20MEC
RRRRRRRRRRRRRRRR#N#CRs0w1qp R
RRRRRRRRRRRRRRRRRRRRRRRRRRCRsb0FsR3"ZqR)t=vR-q_a]uHQRMQR1h25Z"R
RRRRRRRRRRRRRRRRRRRRRRRRRRCR#PHCs0 $R)))m;R
RRRRRRRRRRRRRRCRs0MksRvBmuXp _pumq5)'j,3jRjj32R;
RRRRRCRRMH8RV
;
RRRRRRRR-B-RFklb0PCRNCDkRsVFRC#bODHNR#ONCR#
RRRRRHRRVRR5Zq3vtRR=jR3jNRM8Z)3qtRR=jR3j2ER0CRM
RRRRRRRRRRRRRsRRCs0kMmRBv upXm_up'q)5jj3,3Rjj
2;RRRRRRRRCRM8H
V;
RRRRRRRRRHV53RZvRqt=qRvau]_QMRN83RZqR)t=3RjjRR20MEC
RRRRRRRRRRRRRRRR0sCkRsMBumvp_ Xuqmp)j'53Rj,j23j;R
RRRRRRMRC8VRH;R

RRRRR-RR-FRBl0bkCNRPDRkCVRFsoCCMsRNDOCN#
RRRRRRRRRZ4:u=Rm)pq__amBumvp5 XZ
2;RRRRRRRRZ:.R=mRBv upX1'5QZh54 3)2m*B1Z]54v3Q2B,RmZ154 3)2Q*1hZ]54v3Q2
2;RRRRRRRRZamzRR:=Bumvp_ Xaum_m)pq52Z.;R
RRRRRRCRs0MksRzZmaR;
RCRRM18RQ
h;
RRRRMVkOF0HMmRB1:5ZRRHMBumvpR X2CRs0MksRvBmuXp R
H#RRRRRRRR-7-RCs#OHHb0F
M:RRRRRRRR-R-RRRRRRCR1CkRVMHO0F8MRCNODsHN0FHMRM RQ 1 R048Rj3(n.g-4gRn
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRhRRF
MCRRRRLHCoM


RRRRRRRR-t-RCP0RNCDkRsVFRC#bODHNR#ONCR#
RRRRRHRRVRR5Zv3QRj=R32jRRC0EMR
RRRRRRRRRRRRRRVRHRZ5R3R) =qRvau]_Qe_m .)_RRFsZ 3)R-=Rv]qa__uQm)e _R.20MEC
RRRRRRRRRRRRRRRRRRRRRRRR0sCkRsMv]qa_ BZ)
m;RRRRRRRRRRRRRRRRCRM8H
V;RRRRRRRRCRM8H
V;
RRRRRRRRR--tRC0PkNDCFRVsCRoMNCsDNRO#RC
RRRRRsRRCs0kMmRBv upXB'5mZ1532) *1Bm]35ZQ,v2RQ-1h35Z)* 21]Qh5QZ3v;22
RRRR8CMR1Bm;R

RVRRk0MOHRFMB5m1ZH:RMmRBv upXm_upRq)2CRs0MksRvBmuXp _pumqH)R#R
RRRRRR-R-R#7CObsH0MHF:R
RRRRRR-R-RRRRRRRR1RCCVOkM0MHFRO8CDNNs0MHFRRHMQ   R810R(4jn-3.4ngg
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRRRN2)kC0sRM#Bumvp_ Xuqmp)35jjj,R3Rj2FCMRsssF
R
RRRRRRNRPsLHNDZCR4Z,R.RR:Bumvp; X
RRRRRRRRsPNHDNLCmRZz:aRRvBmuXp _pumq
);RRRRLHCoMR
RRRRRR-R-RCBEOP	RN8DHHR0$FHVRM0bkRoNskMlC0R#
RRRRRHRRVRR5Z)3qtRR=-avq]Q_uR02RE
CMRRRRRRRRRRRRRRRRNC##sw0Rq p1
RRRRRRRRRRRRRRRRRRRRRRRRRRRRbsCFRs0"qZ3)=tRRq-vau]_QMRHR1Bm5"Z2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRP#CC0sH$)R );m)
RRRRRRRRRRRRRRRR0sCkRsMBumvp_ Xuqmp)j'53Rj,j23j;R
RRRRRRMRC8VRH;R

RRRRR-RR-FRBl0bkCNRPDRkCVRFs#ObCHRNDOCN##R
RRRRRRVRHRZ5R3tvqRv=Rq_a]umQ_e_ ).MRN83RZqR)t=3RjjRR20MEC
RRRRRRRRRRRRRRRR0sCkRsMBumvp_ Xuqmp)j'53Rj,j23j;R
RRRRRRMRC8VRH;R

RRRRRHRRVRR5Zq3vtRR=v]qa__uQm)e _N.RMZ8R3tq)Rv=Rq_a]u2QRRC0EMR
RRRRRRRRRRRRRRCRs0MksRvBmuXp _pumq5)'j,3jRjj32R;
RRRRRCRRMH8RV
;
RRRRRRRR-B-RFklb0PCRNCDkRsVFRMoCCDsNR#ONCR
RRRRRR4RZRR:=uqmp)m_a_vBmuXp 5;Z2
RRRRRRRRRZ.:B=Rmpvu 5X'B5m1Z)43 B2*m51]ZQ43vR2,-h1Q53Z4)* 21]Qh53Z4Q2v2;R
RRRRRRmRZz:aR=mRBv upXm_a_pumqZ)5.
2;RRRRRRRRskC0sZMRm;za
RRRR8CMR1Bm;R

RVRRk0MOHRFM1]Qh5RZ:HBMRmpvu 2XRR0sCkRsMBumvpR XHR#
RRRRR-RR-CR7#HOsbF0HMR:
RRRRR-RR-RRRRRRRRC1CRMVkOF0HMCR8OsDNNF0HMMRHR Q  0R18jR4(.n3-g4gnR
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRRFRhMRC
RLRRCMoH
RRRRRRRRR--tRC0PkNDCFRVsbR#CNOHDNRO#
C#RRRRRRRRH5VRR)Z3 RR=jR3j2ER0CRM
RRRRRRRRRRRRRHRRVRR5Zv3QRj=R3FjRs3RZQ=vRRavq]Q_uR02RE
CMRRRRRRRRRRRRRRRRRRRRRRRRskC0svMRq_a]B)Z mR;
RRRRRRRRRRRRRCRRMH8RV
;

R
RRRRRRRRRRRRRRVRHRZ5R3RQv=qRvau]_Qe_m .)_R02RE
CMRRRRRRRRRRRRRRRRRRRRRRRRskC0svMRq_a]B1Aq ;_K
RRRRRRRRRRRRRRRR8CMR;HV
R
RRRRRRRRRRRRRRVRHRZ5R3RQv=vR-q_a]umQ_e_ ).RR20MEC
RRRRRRRRRRRRRRRRRRRRRRRR0sCkRsM-avq]A_Bq_1 KR;
RRRRRRRRRRRRRCRRMH8RVR;
RRRRRCRRMH8RV
;
RRRRRRRR-t-RCP0RNCDkRsVFRMoCCDsNR#ONCR
RRRRRRCRs0MksRvBmuXp 'Q51hZ]532) *1Bm5QZ3vR2,B]m15)Z3 12*QZh532Qv2R;
RCRRM18RQ;h]
R
RRkRVMHO0F1MRQ5h]ZH:RMmRBv upXm_upRq)2CRs0MksRvBmuXp _pumqH)R#R
RRRRRR-R-R#7CObsH0MHF:R
RRRRRR-R-RRRRRRRR1RCCVOkM0MHFRO8CDNNs0MHFRRHMQ   R810R(4jn-3.4ngg
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRRRN2)kC0sRM#Bumvp_ Xuqmp)35jjj,R3Rj2FCMRsssF
R
RRRRRRNRPsLHNDZCR4Z,R.RR:Bumvp; X
RRRRRRRRsPNHDNLCmRZz:aRRvBmuXp _pumq
);RRRRLHCoMR
RRRRRR-R-RCBEOP	RN8DHHR0$FHVRM0bkRoNskMlC0R#
RRRRRHRRVRR5Z)3qtRR=-avq]Q_uR02RE
CMRRRRRRRRRRRRRRRRNC##sw0Rq p1
RRRRRRRRRRRRRRRRRRRRRRRRRRRRbsCFRs0"qZ3)=tRRq-vau]_QMRHRh1Q]25Z"R
RRRRRRRRRRRRRRRRRRRRRRRRRRCR#PHCs0 $R)))m;R
RRRRRRRRRRRRRRCRs0MksRvBmuXp _pumq5)'j,3jRjj32R;
RRRRRCRRMH8RV
;
RRRRRRRR-B-RFklb0PCRNCDkRsVFRC#bODHNR#ONCR#
RRRRRHRRVRR5Zq3vtRR=jR3jNRM8Z)3qtRR=jR3j2ER0CRM
RRRRRRRRRRRRRsRRCs0kMmRBv upXm_up'q)5jj3,3Rjj
2;RRRRRRRRCRM8H
V;
RRRRRRRRRHV53RZvRqt=qRvau]_QMRN83RZqR)t=qRvau]_Qe_m .)_R02RE
CMRRRRRRRRRRRRRRRRskC0sBMRmpvu uX_m)pq'35jjj,R3;j2
RRRRRRRR8CMR;HV
R
RRRRRRVRHRZ5R3tvqRv=Rq_a]umQ_e_ ).MRN83RZqR)t=qRvau]_Qe_m .)_R02RE
CMRRRRRRRRRRRRRRRRskC0sBMRmpvu uX_m)pq'354jv,Rq_a]umQ_e_ ).
2;RRRRRRRRCRM8H
V;
RRRRRRRRRHV53RZvRqt=qRvau]_Qe_m .)_R8NMRqZ3)=tRRq-vau]_Qe_m .)_R02RE
CMRRRRRRRRRRRRRRRRskC0sBMRmpvu uX_m)pq'354j-,Rv]qa__uQm)e _;.2
RRRRRRRR8CMR;HV
R
RRRRRR-R-RlBFbCk0RDPNkVCRFosRCsMCNODRN
#CRRRRRRRRZ:4R=mRup_q)aBm_mpvu ZX52R;
RRRRRZRR.=R:RvBmuXp 'Q51hZ]54 3)2m*B145Z32Qv,mRB1Z]54 3)2Q*1h45Z32Qv2R;
RRRRRZRRmRza:B=Rmpvu aX_mm_up5q)Z;.2
RRRRRRRR0sCkRsMZamz;R
RRMRC8QR1h
];
R
RRkRVMHO0FBMRm51]ZH:RMmRBv upXRR2skC0sBMRmpvu HXR#R
RRRRRR-R-R#7CObsH0MHF:R
RRRRRR-R-RRRRRRRR1RCCVOkM0MHFRO8CDNNs0MHFRRHMQ   R810R(4jn-3.4ngg
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRRMhFCR
RRCRLo
HMRRRRRRRR-t-RCP0RNCDkRsVFRC#bODHNR#ONCR#
RRRRRHRRVRR5Z 3)Rj=R32jRRC0EMR
RRRRRRRRRRRRRRVRHRZ5R3RQv=3RjjRR20MEC
RRRRRRRRRRRRRRRRRRRRRRRR0sCkRsMv]qa_qBA14 _;R
RRRRRRRRRRRRRRMRC8VRH;R

RRRRRRRRRRRRRHRRVRR5Zv3QRv=Rq_a]u2QRRC0EMR
RRRRRRRRRRRRRRRRRRRRRRCRs0MksRq-vaB]_A q1_
4;RRRRRRRRRRRRRRRRCRM8H
V;
RRRRRRRRRRRRRRRRRHV53RZQ=vRRavq]Q_u_ me)R_.FZsR3RQv=vR-q_a]umQ_e_ ).RR20MEC
RRRRRRRRRRRRRRRRRRRRRRRR0sCkRsMv]qa_ BZ)
m;RRRRRRRRRRRRRRRRCRM8H
V;RRRRRRRRCRM8H
V;
RRRRRRRRR--tRC0PkNDCFRVsCRoMNCsDNRO#RC
RRRRRsRRCs0kMmRBv upXB'5m51]Z 3)2m*B135ZQ,v2Rh1Q]35Z)* 215QhZv3Q2
2;RRRRCRM8B]m1;R

RVRRk0MOHRFMB]m15RZ:HBMRmpvu uX_m)pqRs2RCs0kMmRBv upXm_upRq)HR#
RRRRR-RR-CR7#HOsbF0HMR:
RRRRR-RR-RRRRRRRRC1CRMVkOF0HMCR8OsDNNF0HMMRHR Q  0R18jR4(.n3-g4gnR
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRR2RNR0)Ck#sMRvBmuXp _pumqj)53Rj,j23jRRFMCFsssR

RRRRRPRRNNsHLRDCZR4,Z:.RRvBmuXp ;R
RRRRRRNRPsLHNDZCRmRza:mRBv upXm_up;q)
RRRRoLCHRM
RRRRR-RR-ERBCRO	PHND8$H0RRFVHkMb0sRNoCklM
0#RRRRRRRRH5VRRqZ3)=tRRq-vau]_QRR20MEC
RRRRRRRRRRRRRRRR#N#CRs0w1qp R
RRRRRRRRRRRRRRRRRRRRRRRRRRCRsb0FsR3"ZqR)t=vR-q_a]uHQRMmRB1Z]52R"
RRRRRRRRRRRRRRRRRRRRRRRRR#RRCsPCHR0$ m)))R;
RRRRRRRRRRRRRsRRCs0kMmRBv upXm_up'q)5jj3,3Rjj
2;RRRRRRRRCRM8H
V;
RRRRRRRRR--BbFlkR0CPkNDCFRVsbR#CNOHDNRO#
C#RRRRRRRRH5VRRvZ3q=tRRjj3R8NMRqZ3)=tRRjj3R02RE
CMRRRRRRRRRRRRRRRRskC0sBMRmpvu uX_m)pq'354jj,R3;j2
RRRRRRRR8CMR;HV
R
RRRRRRVRHRZ5R3tvqRv=Rq_a]uNQRMZ8R3tq)Rv=Rq_a]umQ_e_ ).RR20MEC
RRRRRRRRRRRRRRRR0sCkRsMBumvp_ Xuqmp)4'53Rj,v]qa_2uQ;R
RRRRRRMRC8VRH;R

RRRRRHRRVRR5Zq3vtRR=v]qa__uQm)e _N.RMZ8R3tq)Rv=Rq_a]umQ_e_ ).RR20MEC
RRRRRRRRRRRRRRRR0sCkRsMBumvp_ Xuqmp)j'53Rj,j23j;R
RRRRRRMRC8VRH;R

RRRRRHRRVRR5Zq3vtRR=v]qa__uQm)e _N.RMZ8R3tq)R-=Rv]qa__uQm)e _2.RRC0EMR
RRRRRRRRRRRRRRCRs0MksRvBmuXp _pumq5)'j,3jRjj32R;
RRRRRCRRMH8RV
;
RRRRRRRR-B-RFklb0PCRNCDkRsVFRMoCCDsNR#ONCR
RRRRRR4RZRR:=uqmp)m_a_vBmuXp 5;Z2
RRRRRRRRRZ.:B=Rmpvu 5X'B]m153Z4)* 2B5m1ZQ43vR2,1]Qh53Z4)* 215QhZQ43v;22
RRRRRRRRzZma=R:RvBmuXp __amuqmp).5Z2R;
RRRRRsRRCs0kMmRZz
a;RRRRCRM8B]m1;


RRRR-R-
R-RR-sRqHl0ECO0HRCmbsFN0sR#
R-RR-R
RRkRVMHO0F"MR+5"RRRp:HBMRmpvu RX;RR):HBMRmpvu 2XRR0sCkRsMBumvpR XHR#
RRRRR-RR-CR7#HOsbF0HMR:
RRRRR-RR-RRRRRRRRC1CRMVkOF0HMCR8OsDNNF0HMMRHR Q  0R18jR4(.n3-g4gnR
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRRFRhMRC
RLRRCMoH
RRRRRRRR0sCkRsMBumvp' X5)p3 RR+) 3),3RpQ+vRRQ)3v
2;RRRRCRM8";+"
R
RRkRVMHO0F"MR+5"RRRp:H)MR ;qpRR):HBMRmpvu 2XRR0sCkRsMBumvpR XHR#
RRRRR-RR-CR7#HOsbF0HMR:
RRRRR-RR-RRRRRRRRC1CRMVkOF0HMCR8OsDNNF0HMMRHR Q  0R18jR4(.n3-g4gnR
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRRFRhMRC
RLRRCMoH
RRRRRRRR0sCkRsMBumvp' X5+pRR))3 ),R32Qv;R
RRMRC8+R""
;
RRRRVOkM0MHFR""+Rp5R:MRHRvBmuXp ;)RR:MRHRq) pRR2RsRRCs0kMmRBv upX#RH
RRRRRRRRR--7OC#s0HbH:FM
RRRRRRRRR--RRRRR1RRCVCRk0MOHRFM8DCON0sNHRFMHQMR R  1R084nj(34.-g
gnRRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRhCFM
RRRRoLCHRM
RRRRRsRRCs0kMmRBv upXp'53R) +,R)RQp3v
2;RRRRCRM8";+"
R
RRkRVMHO0F"MR+5"RpH:RMmRBv upXm_up;q)RR):HBMRmpvu uX_m)pq2R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRCRs0MksRvBmuXp _pumqH)R#R
RRRRRR-R-R#7CObsH0MHF:R
RRRRRR-R-RRRRRRRR1RCCVOkM0MHFRO8CDNNs0MHFRRHMQ   R810R(4jn-3.4ngg
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRRRN2)kC0sRM#Bumvp_ Xuqmp)j'53Rj,j23jRRFMCFsssR
RRRRRR-R-
RRRRRRRRsPNHDNLCpRZ,)RZRB:Rmpvu 
X;RRRRRRRRPHNsNCLDRzZmaRR:Bumvp_ Xuqmp)R;
RLRRCMoH
RRRRRRRRR--BOEC	NRPDHH80F$RVMRHbRk0Nksol0CM#R
RRRRRRVRHRp5R3tq)R-=Rv]qa_RuQ2ER0CRM
RRRRRRRRRRRRRNRR#s#C0qRwp
1 RRRRRRRRRRRRRRRRRRRRRRRRRRRRsFCbs"0Rp)3qtRR=-avq]Q_uRRHM+,5p)
2"RRRRRRRRRRRRRRRRRRRRRRRRRRRR#CCPs$H0R) )m
);RRRRRRRRRRRRRRRRskC0sBMRmpvu uX_m)pq'35jjj,R3;j2
RRRRRRRR8CMR;HV
R

RRRRRHRRVRR5))3qtRR=-avq]Q_uR02RE
CMRRRRRRRRRRRRRRRRNC##sw0Rq p1
RRRRRRRRRRRRRRRRRRRRRRRRRRRRbsCFRs0"q)3)=tRRq-vau]_QMRHRp+5,")2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRP#CC0sH$)R );m)
RRRRRRRRRRRRRRRR0sCkRsMBumvp_ Xuqmp)j'53Rj,j23j;R
RRRRRRMRC8VRH;R

RRRRR-RR-CRt0sRbHHMObRNDPkNDCR
RRRRRRpRZRR:=uqmp)m_a_vBmuXp 5RRp2R;
RRRRRZRR)=R:Rpumqa)_mm_Bv upX)5RR
2;RRRRRRRRZamzRR:=Bumvp_ Xaum_m)pq5vBmuXp 'p5Z3R) +)RZ3,) R3ZpQ+vRZQ)3v;22
RRRRRRRR0sCkRsMZamz;R
RRMRC8+R""
;
RRRRVOkM0MHFR""+Rp5R:MRHRq) pR;R)H:RMmRBv upXm_up2q)R0sCkRsMBumvp_ Xuqmp)#RH
RRRRRRRRR--7OC#s0HbH:FM
RRRRRRRRR--RRRRR1RRCVCRk0MOHRFM8DCON0sNHRFMHQMR R  1R084nj(34.-g
gnRRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRN)2RCs0kMB#Rmpvu uX_m)pq'35jjj,R3Rj2FCMRsssF
RRRRRRRRsPNHDNLC)RZRB:Rmpvu 
X;RRRRRRRRPHNsNCLDRzZmaRR:Bumvp_ Xuqmp)R;
RLRRCMoH
RRRRRRRRR--BOEC	NRPDHH80F$RVMRHbRk0Nksol0CM#R
RRRRRRVRHR)5R3tq)R-=Rv]qa_RuQ2ER0CRM
RRRRRRRRRRRRRNRR#s#C0qRwp
1 RRRRRRRRRRRRRRRRRRRRRRRRRRRRsFCbs"0R))3qtRR=-avq]Q_uRRHM+,5p)
2"RRRRRRRRRRRRRRRRRRRRRRRRRRRR#CCPs$H0R) )m
);RRRRRRRRRRRRRRRRskC0sBMRmpvu uX_m)pq'35jjj,R3;j2
RRRRRRRR8CMR;HV
R
RRRRRR-R-R0tCRHbsMbOHNPDRNCDk
RRRRRRRRRZ):u=Rm)pq__amBumvp5 XR2)R;R
RRRRRRmRZz:aR=mRBv upXm_a_pumqB)5mpvu 5X'pRR+Z))3 Z,R)v3Q2
2;RRRRRRRRskC0sZMRm;za
RRRR8CMR""+;R

RVRRk0MOHRFM"R+"5:RpRRHMBumvp_ Xuqmp)R;R)H:RM R)qRp2skC0sBMRmpvu uX_m)pqR
H#RRRRRRRR-7-RCs#OHHb0F
M:RRRRRRRR-R-RRRRRRCR1CkRVMHO0F8MRCNODsHN0FHMRM RQ 1 R048Rj3(n.g-4gRn
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRNRR2CR)0Mks#mRBv upXm_up'q)5jj3,3RjjF2RMsRCs
FsRRRRRRRR-R-
RRRRRPRRNNsHLRDCZ:pRRvBmuXp ;R
RRRRRRNRPsLHNDZCRmRza:mRBv upXm_up;q)
RRRRoLCHRM
RRRRR-RR-ERBCRO	PHND8$H0RRFVHkMb0sRNoCklM
0#RRRRRRRRH5VRRqp3)=tRRq-vau]_QRR20MEC
RRRRRRRRRRRRRRRR#N#CRs0w1qp R
RRRRRRRRRRRRRRRRRRRRRRRRRRCRsb0FsR3"pqR)t=vR-q_a]uHQRM5R+p2,)"R
RRRRRRRRRRRRRRRRRRRRRRRRRRCR#PHCs0 $R)))m;R
RRRRRRRRRRRRRRCRs0MksRvBmuXp _pumq5)'j,3jRjj32R;
RRRRRCRRMH8RV
;
RRRRRRRR-t-RCb0RsOHMHDbNRDPNkRC
RRRRRZRRp=R:Rpumqa)_mm_Bv upXp5RR
2;RRRRRRRRZamzRR:=Bumvp_ Xaum_m)pq5vBmuXp 'p5Z3R) +,R)R3ZpQ2v2;R
RRRRRRCRs0MksRzZmaR;
RCRRM"8R+
";
RRRRMVkOF0HM-R""RR5pH:RMmRBv upXR;R)H:RMmRBv upXRR2skC0sBMRmpvu HXR#R
RRRRRR-R-R#7CObsH0MHF:R
RRRRRR-R-RRRRRRRR1RCCVOkM0MHFRO8CDNNs0MHFRRHMQ   R810R(4jn-3.4ngg
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRRMhFCR
RRCRLo
HMRRRRRRRRskC0sBMRmpvu 5X'p 3)R)-R3,) RQp3vRR-)v3Q2R;
RCRRM"8R-
";
RRRRMVkOF0HM-R""RR5pH:RM R)qRp;RRRR)H:RMmRBv upXRR2skC0sBMRmpvu HXR#R
RRRRRR-R-R#7CObsH0MHF:R
RRRRRR-R-RRRRRRRR1RCCVOkM0MHFRO8CDNNs0MHFRRHMQ   R810R(4jn-3.4ngg
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRRMhFCR
RRCRLo
HMRRRRRRRRskC0sBMRmpvu 5X'pRR-) 3),4R-3*jRRQ)3v
2;RRRRCRM8";-"
R
RRkRVMHO0F"MR-5"RRRp:HBMRmpvu RX;RR):H)MR Rqp2RRRR0sCkRsMBumvpR XHR#
RRRRR-RR-CR7#HOsbF0HMR:
RRRRR-RR-RRRRRRRRC1CRMVkOF0HMCR8OsDNNF0HMMRHR Q  0R18jR4(.n3-g4gnR
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRRFRhMRC
RLRRCMoH
RRRRRRRR0sCkRsMBumvp' X5)p3 RR-)p,R32Qv;R
RRMRC8-R""
;
RRRRVOkM0MHFR""-Rp5R:MRHRvBmuXp _pumqR);)H:RMmRBv upXm_up2q)
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR0sCkRsMBumvp_ Xuqmp)#RH
RRRRRRRRR--7OC#s0HbH:FM
RRRRRRRRR--RRRRR1RRCVCRk0MOHRFM8DCON0sNHRFMHQMR R  1R084nj(34.-g
gnRRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRN)2RCs0kMB#Rmpvu uX_m)pq'35jjj,R3Rj2FCMRsssF
RRRRRRRR
--RRRRRRRRPHNsNCLDR,ZpRRZ):mRBv upXR;
RRRRRPRRNNsHLRDCZamzRB:Rmpvu uX_m)pq;R
RRCRLo
HMRRRRRRRR-B-RE	CORDPNH08H$VRFRbHMkN0RslokC#M0
RRRRRRRRRHV53RpqR)t=vR-q_a]u2QRRC0EMR
RRRRRRRRRRRRRR#RN#0CsRpwq1R 
RRRRRRRRRRRRRRRRRRRRRRRRRsRRCsbF0pR"3tq)R-=Rv]qa_RuQH-MR5)p,2R"
RRRRRRRRRRRRRRRRRRRRRRRRR#RRCsPCHR0$ m)))R;
RRRRRRRRRRRRRsRRCs0kMmRBv upXm_up'q)5jj3,3Rjj
2;RRRRRRRRCRM8H
V;
RRRRRRRRRHV53R)qR)t=vR-q_a]u2QRRC0EMR
RRRRRRRRRRRRRR#RN#0CsRpwq1R 
RRRRRRRRRRRRRRRRRRRRRRRRRsRRCsbF0)R"3tq)R-=Rv]qa_RuQH-MR5)p,2R"
RRRRRRRRRRRRRRRRRRRRRRRRR#RRCsPCHR0$ m)))R;
RRRRRRRRRRRRRsRRCs0kMmRBv upXm_up'q)5jj3,3Rjj
2;RRRRRRRRCRM8H
V;RRRRRRRR-t-RCb0RsOHMHDbNRDPNkRC
RRRRRZRRp=R:Rpumqa)_mm_Bv upXp5RR
2;RRRRRRRRZ:)R=mRup_q)aBm_mpvu RX5);R2
RRRRRRRRzZma=R:RvBmuXp __amuqmp)m5Bv upXZ'5p 3)RZ-R) 3),pRZ3RQv-3Z)Q2v2;R
RRRRRRCRs0MksRzZmaR;
RCRRM"8R-
";
RRRRMVkOF0HM-R""RR5pH:RM R)qRp;RR):HBMRmpvu uX_m)pq2CRs0MksRvBmuXp _pumqH)R#R
RRRRRR-R-R#7CObsH0MHF:R
RRRRRR-R-RRRRRRRR1RCCVOkM0MHFRO8CDNNs0MHFRRHMQ   R810R(4jn-3.4ngg
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRRRN2)kC0sRM#Bumvp_ Xuqmp)j'53Rj,j23jRRFMCFsssR
RRRRRR-R-
RRRRRRRRsPNHDNLC)RZRB:Rmpvu 
X;RRRRRRRRPHNsNCLDRzZmaRR:Bumvp_ Xuqmp)R;
RLRRCMoH
RRRRRRRRR--BOEC	NRPDHH80F$RVMRHbRk0Nksol0CM#R
RRRRRRVRHR)5R3tq)R-=Rv]qa_RuQ2ER0CRM
RRRRRRRRRRRRRNRR#s#C0qRwp
1 RRRRRRRRRRRRRRRRRRRRRRRRRRRRsFCbs"0R))3qtRR=-avq]Q_uRRHM-,5p)
2"RRRRRRRRRRRRRRRRRRRRRRRRRRRR#CCPs$H0R) )m
);RRRRRRRRRRRRRRRRskC0sBMRmpvu uX_m)pq'35jjj,R3;j2
RRRRRRRR8CMR;HV
R
RRRRRR-R-R0tCRHbsMbOHNPDRNCDk
RRRRRRRRRZ):u=Rm)pq__amBumvp5 XR2)R;R
RRRRRRmRZz:aR=mRBv upXm_a_pumqB)5mpvu 5X'pRR-Z))3 -,R4*3jZQ)3v;22
RRRRRRRR0sCkRsMZamz;R
RRMRC8-R""
;
RRRRVOkM0MHFR""-Rp5R:MRHRvBmuXp _pumqR);RR):H)MR 2qpR0sCkRsMBumvp_ Xuqmp)#RH
RRRRRRRRR--7OC#s0HbH:FM
RRRRRRRRR--RRRRR1RRCVCRk0MOHRFM8DCON0sNHRFMHQMR R  1R084nj(34.-g
gnRRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRN)2RCs0kMB#Rmpvu uX_m)pq'35jjj,R3Rj2FCMRsssF
RRRRRRRR
--RRRRRRRRPHNsNCLDRRZp:mRBv upXR;
RRRRRPRRNNsHLRDCZamzRB:Rmpvu uX_m)pq;R
RRCRLo
HMRRRRRRRR-B-RE	CORDPNH08H$VRFRbHMkN0RslokC#M0
RRRRRRRRRHV53RpqR)t=vR-q_a]u2QRRC0EMR
RRRRRRRRRRRRRR#RN#0CsRpwq1R 
RRRRRRRRRRRRRRRRRRRRRRRRRsRRCsbF0pR"3tq)R-=Rv]qa_RuQH-MR5)p,2R"
RRRRRRRRRRRRRRRRRRRRRRRRR#RRCsPCHR0$ m)))R;
RRRRRRRRRRRRRsRRCs0kMmRBv upXm_up'q)5jj3,3Rjj
2;RRRRRRRRCRM8H
V;
RRRRRRRRR--tRC0bMsHONHbDNRPD
kCRRRRRRRRZ:pR=mRup_q)aBm_mpvu RX5p;R2
RRRRRRRRzZma=R:RvBmuXp __amuqmp)m5Bv upXZ'5p 3)R)-R,pRZ32Qv2R;
RRRRRsRRCs0kMmRZz
a;RRRRCRM8";-"
R

RVRRk0MOHRFM"R*"5:RpRRHMBumvp; XR:R)RRHMBumvpR X2CRs0MksRvBmuXp R
H#RRRRRRRR-7-RCs#OHHb0F
M:RRRRRRRR-R-RRRRRRCR1CkRVMHO0F8MRCNODsHN0FHMRM RQ 1 R048Rj3(n.g-4gRn
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRhRRF
MCRRRRLHCoMR
RRRRRRCRs0MksRvBmuXp '35p)* RR))3 RR-pv3QR)*R3,QvR)p3 RR*)v3QRp+R3RQv*3R)); 2
RRRR8CMR""*;


RRRRVOkM0MHFR""*Rp5R:MRHRq) pR;R)H:RMmRBv upXRR2skC0sBMRmpvu HXR#R
RRRRRR-R-R#7CObsH0MHF:R
RRRRRR-R-RRRRRRRR1RCCVOkM0MHFRO8CDNNs0MHFRRHMQ   R810R(4jn-3.4ngg
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRRMhFCR
RRCRLo
HMRRRRRRRRskC0sBMRmpvu 5X'pRR*) 3),RRp*3R)Q;v2
RRRR8CMR""*;R

RVRRk0MOHRFM"R*"5:RpRRHMBumvp; XR:R)RRHM)p qRR2RRCRs0MksRvBmuXp R
H#RRRRRRRR-7-RCs#OHHb0F
M:RRRRRRRR-R-RRRRRRCR1CkRVMHO0F8MRCNODsHN0FHMRM RQ 1 R048Rj3(n.g-4gRn
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRhRRF
MCRRRRLHCoMR
RRRRRRCRs0MksRvBmuXp '35p)* RRR),pv3QR)*R2R;
RCRRM"8R*
";
RRRRMVkOF0HM*R""RR5pH:RMmRBv upXm_up;q)RR):HBMRmpvu uX_m)pq2R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRCRs0MksRvBmuXp _pumqH)R#R
RRRRRR-R-R#7CObsH0MHF:R
RRRRRR-R-RRRRRRRR1RCCVOkM0MHFRO8CDNNs0MHFRRHMQ   R810R(4jn-3.4ngg
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRRRN2)kC0sRM#Bumvp_ Xuqmp)j'53Rj,j23jRRFMCFsssR
RRRRRR-R-
RRRRRRRRsPNHDNLCmRZz:aRRvBmuXp _pumq
);RRRRLHCoMR
RRRRRR-R-RCBEOP	RN8DHHR0$FHVRM0bkRoNskMlC0R#
RRRRRHRRVRR5p)3qtRR=-avq]Q_uR02RE
CMRRRRRRRRRRRRRRRRNC##sw0Rq p1
RRRRRRRRRRRRRRRRRRRRRRRRRRRRbsCFRs0"qp3)=tRRq-vau]_QMRHRp*5,")2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRP#CC0sH$)R );m)
RRRRRRRRRRRRRRRR0sCkRsMBumvp_ Xuqmp)j'53Rj,j23j;R
RRRRRRMRC8VRH;R

RRRRRHRRVRR5))3qtRR=-avq]Q_uR02RE
CMRRRRRRRRRRRRRRRRNC##sw0Rq p1
RRRRRRRRRRRRRRRRRRRRRRRRRRRRbsCFRs0"q)3)=tRRq-vau]_QMRHRp*5,")2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRP#CC0sH$)R );m)
RRRRRRRRRRRRRRRR0sCkRsMBumvp_ Xuqmp)j'53Rj,j23j;R
RRRRRRMRC8VRH;R

RRRRR-RR-CRt0sRbHHMObRNDPkNDCR
RRRRRRmRZzva3q:tR=3RpvRqt*3R)v;qt
RRRRRRRRzZma)3qt=R:Rat _Qu)huBQqep_q pz5qp3)+tRRq)3);t2
R
RRRRRRCRs0MksRzZmaR;
RCRRM"8R*
";
RRRRMVkOF0HM*R""RR5pH:RM R)qRp;RR):HBMRmpvu uX_m)pq2CRs0MksRvBmuXp _pumqH)R#R
RRRRRR-R-R#7CObsH0MHF:R
RRRRRR-R-RRRRRRRR1RCCVOkM0MHFRO8CDNNs0MHFRRHMQ   R810R(4jn-3.4ngg
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRRRN2)kC0sRM#Bumvp_ Xuqmp)j'53Rj,j23jRRFMCFsssR
RRRRRR-R-
RRRRRRRRRRRRsPNHDNLCpRZRB:Rmpvu uX_m)pq;R
RRRRRRNRPsLHNDZCRmRza:mRBv upXm_up;q)
RRRRoLCHRM
RRRRR-RR-ERBCRO	PHND8$H0RRFVHkMb0sRNoCklM
0#RRRRRRRRH5VRRq)3)=tRRq-vau]_QRR20MEC
RRRRRRRRRRRRRRRR#N#CRs0w1qp R
RRRRRRRRRRRRRRRRRRRRRRRRRRCRsb0FsR3")qR)t=vR-q_a]uHQRM5R*p2,)"R
RRRRRRRRRRRRRRRRRRRRRRRRRRCR#PHCs0 $R)))m;R
RRRRRRRRRRRRRRCRs0MksRvBmuXp _pumq5)'j,3jRjj32R;
RRRRRCRRMH8RV
;
RRRRRRRR-t-RCb0RsOHMHDbNRDPNkRC
RRRRRZRRpq3vt=R:R1umQeaQ  _)q5p'q5A1p;22
RRRRRRRRRHV5RRp<3RjjRR20MEC
RRRRRRRRRRRRRRRR3ZpqR)t:v=Rq_a]u
Q;RRRRRRRRCCD#
RRRRRRRRRRRRRRRR3ZpqR)t:j=R3
j;RRRRRRRRCRM8H
V;
RRRRRRRRzZmaq3vt=R:R3ZpvRqt*3R)v;qt
RRRRRRRRzZma)3qt=R:Rat _Qu)huBQqep_q pz53ZpqR)t+3R)q2)t;R

RRRRRsRRCs0kMmRZz
a;RRRRCRM8";*"
R
RRkRVMHO0F"MR*5"RRRp:HBMRmpvu uX_m)pq;)RR:MRHRq) ps2RCs0kMmRBv upXm_upRq)HR#
RRRRR-RR-CR7#HOsbF0HMR:
RRRRR-RR-RRRRRRRRC1CRMVkOF0HMCR8OsDNNF0HMMRHR Q  0R18jR4(.n3-g4gnR
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRR2RNR0)Ck#sMRvBmuXp _pumq5)'j,3jRjj32MRFRsCsFRs
RRRRR-RR-R
RRRRRRNRPsLHNDZCR)RR:Bumvp_ Xuqmp)R;
RRRRRPRRNNsHLRDCZamzRB:Rmpvu uX_m)pq;R
RRCRLo
HMRRRRRRRR-B-RE	CORDPNH08H$VRFRbHMkN0RslokC#M0
RRRRRRRRRHV53RpqR)t=vR-q_a]u2QRRC0EMR
RRRRRRRRRRRRRR#RN#0CsRpwq1R 
RRRRRRRRRRRRRRRRRRRRRRRRRsRRCsbF0pR"3tq)R-=Rv]qa_RuQH*MR5)p,2R"
RRRRRRRRRRRRRRRRRRRRRRRRR#RRCsPCHR0$ m)))R;
RRRRRRRRRRRRRsRRCs0kMmRBv upXm_up'q)5jj3,3Rjj
2;RRRRRRRRCRM8H
V;
RRRRRRRRR--tRC0bMsHONHbDNRPD
kCRRRRRRRRZv)3q:tR=mRu1QQae) _ 'qp51qA52)2;R
RRRRRRVRHR)5RRj<R32jRRC0EMR
RRRRRRRRRRRRRR)RZ3tq)RR:=v]qa_;uQ
RRRRRRRR#CDCR
RRRRRRRRRRRRRR)RZ3tq)RR:=j;3j
RRRRRRRR8CMR;HV
R
RRRRRRmRZzva3q:tR=3RpvRqt*)RZ3tvq;R
RRRRRRmRZzqa3):tR= Rta)_uQQhBu_qpezqp 35pqR)t+)RZ3tq)2
;
RRRRRRRRskC0sZMRm;za
RRRR8CMR""*;R

RkRVMHO0F"MR/5"RRRp:HBMRmpvu RX;RR):HBMRmpvu 2XRR0sCkRsMBumvpR XHR#
RRRRR-RR-CR7#HOsbF0HMR:
RRRRR-RR-RRRRRRRRC1CRMVkOF0HMCR8OsDNNF0HMMRHR Q  0R18jR4(.n3-g4gnR
RRRRRR-R-R0hFC
#:RRRRRRRR-R-RRRRRR2RNR0)Ck#sMRvBmuXp ' 5)q]p'Q,t]Rjj32MRFRsCsFRs
RRRRR-RR-R
RRRRRRNRPsLHNDaCR Rvu: R)q:pR=3R))) *3R) +3R)Q)v*3;Qv
RRRLHCoMR
RRRRRR-R-RCBEOP	RN8DHHR0$FHVRM0bkRoNskMlC0R#
RRRRRHRRVaR5 Rvu=3Rjj02RE
CMRRRRRRRRRRRRRRRRR#N#CRs0w1qp R
RRRRRRRRRRRRRRRRRRRRRRCRsb0FsR0"q0bCl0FR0RP8HHR8CBumvpR XL5$Rj,3jRjj32R"
RRRRRRRRRRRRRRRRRRRRR#RRCsPCHR0$ m)))R;
RRRRRRRRRRRRRRRRskC0sBMRmpvu 5X')p q't]Q]j,R3;j2
RRRRRRRR8CMR;HV
R
RRRRRR-R-R0tCRDPNkRC
RRRRRsRRCs0kMmRBv upXR'55)p3 RR*) 3)Rp+R3RQv*3R)QRv2/ Rav
u,RRRRRRRRRRRRRRRRRRRRRRRRR35pQ*vRR))3 RR-p 3)R)*R32QvRa/R 2vu;R
RRMRC8/R""
;
RVRRk0MOHRFM"R/"5:RpRRHM)p q;)RR:MRHRvBmuXp Rs2RCs0kMmRBv upX#RH
RRRRRRRRR--7OC#s0HbH:FM
RRRRRRRRR--RRRRR1RRCVCRk0MOHRFM8DCON0sNHRFMHQMR R  1R084nj(34.-g
gnRRRRRRRR-h-RF#0C:R
RRRRRR-R-RRRRRRRRN)2RCs0kMB#Rmpvu 5X')p q't]Q]j,R3Rj2FCMRsssF
RRRRRRRR
--RRRRRRRRPHNsNCLDRva uRR:)p qRR:=) 3)*))3 RR+)v3Q*Q)3vR;
RLRRCMoH
RRRRRRRRR--BOEC	NRPDHH80F$RVMRHbRk0Nksol0CM#R
RRRRRRVRHR 5av=uRRjj32ER0CRM
RRRRRRRRRRRRRRRRNC##sw0Rq p1
RRRRRRRRRRRRRRRRRRRRRRRRbsCFRs0"0q0C0lbRR0F8HHP8BCRmpvu LXR$jR53Rj,j23j"R
RRRRRRRRRRRRRRRRRRRRRRCR#PHCs0 $R)))m;R
RRRRRRRRRRRRRRsRRCs0kMmRBv upX)'5 'qp]]Qt,3Rjj
2;RRRRRRRRCRM8H
V;
RRRRRRRRR--tRC0PkNDCR
RRRRRR Rav:uR=RRp/ Rav
u;RRRRRRRRskC0sRMRBumvp' X5 Rav*uRR))3 -,Rau vR)*R3RQv2R;
RCRRM"8R/
";
RRRRMVkOF0HM/R""RR5pH:RMmRBv upXR;R)H:RM R)q2pRRRRRskC0sBMRmpvu HXR#R
RRRRRR-R-R#7CObsH0MHF:R
RRRRRR-R-RRRRRRRR1RCCVOkM0MHFRO8CDNNs0MHFRRHMQ   R810R(4jn-3.4ngg
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRRRN2)kC0sRM#Bumvp' X5q) pQ']tR],j23jRRFMCFsssR
RRCRLo
HMRRRRRRRR-B-RE	CORDPNH08H$VRFRbHMkN0RslokC#M0
RRRRRRRRRHV5=)RRjj32ER0CRM
RRRRRRRRRRRRRRRRNC##sw0Rq p1
RRRRRRRRRRRRRRRRRRRRRRRRbsCFRs0"0q0C0lbRR0F8HHP8BCRmpvu LXR$3RjjR"
RRRRRRRRRRRRRRRRRRRRR#RRCsPCHR0$ m)))R;
RRRRRRRRRRRRRRRRskC0sBMRmpvu 5X')p q't]Q]j,R3;j2
RRRRRRRR8CMR;HV
R
RRRRRR-R-R0tCRDPNkRC
RRRRRsRRCs0kMmRBv upXp'53R) /,R)RQp3vRR/)
2;RRRRCRM8";/"
R

RVRRk0MOHRFM"R/"5:RpRRHMBumvp_ Xuqmp));R:MRHRvBmuXp _pumq
)2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRskC0sBMRmpvu uX_m)pqR
H#RRRRRRRR-7-RCs#OHHb0F
M:RRRRRRRR-R-RRRRRRCR1CkRVMHO0F8MRCNODsHN0FHMRM RQ 1 R048Rj3(n.g-4gRn
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRNRR2CR)0Mks#mRBv upXm_up'q)5q) pQ']tR],j23jRRFMCFsssR
RRRRRR-R-
RRRRRRRRsPNHDNLCmRZz:aRRvBmuXp _pumq
);RRRRLHCoMR
RRRRRR-R-RCBEOP	RN8DHHR0$FHVRM0bkRoNskMlC0R#
RRRRRHRRV)R53tvqRj=R3Rj20MEC
RRRRRRRRRRRRRRRR#N#CRs0w1qp R
RRRRRRRRRRRRRRRRRRRRRRCRsb0FsR0"q0bCl0FR0RP8HHR8CBumvp_ Xuqmp)$RLR35jjj,R3"j2
RRRRRRRRRRRRRRRRRRRRRRRRP#CC0sH$)R );m)
RRRRRRRRRRRRRRRR0sCkRsMBumvp_ Xuqmp))'5 'qp]]Qt,3Rjj
2;RRRRRRRRCRM8H
V;
RRRRRRRRRHV53RpqR)t=vR-q_a]u2QRRC0EMR
RRRRRRRRRRRRRR#RN#0CsRpwq1R 
RRRRRRRRRRRRRRRRRRRRRsRRCsbF0pR"3tq)R-=Rv]qa_RuQH/MR5)p,2R"
RRRRRRRRRRRRRRRRRRRRR#RRCsPCHR0$ m)))R;
RRRRRRRRRRRRRsRRCs0kMmRBv upXm_up'q)5q) pQ']tR],j23j;R
RRRRRRMRC8VRH;R

RRRRRHRRVRR5))3qtRR=-avq]Q_uR02RE
CMRRRRRRRRRRRRRRRRNC##sw0Rq p1
RRRRRRRRRRRRRRRRRRRRRRRRbsCFRs0"q)3)=tRRq-vau]_QMRHRp/5,")2
RRRRRRRRRRRRRRRRRRRRRRRRP#CC0sH$)R );m)
RRRRRRRRRRRRRRRR0sCkRsMBumvp_ Xuqmp)j'53Rj,j23j;R
RRRRRRMRC8VRH;R

RRRRR-RR-CRt0sRbHHMObRNDPkNDCR
RRRRRRmRZzva3q:tR=3Rpv/qt)q3vtR;
RRRRRZRRm3zaqR)t:t=R ua_)BQhQpuq_peqzp 53tq)R)-R3tq)2
;
RRRRRRRRskC0sZMRm;za
RRRR8CMR""/;R

RVRRk0MOHRFM"R/"5:RpRRHMBumvp_ Xuqmp)R;R)H:RM R)qRp2skC0sBMRmpvu uX_m)pqR
H#RRRRRRRR-7-RCs#OHHb0F
M:RRRRRRRR-R-RRRRRRCR1CkRVMHO0F8MRCNODsHN0FHMRM RQ 1 R048Rj3(n.g-4gRn
RRRRR-RR-FRh0:C#
RRRRRRRRR--RRRRRNRR2CR)0Mks#mRBv upXm_up'q)5q) pQ']tR],j23jRRFMCFsssR
RRRRRR-R-
RRRRRRRRsPNHDNLC)RZRB:Rmpvu uX_m)pq;R
RRRRRRNRPsLHNDZCRmRza:mRBv upXm_up;q)
RRRRoLCHRM
RRRRR-RR-ERBCRO	PHND8$H0RRFVHkMb0sRNoCklM
0#RRRRRRRRH5VR)RR=j23jRC0EMR
RRRRRRRRRRRRRR#RN#0CsRpwq1R 
RRRRRRRRRRRRRRRRRRRRRsRRCsbF0qR"0l0Cb00RFHR8PCH8RvBmuXp _pumqL)R$3RjjR"
RRRRRRRRRRRRRRRRRRRRR#RRCsPCHR0$ m)))R;
RRRRRRRRRRRRRsRRCs0kMmRBv upXm_up'q)5q) pQ']tR],j23j;R
RRRRRRMRC8VRH;R

RRRRRHRRVRR5p)3qtRR=-avq]Q_uR02RE
CMRRRRRRRRRRRRRRRRNC##sw0Rq p1
RRRRRRRRRRRRRRRRRRRRRRRRbsCFRs0"qp3)=tRRq-vau]_QMRHRp/5,")2
RRRRRRRRRRRRRRRRRRRRRRRRP#CC0sH$)R );m)
RRRRRRRRRRRRRRRR0sCkRsMBumvp_ Xuqmp))'5 'qp]]Qt,3Rjj
2;RRRRRRRRCRM8H
V;
RRRRRRRRR--tRC0bMsHONHbDNRPD
kCRRRRRRRRZv)3q:tR=mRu1QQae) _ 'qp51qA52)2;R
RRRRRRVRHR<)RRjj3RC0EMR
RRRRRRRRRRRRRR)RZ3tq)RR:=v]qa_;uQ
RRRRRRRR#CDCR
RRRRRRRRRRRRRR)RZ3tq)RR:=j;3j
RRRRRRRR8CMR;HV
R
RRRRRRmRZzva3q:tR=3Rpv/qtZv)3q
t;RRRRRRRRZamz3tq)RR:=t_ auh)QBqQupq_ep5z p)3qtRR-Zq)3);t2
R
RRRRRRCRs0MksRzZmaR;
RCRRM"8R/
";
RRRRMVkOF0HM/R""RR5pH:RM R)qRp;RR):HBMRmpvu uX_m)pq2CRs0MksRvBmuXp _pumqH)R#R
RRRRRR-R-R#7CObsH0MHF:R
RRRRRR-R-RRRRRRRR1RCCVOkM0MHFRO8CDNNs0MHFRRHMQ   R810R(4jn-3.4ngg
RRRRRRRRR--hCF0#R:
RRRRR-RR-RRRRRRRRRN2)kC0sRM#Bumvp_ Xuqmp))'5 'qp]]Qt,3RjjF2RMsRCs
FsRRRRRRRR-R-
RRRRRPRRNNsHLRDCZ:pRRvBmuXp _pumq
);RRRRRRRRPHNsNCLDRzZmaRR:Bumvp_ Xuqmp)R;
RLRRCMoH
RRRRRRRRR--BOEC	NRPDHH80F$RVMRHbRk0Nksol0CM#R
RRRRRRVRHR35)vRqt=3Rjj02RE
CMRRRRRRRRRRRRRRRRNC##sw0Rq p1
RRRRRRRRRRRRRRRRRRRRRRRRbsCFRs0"0q0C0lbRR0F8HHP8BCRmpvu uX_m)pqRRL$5jj3,3Rjj
2"RRRRRRRRRRRRRRRRRRRRRRRR#CCPs$H0R) )m
);RRRRRRRRRRRRRRRRskC0sBMRmpvu uX_m)pq' 5)q]p'Q,t]Rjj32R;
RRRRRCRRMH8RV
;
RRRRRRRRH5VRRq)3)=tRRq-vau]_QRR20MEC
RRRRRRRRRRRRRRRR#N#CRs0w1qp R
RRRRRRRRRRRRRRRRRRRRRRCRsb0FsR3")qR)t=vR-q_a]uMRHRp/5,")2
RRRRRRRRRRRRRRRRRRRRRRRRP#CC0sH$)R );m)
RRRRRRRRRRRRRRRR0sCkRsMBumvp_ Xuqmp)j'53Rj,j23j;R
RRRRRRMRC8VRH;R

RRRRR-RR-CRt0sRbHHMObRNDPkNDCR
RRRRRRpRZ3tvqRR:=uQm1a Qe_q) pq'5Ap152
2;RRRRRRRRHpVRRj<R30jRE
CMRRRRRRRRRRRRRRRRZqp3):tR=qRvau]_QR;
RRRRRCRRD
#CRRRRRRRRRRRRRRRRZqp3):tR=3RjjR;
RRRRRCRRMH8RV
;
RRRRRRRRZamz3tvqRR:=Zvp3q)t/3tvq;R
RRRRRRmRZzqa3):tR= Rta)_uQQhBu_qpezqp p5Z3tq)R)-R3tq)2
;
RRRRRRRRskC0sZMRm;za
RRRR8CMR""/;C

MR8Rv]qa_vBmuXp ;



