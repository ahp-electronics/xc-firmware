--******************************************************
@Ea--HC0D:RRRR_#LH_OCObFlFMMC0##_$PM3E
8R-k-q0sEF:RRR[FoDM-o
-MwkOF0HMH:RMN#0MN0H0NCRD0DREOCRC#DDRRFV0REC#HL_O#C_$PM3RLDHs$NsR-
-BbFlN:M$RHR1DFHOMkADCCRaOFEMDHFoCR#,Q3MO
Q--h:QaRRRRRLwCR,4URj.jU-
-)HCP#MHFR#]H0$Fs:-
-Roqkj.n,jR46BsFsCRO01QA_md_QBHRbMHR8s0COH3FMR$KNNl	kN1sRkNM8s3Nl
R--qjko(j,.4q6R818RA _7p_qY61jhR8NMR_1AwaQp 6)_j3h1RHAsNaMRN
H3-q-RkUo4,4.j68Rq8RC81_BpQzhuaQ_wp)a  N7R0H0sLFR0R_1AQ3.BwRHGlFHMs#RH##kC3NRK$kN	lRNs18kMNlsN3-
-*****************************************************
*
DsHLNRs$HCCCRk;
#HCRC3CC#_08DHFoO4_4nNc3D
D;
ObN	CNoRvBmu mhhRa1HN#
0H0sLCk0RM#$_NLDOL	_F:GRRFLFDMCN;0
N0LsHkR0C#_$MD_HLODCDRL:RFCFDN
M;Ns00H0LkCORG_blNR#:R0MsHoN;
0H0sLCk0RNLDOL	_FbG_Nb8_H:MRRs#0H;Mo
0N0skHL0#CR$LM_D	NO_GLFRRFVObFlFMMC0:#RRObN	CNoRRH#0Csk;0
N0LsHkR0C#_$MD_HLODCDRRFVObFlFMMC0:#RRObN	CNoRRH#0Csk;0
N0LsHkR0C)amz ]_a)tmz]q_wAB)QRL:RFCFDN
M;Ns00H0LkC7R1qh_Qu_za7q pYR 7:FRLFNDCMN;
0H0sLCk0Rq17_amzu_za7q pYR 7:FRLFNDCMN;
0H0sLCk0Rp1B_uQhzwa_Q pa)R 7:FRLFNDCMN;
0H0sLCk0Rp1B_pwQa  )7RR:LDFFC;NM
0N0skHL0QCR.BB_p7i_Q7eQ :)RR0HMCsoC;0
N0LsHkR0CQ_.BwmQw_A hR#:R0MsHoN;
0H0sLCk0R1a au_1)Rqv:0R#soHM;F
OlMbFCRM01BA_qY))RR
RRRRRRRRRb0Fs5RR
RRRRRRRRRRRRRBRRmRR:FRk0#_08DHFoO;RR
RRRRRRRRRRRRRRRRRQj:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRR4RQ:HRRM#RR0D8_FOoHRR;
RRRRRRRRRRRRRBRRQRR:HRMR#_08DHFoORR
RRRRRRRRRRRRR;R2
8CMRlOFbCFMM
0;
lOFbCFMM10RAq_B)_)YQvh_zRX
RRRRRRRRRMoCCOsHRB5R_QQhaRR:L_H0P0COFRs548RRF0IMF2RjRR2R;R
RRRRRRRRRb0Fs5RR
RRRRRRRRRRRRRORRN$ss_HHM0k_F0RR:R0FkR8#0_oDFH;OR
RRRRRRRRRRRRRRRRsONsH$_M_H0HRMR:HRRM#RR0D8_FOoHRR
RRRRRRRRRRRRRR
2;CRM8ObFlFMMC0
;
ObFlFMMC0AR1_apzcR
RRRRRRRRRoCCMsRHO5zRpah_QQ:aRR0LH_OPC05FsRR46RI8FMR0Fj22RRR;
RRRRRRRRRsbF0
5RRRRRRRRRRRRRRRRRm:RRR0FkR8#0_oDFH;OR
RRRRRRRRRRRRRRRRRQj:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRR4RQRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRRQRR.RR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRRQ:dRRRHMR8#0_oDFH
ORRRRRRRRRRRRRR2RR;M
C8FROlMbFC;M0
0N0skHL0GCRON_lbVRFR_1ApczaRO:RFFlbM0CMRRH#"0Dk"
;
ObFlFMMC0AR1_w7w
RRRRRRRRbRRF5s0RR
RRRRRRRRRRRRRRRRT:kRF00R#8F_DoRHO;R
RRRRRRRRRRRRRRRRB:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRRR7:MRHR0R#8F_DoRHO
RRRRRRRRRRRRRRR2C;
MO8RFFlbM0CM;O

FFlbM0CMR_1A71ww)R
RRRRRRRRRb0Fs5RR
RRRRRRRRRRRRRTRRRF:Rk#0R0D8_FOoHRR;
RRRRRRRRRRRRRBRRRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRR7RRRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRR)RRRH:RM#RR0D8_FOoHRR
RRRRRRRRRRRRRR
2;CRM8ObFlFMMC0
;
ObFlFMMC0AR1_w7w1R1
RRRRRRRRRsbF0
5RRRRRRRRRRRRRRRRRTRR:FRk0#_08DHFoO
R;RRRRRRRRRRRRRRRRBRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRR7RR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRR1RR:HRMR#_08DHFoORR
RRRRRRRRRRRRR;R2
8CMRlOFbCFMM
0;
lOFbCFMM10RAw_7wR)
RRRRRRRRRsbF0
5RRRRRRRRRRRRRRRRRTRR:FRk0#_08DHFoO
R;RRRRRRRRRRRRRRRRBRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRR7RR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRR)RR:HRMR#_08DHFoORR
RRRRRRRRRRRRR;R2
8CMRlOFbCFMM
0;
lOFbCFMM10RAw_7wR1
RRRRRRRRRsbF0
5RRRRRRRRRRRRRRRRRTRR:FRk0#_08DHFoO
R;RRRRRRRRRRRRRRRRBRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRR7RR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRR1RR:HRMR#_08DHFoORR
RRRRRRRRRRRRR;R2
8CMRlOFbCFMM
0;
lOFbCFMM10RAw_7wR 
RRRRRRRRRsbF0
5RRRRRRRRRRRRRRRRRTRR:FRk0#_08DHFoO
R;RRRRRRRRRRRRRRRRBRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRR RR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRR7RR:HRMR#_08DHFoORR
RRRRRRRRRRRRR;R2
8CMRlOFbCFMM
0;
lOFbCFMM10RAw_7w) 1
RRRRRRRRbRRF5s0RR
RRRRRRRRRRRRRRRRT:kRF00R#8F_DoRHO;R
RRRRRRRRRRRRRRRRB:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRRR :MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRRR7:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRRR):MRHR0R#8F_DoRHO
RRRRRRRRRRRRRRR2C;
MO8RFFlbM0CM;O

FFlbM0CMR_1A7 ww1R1
RRRRRRRRRsbF0
5RRRRRRRRRRRRRRRRRTRR:FRk0#_08DHFoO
R;RRRRRRRRRRRRRRRRBRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRR RR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRR7RR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRR1RR:HRMR#_08DHFoORR
RRRRRRRRRRRRR;R2
8CMRlOFbCFMM
0;
lOFbCFMM10RAw_7w
 )RRRRRRRRRFRbsR05
RRRRRRRRRRRRRRRR:TRR0FkR8#0_oDFH;OR
RRRRRRRRRRRRRRRR:BRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRR: RRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRR:7RRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRR:)RRRHMR8#0_oDFH
ORRRRRRRRRRRRRR2RR;M
C8FROlMbFC;M0
F
OlMbFCRM017A_w1w 
RRRRRRRRbRRF5s0RR
RRRRRRRRRRRRRRRRT:kRF00R#8F_DoRHO;R
RRRRRRRRRRRRRRRRB:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRRR :MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRRR7:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRRR1:MRHR0R#8F_DoRHO
RRRRRRRRRRRRRRR2C;
MO8RFFlbM0CM;O

FFlbM0CMR_1A7hww
RRRRRRRRbRRF5s0RR
RRRRRRRRRRRRRRRRT:kRF00R#8F_DoRHO;R
RRRRRRRRRRRRRRRRB:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRRR7:MRHR0R#8F_DoRHO
RRRRRRRRRRRRRRR2C;
MO8RFFlbM0CM;O

FFlbM0CMR_1A7hww1R)
RRRRRRRRRsbF0
5RRRRRRRRRRRRRRRRRTRR:FRk0#_08DHFoO
R;RRRRRRRRRRRRRRRRBRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRR7RR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRR)RR:HRMR#_08DHFoORR
RRRRRRRRRRRRR;R2
8CMRlOFbCFMM
0;
lOFbCFMM10RAw_7w1h1
RRRRRRRRbRRF5s0RR
RRRRRRRRRRRRRRRRT:kRF00R#8F_DoRHO;R
RRRRRRRRRRRRRRRRB:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRRR7:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRRR1:MRHR0R#8F_DoRHO
RRRRRRRRRRRRRRR2C;
MO8RFFlbM0CM;O

FFlbM0CMR_1A7hww)R
RRRRRRRRRb0Fs5RR
RRRRRRRRRRRRRTRRRF:Rk#0R0D8_FOoHRR;
RRRRRRRRRRRRRBRRRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRR7RRRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRR)RRRH:RM#RR0D8_FOoHRR
RRRRRRRRRRRRRR
2;CRM8ObFlFMMC0
;
ObFlFMMC0AR1_w7whR1
RRRRRRRRRsbF0
5RRRRRRRRRRRRRRRRRTRR:FRk0#_08DHFoO
R;RRRRRRRRRRRRRRRRBRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRR7RR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRR1RR:HRMR#_08DHFoORR
RRRRRRRRRRRRR;R2
8CMRlOFbCFMM
0;
lOFbCFMM10RAw_7w
h RRRRRRRRRFRbsR05
RRRRRRRRRRRRRRRR:TRR0FkR8#0_oDFH;OR
RRRRRRRRRRRRRRRR:BRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRR: RRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRR:7RRRHMR8#0_oDFH
ORRRRRRRRRRRRRR2RR;M
C8FROlMbFC;M0
F
OlMbFCRM017A_w wh1R)
RRRRRRRRRsbF0
5RRRRRRRRRRRRRRRRRTRR:FRk0#_08DHFoO
R;RRRRRRRRRRRRRRRRBRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRR RR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRR7RR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRR)RR:HRMR#_08DHFoORR
RRRRRRRRRRRRR;R2
8CMRlOFbCFMM
0;
lOFbCFMM10RAw_7w1h 1R
RRRRRRRRRb0Fs5RR
RRRRRRRRRRRRRTRRRF:Rk#0R0D8_FOoHRR;
RRRRRRRRRRRRRBRRRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRR RRRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRR7RRRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRR1RRRH:RM#RR0D8_FOoHRR
RRRRRRRRRRRRRR
2;CRM8ObFlFMMC0
;
ObFlFMMC0AR1_w7wh
 )RRRRRRRRRFRbsR05
RRRRRRRRRRRRRRRR:TRR0FkR8#0_oDFH;OR
RRRRRRRRRRRRRRRR:BRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRR: RRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRR:7RRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRR:)RRRHMR8#0_oDFH
ORRRRRRRRRRRRRR2RR;M
C8FROlMbFC;M0
F
OlMbFCRM017A_w wh1R
RRRRRRRRRb0Fs5RR
RRRRRRRRRRRRRTRRRF:Rk#0R0D8_FOoHRR;
RRRRRRRRRRRRRBRRRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRR RRRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRR7RRRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRR1RRRH:RM#RR0D8_FOoHRR
RRRRRRRRRRRRRR
2;CRM8ObFlFMMC0
;
ObFlFMMC0AR1_v)qccj_iR
RRRRRRRRRoCCMsRHO5)RWQ_a v m7RH:RMo0CC:sR=;Rj
RRRRRRRRRRRRRRRRRRRRq) 7m_v7: RR0HMCsoCRR:=jR;
RRRRRRRRRRRRRRRRRQRRh_QajRR:L_H0P0COFRs5.R66RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRRRRRQQhaR_4:HRL0C_POs0F56R.68RRF0IMF2RjR
;RRRRRRRRRRRRRRRRRRRRRQahQ_:.RR0LH_OPC05FsR6.6RFR8IFM0RRj2;RR
RRRRRRRRRRRRRRRRRQRRh_QadRR:L_H0P0COFRs5.R66RI8FMR0Fj;2RRR
RRRRRRRRRRRRRRRRRRhRQQca_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2RR;
RRRRRRRRRRRRRRRRRRRRQQhaR_6:HRL0C_POs0F56R.68RRF0IMF2RjRR;
RRRRRRRRRRRRRRRRRQRRh_QanRR:L_H0P0COFRs5.R66RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRRRRRQQhaR_(:HRL0C_POs0F56R.68RRF0IMF2RjRR;
RRRRRRRRRRRRRRRRRQRRh_QaURR:L_H0P0COFRs5.R66RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRRRRRQQhaR_g:HRL0C_POs0F56R.68RRF0IMF2RjRR;
RRRRRRRRRRRRRRRRRQRRh_QaqRR:L_H0P0COFRs5.R66RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRRRRRQQhaR_A:HRL0C_POs0F56R.68RRF0IMF2RjRR;
RRRRRRRRRRRRRRRRRQRRh_QaBRR:L_H0P0COFRs5.R66RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRRRRRQQhaR_7:HRL0C_POs0F56R.68RRF0IMF2RjRR;
RRRRRRRRRRRRRRRRRQRRh_Qa RR:L_H0P0COFRs5.R66RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRRRRRQQhaR_w:HRL0C_POs0F56R.68RRF0IMF2RjRR
RRRRRRRRRRRRRRRRR2
R;RRRRRRRRRFRbsR05
RRRRRRRRRRRRRRRRq)7a:qRR0FkR8#0_oDFHPO_CFO0s45R68RRF0IMF2RjRR;
RRRRRRRRRRRRR)RRBRpi:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRBR)pRi :MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRR R)RRRR:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRqR)7R7):MRHR0R#8F_Do_HOP0COFRs54RjR8MFI0jFR2
R;RRRRRRRRRRRRRRRRWiBpRRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRRWiBp RR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRRWR RRRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRRW7q7)RR:HRMR#_08DHFoOC_POs0F5jR4RFR8IFM0RRj2;R
RRRRRRRRRRRRRRqRv1RiR:MRHR0R#8F_Do_HOP0COFRs54R6R8MFI0jFR2
R;RRRRRRRRRRRRRRRRWa7qqRR:HRMR#_08DHFoOC_POs0F56R4RFR8IFM0R
j2RRRRRRRRRRRRR2RR;M
C8FROlMbFC;M0
O

FFlbM0CMR_1A)cqvji_chR)
RRRRRRRRRMoCCOsHRW5R) Qa_7vm RR:HCM0oRCs:j=R;R
RRRRRRRRRRRRRRRRRR R)qv7_mR7 :MRH0CCos=R:R
j;RRRRRRRRRRRRRRRRRRRRQahQ_:jRR0LH_OPC05FsR6.6RFR8IFM0RRj2;R
RRRRRRRRRRRRRRRRRRhRQQ4a_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2RR;
RRRRRRRRRRRRRRRRRRRRQQhaR_.:HRL0C_POs0F56R.68RRF0IMF2RjR
;RRRRRRRRRRRRRRRRRRRRRQahQ_:dRR0LH_OPC05FsR6.6RFR8IFM0RRj2;RR
RRRRRRRRRRRRRRRRRQRRh_QacRR:L_H0P0COFRs5.R66RI8FMR0Fj;2RRR
RRRRRRRRRRRRRRRRRRhRQQ6a_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2
R;RRRRRRRRRRRRRRRRRRRRQahQ_:nRR0LH_OPC05FsR6.6RFR8IFM0RRj2;R
RRRRRRRRRRRRRRRRRRhRQQ(a_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2
R;RRRRRRRRRRRRRRRRRRRRQahQ_:URR0LH_OPC05FsR6.6RFR8IFM0RRj2;R
RRRRRRRRRRRRRRRRRRhRQQga_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2
R;RRRRRRRRRRRRRRRRRRRRQahQ_:qRR0LH_OPC05FsR6.6RFR8IFM0RRj2;R
RRRRRRRRRRRRRRRRRRhRQQAa_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2
R;RRRRRRRRRRRRRRRRRRRRQahQ_:BRR0LH_OPC05FsR6.6RFR8IFM0RRj2;R
RRRRRRRRRRRRRRRRRRhRQQ7a_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2
R;RRRRRRRRRRRRRRRRRRRRQahQ_: RR0LH_OPC05FsR6.6RFR8IFM0RRj2;R
RRRRRRRRRRRRRRRRRRhRQQwa_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2RR
RRRRRRRRRRRRRRRRR;2R
RRRRRRRRbRRF5s0RR
RRRRRRRRRRRRRR7R)qRaq:kRF00R#8F_Do_HOP0COFRs54R6R8MFI0jFR2
R;RRRRRRRRRRRRRRRR)iBphRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRR)iBp RR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRR)R RRRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRR)7q7)RR:HRMR#_08DHFoOC_POs0F5jR4RFR8IFM0RRj2;R
RRRRRRRRRRRRRRBRWpRiR:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRBRWpRi :MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRR RWRRRR:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRqRW7R7):MRHR0R#8F_Do_HOP0COFRs54RjR8MFI0jFR2
R;RRRRRRRRRRRRRRRRviq1RRR:HRMR#_08DHFoOC_POs0F56R4RFR8IFM0RRj2;R
RRRRRRRRRRRRRR7RWqRaq:MRHR0R#8F_Do_HOP0COFRs54R6R8MFI0jFR2R
RRRRRRRRRRRRRR
2;CRM8ObFlFMMC0
;

lOFbCFMM10RAq_)v_cjcWih
RRRRRRRRoRRCsMCH5ORRQW)av _mR7 :MRH0CCos=R:R
j;RRRRRRRRRRRRRRRRRRRR)7 q_7vm RR:HCM0oRCs:j=R;R
RRRRRRRRRRRRRRRRRRhRQQja_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2
R;RRRRRRRRRRRRRRRRRRRRQahQ_:4RR0LH_OPC05FsR6.6RFR8IFM0RRj2;RR
RRRRRRRRRRRRRRRRRQRRh_Qa.RR:L_H0P0COFRs5.R66RI8FMR0Fj;2RRR
RRRRRRRRRRRRRRRRRRhRQQda_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2RR;
RRRRRRRRRRRRRRRRRRRRQQhaR_c:HRL0C_POs0F56R.68RRF0IMF2RjR
;RRRRRRRRRRRRRRRRRRRRRQahQ_:6RR0LH_OPC05FsR6.6RFR8IFM0RRj2;R
RRRRRRRRRRRRRRRRRRhRQQna_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2
R;RRRRRRRRRRRRRRRRRRRRQahQ_:(RR0LH_OPC05FsR6.6RFR8IFM0RRj2;R
RRRRRRRRRRRRRRRRRRhRQQUa_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2
R;RRRRRRRRRRRRRRRRRRRRQahQ_:gRR0LH_OPC05FsR6.6RFR8IFM0RRj2;R
RRRRRRRRRRRRRRRRRRhRQQqa_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2
R;RRRRRRRRRRRRRRRRRRRRQahQ_:ARR0LH_OPC05FsR6.6RFR8IFM0RRj2;R
RRRRRRRRRRRRRRRRRRhRQQBa_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2
R;RRRRRRRRRRRRRRRRRRRRQahQ_:7RR0LH_OPC05FsR6.6RFR8IFM0RRj2;R
RRRRRRRRRRRRRRRRRRhRQQ a_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2
R;RRRRRRRRRRRRRRRRRRRRQahQ_:wRR0LH_OPC05FsR6.6RFR8IFM0RRj2
RRRRRRRRRRRRRRRR2RRRR;
RRRRRRRRRsbF0
5RRRRRRRRRRRRRRRRR)a7qqRR:FRk0#_08DHFoOC_POs0F56R4RFR8IFM0RRj2;R
RRRRRRRRRRRRRRBR)p:iRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRp)Bi: RRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRR) R:RRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRR7)q7:)RRRHMR8#0_oDFHPO_CFO0s45Rj8RRF0IMF2RjRR;
RRRRRRRRRRRRRWRRBhpiRRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRRWiBp RR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRRWR RRRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRRW7q7)RR:HRMR#_08DHFoOC_POs0F5jR4RFR8IFM0RRj2;R
RRRRRRRRRRRRRRqRv1RiR:MRHR0R#8F_Do_HOP0COFRs54R6R8MFI0jFR2
R;RRRRRRRRRRRRRRRRWa7qqRR:HRMR#_08DHFoOC_POs0F56R4RFR8IFM0R
j2RRRRRRRRRRRRR2RR;M
C8FROlMbFC;M0
O

FFlbM0CMR_1A)cqvji_chW)h
RRRRRRRRoRRCsMCH5ORRQW)av _mR7 :MRH0CCos=R:R
j;RRRRRRRRRRRRRRRRRRRR)7 q_7vm RR:HCM0oRCs:j=R;R
RRRRRRRRRRRRRRRRRRhRQQja_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2
R;RRRRRRRRRRRRRRRRRRRRQahQ_:4RR0LH_OPC05FsR6.6RFR8IFM0RRj2;RR
RRRRRRRRRRRRRRRRRQRRh_Qa.RR:L_H0P0COFRs5.R66RI8FMR0Fj;2RRR
RRRRRRRRRRRRRRRRRRhRQQda_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2RR;
RRRRRRRRRRRRRRRRRRRRQQhaR_c:HRL0C_POs0F56R.68RRF0IMF2RjR
;RRRRRRRRRRRRRRRRRRRRRQahQ_:6RR0LH_OPC05FsR6.6RFR8IFM0RRj2;R
RRRRRRRRRRRRRRRRRRhRQQna_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2
R;RRRRRRRRRRRRRRRRRRRRQahQ_:(RR0LH_OPC05FsR6.6RFR8IFM0RRj2;R
RRRRRRRRRRRRRRRRRRhRQQUa_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2
R;RRRRRRRRRRRRRRRRRRRRQahQ_:gRR0LH_OPC05FsR6.6RFR8IFM0RRj2;R
RRRRRRRRRRRRRRRRRRhRQQqa_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2
R;RRRRRRRRRRRRRRRRRRRRQahQ_:ARR0LH_OPC05FsR6.6RFR8IFM0RRj2;R
RRRRRRRRRRRRRRRRRRhRQQBa_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2
R;RRRRRRRRRRRRRRRRRRRRQahQ_:7RR0LH_OPC05FsR6.6RFR8IFM0RRj2;R
RRRRRRRRRRRRRRRRRRhRQQ a_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2
R;RRRRRRRRRRRRRRRRRRRRQahQ_:wRR0LH_OPC05FsR6.6RFR8IFM0RRj2
RRRRRRRRRRRRRRRR2RRRR;
RRRRRRRRRsbF0
5RRRRRRRRRRRRRRRRR)a7qqRR:FRk0#_08DHFoOC_POs0F56R4RFR8IFM0RRj2;R
RRRRRRRRRRRRRRBR)pRih:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRBR)pRi :MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRR R)RRRR:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRqR)7R7):MRHR0R#8F_Do_HOP0COFRs54RjR8MFI0jFR2
R;RRRRRRRRRRRRRRRRWiBph:RRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRpWBi: RRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRRW R:RRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRR7Wq7:)RRRHMR8#0_oDFHPO_CFO0s45Rj8RRF0IMF2RjRR;
RRRRRRRRRRRRRvRRqR1iRH:RM#RR0D8_FOoH_OPC05FsRR46RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRqW7a:qRRRHMR8#0_oDFHPO_CFO0s45R68RRF0IMF2Rj
RRRRRRRRRRRRRRR2C;
MO8RFFlbM0CM;O

FFlbM0CMR_1A).qv64nGnR
RRRRRRRRRoCCMsRHO5hRQQja_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2
R;RRRRRRRRRRRRRRRRRRRRQahQ_:4RR0LH_OPC05FsR6.6RFR8IFM0RRj2;RR
RRRRRRRRRRRRRRRRRQRRh_Qa.RR:L_H0P0COFRs5.R66RI8FMR0Fj;2RRR
RRRRRRRRRRRRRRRRRRhRQQda_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2RR;
RRRRRRRRRRRRRRRRRRRRQQhaR_c:HRL0C_POs0F56R.68RRF0IMF2RjR
;RRRRRRRRRRRRRRRRRRRRRQahQ_:6RR0LH_OPC05FsR6.6RFR8IFM0RRj2;R
RRRRRRRRRRRRRRRRRRhRQQna_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2
R;RRRRRRRRRRRRRRRRRRRRQahQ_:(RR0LH_OPC05FsR6.6RFR8IFM0RRj2;R
RRRRRRRRRRRRRRRRRRhRQQUa_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2
R;RRRRRRRRRRRRRRRRRRRRQahQ_:gRR0LH_OPC05FsR6.6RFR8IFM0RRj2;R
RRRRRRRRRRRRRRRRRRhRQQqa_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2
R;RRRRRRRRRRRRRRRRRRRRQahQ_:ARR0LH_OPC05FsR6.6RFR8IFM0RRj2;R
RRRRRRRRRRRRRRRRRRhRQQBa_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2
R;RRRRRRRRRRRRRRRRRRRRQahQ_:7RR0LH_OPC05FsR6.6RFR8IFM0RRj2;R
RRRRRRRRRRRRRRRRRRhRQQ a_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2
R;RRRRRRRRRRRRRRRRRRRRQahQ_:wRR0LH_OPC05FsR6.6RFR8IFM0RRj2
RRRRRRRRRRRRRRRR2RRRR;
RRRRRRRRRsbF0
5RRRRRRRRRRRRRRRRR)a7qqRR:FRk0#_08DHFoOC_POs0F56R4RFR8IFM0RRj2;R
RRRRRRRRRRRRRRBR)p:iRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRp)Bi: RRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRR) R:RRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRR7)q7:)RRRHMR8#0_oDFHPO_CFO0s(5RRFR8IFM0RRj2;R
RRRRRRRRRRRRRRBRWpRiR:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRBRWpRi :MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRR RWRRRR:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRqRW7R7):MRHR0R#8F_Do_HOP0COFRs5(8RRF0IMF2RjRR;
RRRRRRRRRRRRRvRRqR1iRH:RM#RR0D8_FOoH_OPC05FsRR46RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRqW7a:qRRRHMR8#0_oDFHPO_CFO0s45R68RRF0IMF2Rj
RRRRRRRRRRRRRRR2C;
MO8RFFlbM0CM;O

FFlbM0CMR_1A).qv64nGn
h)RRRRRRRRRCRoMHCsORR5QahQ_:jRR0LH_OPC05FsR6.6RFR8IFM0RRj2;R
RRRRRRRRRRRRRRRRRRhRQQ4a_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2RR;
RRRRRRRRRRRRRRRRRRRRQQhaR_.:HRL0C_POs0F56R.68RRF0IMF2RjR
;RRRRRRRRRRRRRRRRRRRRRQahQ_:dRR0LH_OPC05FsR6.6RFR8IFM0RRj2;RR
RRRRRRRRRRRRRRRRRQRRh_QacRR:L_H0P0COFRs5.R66RI8FMR0Fj;2RRR
RRRRRRRRRRRRRRRRRRhRQQ6a_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2
R;RRRRRRRRRRRRRRRRRRRRQahQ_:nRR0LH_OPC05FsR6.6RFR8IFM0RRj2;R
RRRRRRRRRRRRRRRRRRhRQQ(a_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2
R;RRRRRRRRRRRRRRRRRRRRQahQ_:URR0LH_OPC05FsR6.6RFR8IFM0RRj2;R
RRRRRRRRRRRRRRRRRRhRQQga_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2
R;RRRRRRRRRRRRRRRRRRRRQahQ_:qRR0LH_OPC05FsR6.6RFR8IFM0RRj2;R
RRRRRRRRRRRRRRRRRRhRQQAa_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2
R;RRRRRRRRRRRRRRRRRRRRQahQ_:BRR0LH_OPC05FsR6.6RFR8IFM0RRj2;R
RRRRRRRRRRRRRRRRRRhRQQ7a_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2
R;RRRRRRRRRRRRRRRRRRRRQahQ_: RR0LH_OPC05FsR6.6RFR8IFM0RRj2;R
RRRRRRRRRRRRRRRRRRhRQQwa_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2RR
RRRRRRRRRRRRRRRRR;2R
RRRRRRRRbRRF5s0RR
RRRRRRRRRRRRRR7R)qRaq:kRF00R#8F_Do_HOP0COFRs54R6R8MFI0jFR2
R;RRRRRRRRRRRRRRRR)iBph:RRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRp)Bi: RRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRR) R:RRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRR7)q7:)RRRHMR8#0_oDFHPO_CFO0s(5RRFR8IFM0RRj2;R
RRRRRRRRRRRRRRBRWp:iRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRpWBi: RRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRRW R:RRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRR7Wq7:)RRRHMR8#0_oDFHPO_CFO0s(5RRFR8IFM0RRj2;R
RRRRRRRRRRRRRRqRv1RiR:MRHR0R#8F_Do_HOP0COFRs54R6R8MFI0jFR2
R;RRRRRRRRRRRRRRRRWa7qqRR:HRMR#_08DHFoOC_POs0F56R4RFR8IFM0R
j2RRRRRRRRRRRRR2RR;M
C8FROlMbFC;M0
F
OlMbFCRM01)A_q6v.nnG4hRW
RRRRRRRRRMoCCOsHRQ5Rh_QajRR:L_H0P0COFRs5.R66RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRRRRRQQhaR_4:HRL0C_POs0F56R.68RRF0IMF2RjR
;RRRRRRRRRRRRRRRRRRRRRQahQ_:.RR0LH_OPC05FsR6.6RFR8IFM0RRj2;RR
RRRRRRRRRRRRRRRRRQRRh_QadRR:L_H0P0COFRs5.R66RI8FMR0Fj;2RRR
RRRRRRRRRRRRRRRRRRhRQQca_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2RR;
RRRRRRRRRRRRRRRRRRRRQQhaR_6:HRL0C_POs0F56R.68RRF0IMF2RjRR;
RRRRRRRRRRRRRRRRRQRRh_QanRR:L_H0P0COFRs5.R66RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRRRRRQQhaR_(:HRL0C_POs0F56R.68RRF0IMF2RjRR;
RRRRRRRRRRRRRRRRRQRRh_QaURR:L_H0P0COFRs5.R66RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRRRRRQQhaR_g:HRL0C_POs0F56R.68RRF0IMF2RjRR;
RRRRRRRRRRRRRRRRRQRRh_QaqRR:L_H0P0COFRs5.R66RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRRRRRQQhaR_A:HRL0C_POs0F56R.68RRF0IMF2RjRR;
RRRRRRRRRRRRRRRRRQRRh_QaBRR:L_H0P0COFRs5.R66RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRRRRRQQhaR_7:HRL0C_POs0F56R.68RRF0IMF2RjRR;
RRRRRRRRRRRRRRRRRQRRh_Qa RR:L_H0P0COFRs5.R66RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRRRRRQQhaR_w:HRL0C_POs0F56R.68RRF0IMF2RjRR
RRRRRRRRRRRRRRRRR2
R;RRRRRRRRRFRbsR05
RRRRRRRRRRRRRRRRq)7a:qRR0FkR8#0_oDFHPO_CFO0s45R68RRF0IMF2RjRR;
RRRRRRRRRRRRR)RRBRpi:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRBR)pRi :MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRR R)RRRR:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRqR)7R7):MRHR0R#8F_Do_HOP0COFRs5(8RRF0IMF2RjRR;
RRRRRRRRRRRRRWRRBhpiRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRRWRRB piRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRRWRR RRRRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRRWRRq)77RH:RM#RR0D8_FOoH_OPC05FsRR(R8MFI0jFR2
R;RRRRRRRRRRRRRRRRviq1RRR:HRMR#_08DHFoOC_POs0F56R4RFR8IFM0RRj2;R
RRRRRRRRRRRRRR7RWqRaq:MRHR0R#8F_Do_HOP0COFRs54R6R8MFI0jFR2R
RRRRRRRRRRRRRR
2;CRM8ObFlFMMC0
;
ObFlFMMC0AR1_v)q.G6n4)nhhRW
RRRRRRRRRMoCCOsHRQ5Rh_QajRR:L_H0P0COFRs5.R66RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRRRRRQQhaR_4:HRL0C_POs0F56R.68RRF0IMF2RjR
;RRRRRRRRRRRRRRRRRRRRRQahQ_:.RR0LH_OPC05FsR6.6RFR8IFM0RRj2;RR
RRRRRRRRRRRRRRRRRQRRh_QadRR:L_H0P0COFRs5.R66RI8FMR0Fj;2RRR
RRRRRRRRRRRRRRRRRRhRQQca_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2RR;
RRRRRRRRRRRRRRRRRRRRQQhaR_6:HRL0C_POs0F56R.68RRF0IMF2RjRR;
RRRRRRRRRRRRRRRRRQRRh_QanRR:L_H0P0COFRs5.R66RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRRRRRQQhaR_(:HRL0C_POs0F56R.68RRF0IMF2RjRR;
RRRRRRRRRRRRRRRRRQRRh_QaURR:L_H0P0COFRs5.R66RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRRRRRQQhaR_g:HRL0C_POs0F56R.68RRF0IMF2RjRR;
RRRRRRRRRRRRRRRRRQRRh_QaqRR:L_H0P0COFRs5.R66RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRRRRRQQhaR_A:HRL0C_POs0F56R.68RRF0IMF2RjRR;
RRRRRRRRRRRRRRRRRQRRh_QaBRR:L_H0P0COFRs5.R66RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRRRRRQQhaR_7:HRL0C_POs0F56R.68RRF0IMF2RjRR;
RRRRRRRRRRRRRRRRRQRRh_Qa RR:L_H0P0COFRs5.R66RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRRRRRQQhaR_w:HRL0C_POs0F56R.68RRF0IMF2RjRR
RRRRRRRRRRRRRRRRR2
R;RRRRRRRRRFRbsR05
RRRRRRRRRRRRRRRRq)7a:qRR0FkR8#0_oDFHPO_CFO0s45R68RRF0IMF2RjRR;
RRRRRRRRRRRRR)RRBhpiRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRR)RRB piRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRR)RR RRRRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRR)RRq)77RH:RM#RR0D8_FOoH_OPC05FsRR(R8MFI0jFR2
R;RRRRRRRRRRRRRRRRWiBph:RRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRpWBi: RRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRRW R:RRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRR7Wq7:)RRRHMR8#0_oDFHPO_CFO0s(5RRFR8IFM0RRj2;R
RRRRRRRRRRRRRRqRv1RiR:MRHR0R#8F_Do_HOP0COFRs54R6R8MFI0jFR2
R;RRRRRRRRRRRRRRRRWa7qqRR:HRMR#_08DHFoOC_POs0F56R4RFR8IFM0R
j2RRRRRRRRRRRRR2RR;M
C8FROlMbFC;M0
O

FFlbM0CMR_1A)6qv4U.G
RRRRRRRRoRRCsMCH5ORRQQhaR_j:HRL0C_POs0F56R.68RRF0IMF2RjRR;
RRRRRRRRRRRRRRRRRQRRh_Qa4RR:L_H0P0COFRs5.R66RI8FMR0Fj;2RRR
RRRRRRRRRRRRRRRRRRhRQQ.a_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2RR;
RRRRRRRRRRRRRRRRRRRRQQhaR_d:HRL0C_POs0F56R.68RRF0IMF2RjR
;RRRRRRRRRRRRRRRRRRRRRQahQ_:cRR0LH_OPC05FsR6.6RFR8IFM0RRj2;RR
RRRRRRRRRRRRRRRRRQRRh_Qa6RR:L_H0P0COFRs5.R66RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRRRRRQQhaR_n:HRL0C_POs0F56R.68RRF0IMF2RjRR;
RRRRRRRRRRRRRRRRRQRRh_Qa(RR:L_H0P0COFRs5.R66RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRRRRRQQhaR_U:HRL0C_POs0F56R.68RRF0IMF2RjRR;
RRRRRRRRRRRRRRRRRQRRh_QagRR:L_H0P0COFRs5.R66RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRRRRRQQhaR_q:HRL0C_POs0F56R.68RRF0IMF2RjRR;
RRRRRRRRRRRRRRRRRQRRh_QaARR:L_H0P0COFRs5.R66RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRRRRRQQhaR_B:HRL0C_POs0F56R.68RRF0IMF2RjRR;
RRRRRRRRRRRRRRRRRQRRh_Qa7RR:L_H0P0COFRs5.R66RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRRRRRQQhaR_ :HRL0C_POs0F56R.68RRF0IMF2RjRR;
RRRRRRRRRRRRRRRRRQRRh_QawRR:L_H0P0COFRs5.R66RI8FMR0Fj
2RRRRRRRRRRRRRRRRRRRR2;R
RRRRRRRRRb0Fs5RR
RRRRRRRRRRRRR)RR7qqaRF:Rk#0R0D8_FOoH_OPC05FsRR(R8MFI0jFR2
R;RRRRRRRRRRRRRRRR)iBpRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRR)RRB piRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRR)RR RRRRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRR)RRq)77RH:RM#RR0D8_FOoH_OPC05FsRRUR8MFI0jFR2
R;RRRRRRRRRRRRRRRRWiBpRRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRRWiBp RR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRRWR RRRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRRW7q7)RR:HRMR#_08DHFoOC_POs0F5RRURI8FMR0Fj;2R
RRRRRRRRRRRRRRRRqW7a:qRRRHMR8#0_oDFHPO_CFO0s(5RRFR8IFM0R
j2RRRRRRRRRRRRR2RR;M
C8FROlMbFC;M0
O

FFlbM0CMR_1A)6qv4U.GhR)
RRRRRRRRRMoCCOsHRQ5Rh_QajRR:L_H0P0COFRs5.R66RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRRRRRQQhaR_4:HRL0C_POs0F56R.68RRF0IMF2RjR
;RRRRRRRRRRRRRRRRRRRRRQahQ_:.RR0LH_OPC05FsR6.6RFR8IFM0RRj2;RR
RRRRRRRRRRRRRRRRRQRRh_QadRR:L_H0P0COFRs5.R66RI8FMR0Fj;2RRR
RRRRRRRRRRRRRRRRRRhRQQca_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2RR;
RRRRRRRRRRRRRRRRRRRRQQhaR_6:HRL0C_POs0F56R.68RRF0IMF2RjRR;
RRRRRRRRRRRRRRRRRQRRh_QanRR:L_H0P0COFRs5.R66RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRRRRRQQhaR_(:HRL0C_POs0F56R.68RRF0IMF2RjRR;
RRRRRRRRRRRRRRRRRQRRh_QaURR:L_H0P0COFRs5.R66RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRRRRRQQhaR_g:HRL0C_POs0F56R.68RRF0IMF2RjRR;
RRRRRRRRRRRRRRRRRQRRh_QaqRR:L_H0P0COFRs5.R66RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRRRRRQQhaR_A:HRL0C_POs0F56R.68RRF0IMF2RjRR;
RRRRRRRRRRRRRRRRRQRRh_QaBRR:L_H0P0COFRs5.R66RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRRRRRQQhaR_7:HRL0C_POs0F56R.68RRF0IMF2RjRR;
RRRRRRRRRRRRRRRRRQRRh_Qa RR:L_H0P0COFRs5.R66RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRRRRRQQhaR_w:HRL0C_POs0F56R.68RRF0IMF2RjRR
RRRRRRRRRRRRRRRRR2
R;RRRRRRRRRFRbsR05
RRRRRRRRRRRRRRRRq)7a:qRR0FkR8#0_oDFHPO_CFO0s(5RRFR8IFM0RRj2;R
RRRRRRRRRRRRRRBR)pRih:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRBR)pRi :MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRR R)RRRR:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRqR)7R7):MRHR0R#8F_Do_HOP0COFRs5U8RRF0IMF2RjRR;
RRRRRRRRRRRRRWRRBRpiRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRRWRRB piRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRRWRR RRRRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRRWRRq)77RH:RM#RR0D8_FOoH_OPC05FsRRUR8MFI0jFR2
R;RRRRRRRRRRRRRRRRWa7qqRR:HRMR#_08DHFoOC_POs0F5RR(RI8FMR0FjR2
RRRRRRRRRRRRR;R2
8CMRlOFbCFMM
0;
lOFbCFMM10RAq_)v.64GWUh
RRRRRRRRoRRCsMCH5ORRQQhaR_j:HRL0C_POs0F56R.68RRF0IMF2RjRR;
RRRRRRRRRRRRRRRRRQRRh_Qa4RR:L_H0P0COFRs5.R66RI8FMR0Fj;2RRR
RRRRRRRRRRRRRRRRRRhRQQ.a_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2RR;
RRRRRRRRRRRRRRRRRRRRQQhaR_d:HRL0C_POs0F56R.68RRF0IMF2RjR
;RRRRRRRRRRRRRRRRRRRRRQahQ_:cRR0LH_OPC05FsR6.6RFR8IFM0RRj2;RR
RRRRRRRRRRRRRRRRRQRRh_Qa6RR:L_H0P0COFRs5.R66RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRRRRRQQhaR_n:HRL0C_POs0F56R.68RRF0IMF2RjRR;
RRRRRRRRRRRRRRRRRQRRh_Qa(RR:L_H0P0COFRs5.R66RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRRRRRQQhaR_U:HRL0C_POs0F56R.68RRF0IMF2RjRR;
RRRRRRRRRRRRRRRRRQRRh_QagRR:L_H0P0COFRs5.R66RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRRRRRQQhaR_q:HRL0C_POs0F56R.68RRF0IMF2RjRR;
RRRRRRRRRRRRRRRRRQRRh_QaARR:L_H0P0COFRs5.R66RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRRRRRQQhaR_B:HRL0C_POs0F56R.68RRF0IMF2RjRR;
RRRRRRRRRRRRRRRRRQRRh_Qa7RR:L_H0P0COFRs5.R66RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRRRRRQQhaR_ :HRL0C_POs0F56R.68RRF0IMF2RjRR;
RRRRRRRRRRRRRRRRRQRRh_QawRR:L_H0P0COFRs5.R66RI8FMR0Fj
2RRRRRRRRRRRRRRRRRRRR2;R
RRRRRRRRRb0Fs5RR
RRRRRRRRRRRRR)RR7qqaRF:Rk#0R0D8_FOoH_OPC05FsRR(R8MFI0jFR2
R;RRRRRRRRRRRRRRRR)iBpRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRR)RRB piRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRR)RR RRRRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRR)RRq)77RH:RM#RR0D8_FOoH_OPC05FsRRUR8MFI0jFR2
R;RRRRRRRRRRRRRRRRWiBph:RRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRpWBi: RRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRRW R:RRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRR7Wq7:)RRRHMR8#0_oDFHPO_CFO0sU5RRFR8IFM0RRj2;R
RRRRRRRRRRRRRR7RWqRaq:MRHR0R#8F_Do_HOP0COFRs5(8RRF0IMF2Rj
RRRRRRRRRRRRRRR2C;
MO8RFFlbM0CM;O

FFlbM0CMR_1A)6qv4U.GhW)h
RRRRRRRRoRRCsMCH5ORRQQhaR_j:HRL0C_POs0F56R.68RRF0IMF2RjRR;
RRRRRRRRRRRRRRRRRQRRh_Qa4RR:L_H0P0COFRs5.R66RI8FMR0Fj;2RRR
RRRRRRRRRRRRRRRRRRhRQQ.a_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2RR;
RRRRRRRRRRRRRRRRRRRRQQhaR_d:HRL0C_POs0F56R.68RRF0IMF2RjR
;RRRRRRRRRRRRRRRRRRRRRQahQ_:cRR0LH_OPC05FsR6.6RFR8IFM0RRj2;RR
RRRRRRRRRRRRRRRRRQRRh_Qa6RR:L_H0P0COFRs5.R66RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRRRRRQQhaR_n:HRL0C_POs0F56R.68RRF0IMF2RjRR;
RRRRRRRRRRRRRRRRRQRRh_Qa(RR:L_H0P0COFRs5.R66RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRRRRRQQhaR_U:HRL0C_POs0F56R.68RRF0IMF2RjRR;
RRRRRRRRRRRRRRRRRQRRh_QagRR:L_H0P0COFRs5.R66RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRRRRRQQhaR_q:HRL0C_POs0F56R.68RRF0IMF2RjRR;
RRRRRRRRRRRRRRRRRQRRh_QaARR:L_H0P0COFRs5.R66RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRRRRRQQhaR_B:HRL0C_POs0F56R.68RRF0IMF2RjRR;
RRRRRRRRRRRRRRRRRQRRh_Qa7RR:L_H0P0COFRs5.R66RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRRRRRQQhaR_ :HRL0C_POs0F56R.68RRF0IMF2RjRR;
RRRRRRRRRRRRRRRRRQRRh_QawRR:L_H0P0COFRs5.R66RI8FMR0Fj
2RRRRRRRRRRRRRRRRRRRR2;R
RRRRRRRRRb0Fs5RR
RRRRRRRRRRRRR)RR7qqaRF:Rk#0R0D8_FOoH_OPC05FsRR(R8MFI0jFR2
R;RRRRRRRRRRRRRRRR)iBphRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRR)iBp RR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRR)R RRRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRR)7q7)RR:HRMR#_08DHFoOC_POs0F5RRURI8FMR0Fj;2R
RRRRRRRRRRRRRRRRpWBiRhR:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRBRWpRi :MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRR RWRRRR:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRqRW7R7):MRHR0R#8F_Do_HOP0COFRs5U8RRF0IMF2RjRR;
RRRRRRRRRRRRRWRR7qqaRH:RM#RR0D8_FOoH_OPC05FsRR(R8MFI0jFR2R
RRRRRRRRRRRRRR
2;CRM8ObFlFMMC0
;

lOFbCFMM10RAq_)v.4jc
GcRRRRRRRRRCRoMHCsORR5QahQ_:jRR0LH_OPC05FsR6.6RFR8IFM0RRj2;R
RRRRRRRRRRRRRRRRRRhRQQ4a_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2RR;
RRRRRRRRRRRRRRRRRRRRQQhaR_.:HRL0C_POs0F56R.68RRF0IMF2RjR
;RRRRRRRRRRRRRRRRRRRRRQahQ_:dRR0LH_OPC05FsR6.6RFR8IFM0RRj2;RR
RRRRRRRRRRRRRRRRRQRRh_QacRR:L_H0P0COFRs5.R66RI8FMR0Fj;2RRR
RRRRRRRRRRRRRRRRRRhRQQ6a_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2
R;RRRRRRRRRRRRRRRRRRRRQahQ_:nRR0LH_OPC05FsR6.6RFR8IFM0RRj2;R
RRRRRRRRRRRRRRRRRRhRQQ(a_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2
R;RRRRRRRRRRRRRRRRRRRRQahQ_:URR0LH_OPC05FsR6.6RFR8IFM0RRj2;R
RRRRRRRRRRRRRRRRRRhRQQga_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2
R;RRRRRRRRRRRRRRRRRRRRQahQ_:qRR0LH_OPC05FsR6.6RFR8IFM0RRj2;R
RRRRRRRRRRRRRRRRRRhRQQAa_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2
R;RRRRRRRRRRRRRRRRRRRRQahQ_:BRR0LH_OPC05FsR6.6RFR8IFM0RRj2;R
RRRRRRRRRRRRRRRRRRhRQQ7a_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2
R;RRRRRRRRRRRRRRRRRRRRQahQ_: RR0LH_OPC05FsR6.6RFR8IFM0RRj2;R
RRRRRRRRRRRRRRRRRRhRQQwa_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2RR
RRRRRRRRRRRRRRRRR;2R
RRRRRRRRbRRF5s0RR
RRRRRRRRRRRRRR7R)qRaq:kRF00R#8F_Do_HOP0COFRs5d8RRF0IMF2RjRR;
RRRRRRRRRRRRR)RRBRpi:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRBR)pRi :MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRR R)RRRR:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRqR)7R7):MRHR0R#8F_Do_HOP0COFRs5g8RRF0IMF2RjRR;
RRRRRRRRRRRRRWRRBRpiRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRRWRRB piRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRRWRR RRRRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRRWRRq)77RH:RM#RR0D8_FOoH_OPC05FsRRgR8MFI0jFR2
R;RRRRRRRRRRRRRRRRWa7qqRR:HRMR#_08DHFoOC_POs0F5RRdRI8FMR0FjR2
RRRRRRRRRRRRR;R2
8CMRlOFbCFMM
0;
lOFbCFMM10RAq_)v.4jchGc)R
RRRRRRRRRoCCMsRHO5hRQQja_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2
R;RRRRRRRRRRRRRRRRRRRRQahQ_:4RR0LH_OPC05FsR6.6RFR8IFM0RRj2;RR
RRRRRRRRRRRRRRRRRQRRh_Qa.RR:L_H0P0COFRs5.R66RI8FMR0Fj;2RRR
RRRRRRRRRRRRRRRRRRhRQQda_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2RR;
RRRRRRRRRRRRRRRRRRRRQQhaR_c:HRL0C_POs0F56R.68RRF0IMF2RjR
;RRRRRRRRRRRRRRRRRRRRRQahQ_:6RR0LH_OPC05FsR6.6RFR8IFM0RRj2;R
RRRRRRRRRRRRRRRRRRhRQQna_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2
R;RRRRRRRRRRRRRRRRRRRRQahQ_:(RR0LH_OPC05FsR6.6RFR8IFM0RRj2;R
RRRRRRRRRRRRRRRRRRhRQQUa_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2
R;RRRRRRRRRRRRRRRRRRRRQahQ_:gRR0LH_OPC05FsR6.6RFR8IFM0RRj2;R
RRRRRRRRRRRRRRRRRRhRQQqa_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2
R;RRRRRRRRRRRRRRRRRRRRQahQ_:ARR0LH_OPC05FsR6.6RFR8IFM0RRj2;R
RRRRRRRRRRRRRRRRRRhRQQBa_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2
R;RRRRRRRRRRRRRRRRRRRRQahQ_:7RR0LH_OPC05FsR6.6RFR8IFM0RRj2;R
RRRRRRRRRRRRRRRRRRhRQQ a_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2
R;RRRRRRRRRRRRRRRRRRRRQahQ_:wRR0LH_OPC05FsR6.6RFR8IFM0RRj2
RRRRRRRRRRRRRRRR2RRRR;
RRRRRRRRRsbF0
5RRRRRRRRRRRRRRRRR)a7qqRR:FRk0#_08DHFoOC_POs0F5RRdRI8FMR0Fj;2R
RRRRRRRRRRRRRRRRp)Bi:hRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRp)Bi: RRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRR) R:RRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRR7)q7:)RRRHMR8#0_oDFHPO_CFO0sg5RRFR8IFM0RRj2;R
RRRRRRRRRRRRRRBRWpRiR:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRBRWpRi :MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRR RWRRRR:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRqRW7R7):MRHR0R#8F_Do_HOP0COFRs5g8RRF0IMF2RjRR;
RRRRRRRRRRRRRWRR7qqaRH:RM#RR0D8_FOoH_OPC05FsRRdR8MFI0jFR2R
RRRRRRRRRRRRRR
2;CRM8ObFlFMMC0
;
ObFlFMMC0AR1_v)q4cj.GWch
RRRRRRRRoRRCsMCH5ORRQQhaR_j:HRL0C_POs0F56R.68RRF0IMF2RjRR;
RRRRRRRRRRRRRRRRRQRRh_Qa4RR:L_H0P0COFRs5.R66RI8FMR0Fj;2RRR
RRRRRRRRRRRRRRRRRRhRQQ.a_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2RR;
RRRRRRRRRRRRRRRRRRRRQQhaR_d:HRL0C_POs0F56R.68RRF0IMF2RjR
;RRRRRRRRRRRRRRRRRRRRRQahQ_:cRR0LH_OPC05FsR6.6RFR8IFM0RRj2;RR
RRRRRRRRRRRRRRRRRQRRh_Qa6RR:L_H0P0COFRs5.R66RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRRRRRQQhaR_n:HRL0C_POs0F56R.68RRF0IMF2RjRR;
RRRRRRRRRRRRRRRRRQRRh_Qa(RR:L_H0P0COFRs5.R66RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRRRRRQQhaR_U:HRL0C_POs0F56R.68RRF0IMF2RjRR;
RRRRRRRRRRRRRRRRRQRRh_QagRR:L_H0P0COFRs5.R66RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRRRRRQQhaR_q:HRL0C_POs0F56R.68RRF0IMF2RjRR;
RRRRRRRRRRRRRRRRRQRRh_QaARR:L_H0P0COFRs5.R66RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRRRRRQQhaR_B:HRL0C_POs0F56R.68RRF0IMF2RjRR;
RRRRRRRRRRRRRRRRRQRRh_Qa7RR:L_H0P0COFRs5.R66RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRRRRRQQhaR_ :HRL0C_POs0F56R.68RRF0IMF2RjRR;
RRRRRRRRRRRRRRRRRQRRh_QawRR:L_H0P0COFRs5.R66RI8FMR0Fj
2RRRRRRRRRRRRRRRRRRRR2;R
RRRRRRRRRb0Fs5RR
RRRRRRRRRRRRR)RR7qqaRF:Rk#0R0D8_FOoH_OPC05FsRRdR8MFI0jFR2
R;RRRRRRRRRRRRRRRR)iBpRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRR)RRB piRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRR)RR RRRRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRR)RRq)77RH:RM#RR0D8_FOoH_OPC05FsRRgR8MFI0jFR2
R;RRRRRRRRRRRRRRRRWiBph:RRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRpWBi: RRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRRW R:RRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRR7Wq7:)RRRHMR8#0_oDFHPO_CFO0sg5RRFR8IFM0RRj2;R
RRRRRRRRRRRRRR7RWqRaq:MRHR0R#8F_Do_HOP0COFRs5d8RRF0IMF2Rj
RRRRRRRRRRRRRRR2C;
MO8RFFlbM0CM;O

FFlbM0CMR_1A)4qvjG.cchh)WR
RRRRRRRRRoCCMsRHO5hRQQja_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2
R;RRRRRRRRRRRRRRRRRRRRQahQ_:4RR0LH_OPC05FsR6.6RFR8IFM0RRj2;RR
RRRRRRRRRRRRRRRRRQRRh_Qa.RR:L_H0P0COFRs5.R66RI8FMR0Fj;2RRR
RRRRRRRRRRRRRRRRRRhRQQda_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2RR;
RRRRRRRRRRRRRRRRRRRRQQhaR_c:HRL0C_POs0F56R.68RRF0IMF2RjR
;RRRRRRRRRRRRRRRRRRRRRQahQ_:6RR0LH_OPC05FsR6.6RFR8IFM0RRj2;R
RRRRRRRRRRRRRRRRRRhRQQna_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2
R;RRRRRRRRRRRRRRRRRRRRQahQ_:(RR0LH_OPC05FsR6.6RFR8IFM0RRj2;R
RRRRRRRRRRRRRRRRRRhRQQUa_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2
R;RRRRRRRRRRRRRRRRRRRRQahQ_:gRR0LH_OPC05FsR6.6RFR8IFM0RRj2;R
RRRRRRRRRRRRRRRRRRhRQQqa_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2
R;RRRRRRRRRRRRRRRRRRRRQahQ_:ARR0LH_OPC05FsR6.6RFR8IFM0RRj2;R
RRRRRRRRRRRRRRRRRRhRQQBa_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2
R;RRRRRRRRRRRRRRRRRRRRQahQ_:7RR0LH_OPC05FsR6.6RFR8IFM0RRj2;R
RRRRRRRRRRRRRRRRRRhRQQ a_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2
R;RRRRRRRRRRRRRRRRRRRRQahQ_:wRR0LH_OPC05FsR6.6RFR8IFM0RRj2
RRRRRRRRRRRRRRRR2RRRR;
RRRRRRRRRsbF0
5RRRRRRRRRRRRRRRRR)a7qqRR:FRk0#_08DHFoOC_POs0F5RRdRI8FMR0Fj;2R
RRRRRRRRRRRRRRRRp)Bi:hRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRp)Bi: RRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRR) R:RRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRR7)q7:)RRRHMR8#0_oDFHPO_CFO0sg5RRFR8IFM0RRj2;R
RRRRRRRRRRRRRRBRWpRihRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRRWRRB piRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRRWRR RRRRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRRWRRq)77RH:RM#RR0D8_FOoH_OPC05FsRRgR8MFI0jFR2
R;RRRRRRRRRRRRRRRRWa7qqRR:HRMR#_08DHFoOC_POs0F5RRdRI8FMR0FjR2
RRRRRRRRRRRRR;R2
8CMRlOFbCFMM
0;
F
OlMbFCRM01)A_qjv.c.UG
RRRRRRRRoRRCsMCH5ORRQQhaR_j:HRL0C_POs0F56R.68RRF0IMF2RjRR;
RRRRRRRRRRRRRRRRRQRRh_Qa4RR:L_H0P0COFRs5.R66RI8FMR0Fj;2RRR
RRRRRRRRRRRRRRRRRRhRQQ.a_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2RR;
RRRRRRRRRRRRRRRRRRRRQQhaR_d:HRL0C_POs0F56R.68RRF0IMF2RjR
;RRRRRRRRRRRRRRRRRRRRRQahQ_:cRR0LH_OPC05FsR6.6RFR8IFM0RRj2;RR
RRRRRRRRRRRRRRRRRQRRh_Qa6RR:L_H0P0COFRs5.R66RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRRRRRQQhaR_n:HRL0C_POs0F56R.68RRF0IMF2RjRR;
RRRRRRRRRRRRRRRRRQRRh_Qa(RR:L_H0P0COFRs5.R66RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRRRRRQQhaR_U:HRL0C_POs0F56R.68RRF0IMF2RjRR;
RRRRRRRRRRRRRRRRRQRRh_QagRR:L_H0P0COFRs5.R66RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRRRRRQQhaR_q:HRL0C_POs0F56R.68RRF0IMF2RjRR;
RRRRRRRRRRRRRRRRRQRRh_QaARR:L_H0P0COFRs5.R66RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRRRRRQQhaR_B:HRL0C_POs0F56R.68RRF0IMF2RjRR;
RRRRRRRRRRRRRRRRRQRRh_Qa7RR:L_H0P0COFRs5.R66RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRRRRRQQhaR_ :HRL0C_POs0F56R.68RRF0IMF2RjRR;
RRRRRRRRRRRRRRRRRQRRh_QawRR:L_H0P0COFRs5.R66RI8FMR0Fj
2RRRRRRRRRRRRRRRRRRRR2;R
RRRRRRRRRb0Fs5RR
RRRRRRRRRRRRR)RR7qqaRF:Rk#0R0D8_FOoH_OPC05FsRR4R8MFI0jFR2
R;RRRRRRRRRRRRRRRR)iBpRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRR)RRB piRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRR)RR RRRRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRR)RRq)77RH:RM#RR0D8_FOoH_OPC05FsRR4jRI8FMR0Fj;2R
RRRRRRRRRRRRRRRRpWBi:RRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRpWBi: RRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRRW R:RRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRR7Wq7:)RRRHMR8#0_oDFHPO_CFO0s45Rj8RRF0IMF2RjRR;
RRRRRRRRRRRRRWRR7qqaRH:RM#RR0D8_FOoH_OPC05FsRR4R8MFI0jFR2R
RRRRRRRRRRRRRR
2;CRM8ObFlFMMC0
;
ObFlFMMC0AR1_v)q.UjcG).h
RRRRRRRRoRRCsMCH5ORRQQhaR_j:HRL0C_POs0F56R.68RRF0IMF2RjRR;
RRRRRRRRRRRRRRRRRQRRh_Qa4RR:L_H0P0COFRs5.R66RI8FMR0Fj;2RRR
RRRRRRRRRRRRRRRRRRhRQQ.a_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2RR;
RRRRRRRRRRRRRRRRRRRRQQhaR_d:HRL0C_POs0F56R.68RRF0IMF2RjR
;RRRRRRRRRRRRRRRRRRRRRQahQ_:cRR0LH_OPC05FsR6.6RFR8IFM0RRj2;RR
RRRRRRRRRRRRRRRRRQRRh_Qa6RR:L_H0P0COFRs5.R66RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRRRRRQQhaR_n:HRL0C_POs0F56R.68RRF0IMF2RjRR;
RRRRRRRRRRRRRRRRRQRRh_Qa(RR:L_H0P0COFRs5.R66RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRRRRRQQhaR_U:HRL0C_POs0F56R.68RRF0IMF2RjRR;
RRRRRRRRRRRRRRRRRQRRh_QagRR:L_H0P0COFRs5.R66RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRRRRRQQhaR_q:HRL0C_POs0F56R.68RRF0IMF2RjRR;
RRRRRRRRRRRRRRRRRQRRh_QaARR:L_H0P0COFRs5.R66RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRRRRRQQhaR_B:HRL0C_POs0F56R.68RRF0IMF2RjRR;
RRRRRRRRRRRRRRRRRQRRh_Qa7RR:L_H0P0COFRs5.R66RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRRRRRQQhaR_ :HRL0C_POs0F56R.68RRF0IMF2RjRR;
RRRRRRRRRRRRRRRRRQRRh_QawRR:L_H0P0COFRs5.R66RI8FMR0Fj
2RRRRRRRRRRRRRRRRRRRR2;R
RRRRRRRRRb0Fs5RR
RRRRRRRRRRRRR)RR7qqaRF:Rk#0R0D8_FOoH_OPC05FsRR4R8MFI0jFR2
R;RRRRRRRRRRRRRRRR)iBphRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRR)iBp RR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRR)R RRRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRR)7q7)RR:HRMR#_08DHFoOC_POs0F5jR4RFR8IFM0RRj2;R
RRRRRRRRRRRRRRBRWpRiR:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRBRWpRi :MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRR RWRRRR:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRqRW7R7):MRHR0R#8F_Do_HOP0COFRs54RjR8MFI0jFR2
R;RRRRRRRRRRRRRRRRWa7qqRR:HRMR#_08DHFoOC_POs0F5RR4RI8FMR0FjR2
RRRRRRRRRRRRR;R2
8CMRlOFbCFMM
0;
lOFbCFMM10RAq_)vc.jUhG.WR
RRRRRRRRRoCCMsRHO5hRQQja_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2
R;RRRRRRRRRRRRRRRRRRRRQahQ_:4RR0LH_OPC05FsR6.6RFR8IFM0RRj2;RR
RRRRRRRRRRRRRRRRRQRRh_Qa.RR:L_H0P0COFRs5.R66RI8FMR0Fj;2RRR
RRRRRRRRRRRRRRRRRRhRQQda_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2RR;
RRRRRRRRRRRRRRRRRRRRQQhaR_c:HRL0C_POs0F56R.68RRF0IMF2RjR
;RRRRRRRRRRRRRRRRRRRRRQahQ_:6RR0LH_OPC05FsR6.6RFR8IFM0RRj2;R
RRRRRRRRRRRRRRRRRRhRQQna_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2
R;RRRRRRRRRRRRRRRRRRRRQahQ_:(RR0LH_OPC05FsR6.6RFR8IFM0RRj2;R
RRRRRRRRRRRRRRRRRRhRQQUa_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2
R;RRRRRRRRRRRRRRRRRRRRQahQ_:gRR0LH_OPC05FsR6.6RFR8IFM0RRj2;R
RRRRRRRRRRRRRRRRRRhRQQqa_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2
R;RRRRRRRRRRRRRRRRRRRRQahQ_:ARR0LH_OPC05FsR6.6RFR8IFM0RRj2;R
RRRRRRRRRRRRRRRRRRhRQQBa_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2
R;RRRRRRRRRRRRRRRRRRRRQahQ_:7RR0LH_OPC05FsR6.6RFR8IFM0RRj2;R
RRRRRRRRRRRRRRRRRRhRQQ a_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2
R;RRRRRRRRRRRRRRRRRRRRQahQ_:wRR0LH_OPC05FsR6.6RFR8IFM0RRj2
RRRRRRRRRRRRRRRR2RRRR;
RRRRRRRRRsbF0
5RRRRRRRRRRRRRRRRR)a7qqRR:FRk0#_08DHFoOC_POs0F5RR4RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRp)BiRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRR)iBp RR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRR)R RRRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRR)7q7)RR:HRMR#_08DHFoOC_POs0F5jR4RFR8IFM0RRj2;R
RRRRRRRRRRRRRRBRWpRihRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRRWRRB piRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRRWRR RRRRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRRWRRq)77RH:RM#RR0D8_FOoH_OPC05FsRR4jRI8FMR0Fj;2R
RRRRRRRRRRRRRRRRqW7a:qRRRHMR8#0_oDFHPO_CFO0s45RRFR8IFM0R
j2RRRRRRRRRRRRR2RR;M
C8FROlMbFC;M0
F
OlMbFCRM01)A_qjv.c.UGhW)h
RRRRRRRRoRRCsMCH5ORRQQhaR_j:HRL0C_POs0F56R.68RRF0IMF2RjRR;
RRRRRRRRRRRRRRRRRQRRh_Qa4RR:L_H0P0COFRs5.R66RI8FMR0Fj;2RRR
RRRRRRRRRRRRRRRRRRhRQQ.a_RL:RHP0_CFO0s.5R6R6R8MFI0jFR2RR;
RRRRRRRRRRRRRRRRRRRRQQhaR_d:HRL0C_POs0F56R.68RRF0IMF2RjR
;RRRRRRRRRRRRRRRRRRRRRQahQ_:cRR0LH_OPC05FsR6.6RFR8IFM0RRj2;RR
RRRRRRRRRRRRRRRRRQRRh_Qa6RR:L_H0P0COFRs5.R66RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRRRRRQQhaR_n:HRL0C_POs0F56R.68RRF0IMF2RjRR;
RRRRRRRRRRRRRRRRRQRRh_Qa(RR:L_H0P0COFRs5.R66RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRRRRRQQhaR_U:HRL0C_POs0F56R.68RRF0IMF2RjRR;
RRRRRRRRRRRRRRRRRQRRh_QagRR:L_H0P0COFRs5.R66RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRRRRRQQhaR_q:HRL0C_POs0F56R.68RRF0IMF2RjRR;
RRRRRRRRRRRRRRRRRQRRh_QaARR:L_H0P0COFRs5.R66RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRRRRRQQhaR_B:HRL0C_POs0F56R.68RRF0IMF2RjRR;
RRRRRRRRRRRRRRRRRQRRh_Qa7RR:L_H0P0COFRs5.R66RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRRRRRQQhaR_ :HRL0C_POs0F56R.68RRF0IMF2RjRR;
RRRRRRRRRRRRRRRRRQRRh_QawRR:L_H0P0COFRs5.R66RI8FMR0Fj
2RRRRRRRRRRRRRRRRRRRR2;R
RRRRRRRRRb0Fs5RR
RRRRRRRRRRRRR)RR7qqaRF:Rk#0R0D8_FOoH_OPC05FsRR4R8MFI0jFR2
R;RRRRRRRRRRRRRRRR)iBphRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRR)iBp RR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRR)R RRRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRR)7q7)RR:HRMR#_08DHFoOC_POs0F5jR4RFR8IFM0RRj2;R
RRRRRRRRRRRRRRBRWpRihRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRRWRRB piRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRRWRR RRRRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRRWRRq)77RH:RM#RR0D8_FOoH_OPC05FsRR4jRI8FMR0Fj;2R
RRRRRRRRRRRRRRRRqW7a:qRRRHMR8#0_oDFHPO_CFO0s45RRFR8IFM0R
j2RRRRRRRRRRRRR2RR;M
C8FROlMbFC;M0
F
OlMbFCRM01QA_mR
RRRRRRRRRoCCMsRHO5QRuhY_auR RRRR:L_H0P0COFRs568RRF0IMF2Rj;R
RRRRRRRRRRRRRRRRRRzRupupzR:RRR0LH;RR
RRRRRRRRRRRRRRRRRhRR at_)tQt :)RR0LH;RR
RRRRRRRRRRRRRRRRRQRRma_1qqh7):7RRs#0HRMo
RRRRRRRRRRRRRRRR2RRRR;
RRRRRRRRRsbF0
5RRRRRRRRRRRRRRRRRuiqBq_t uRQhRRRRR:RRRFHMk#0R0D8_FOoHRR;
RRRRRRRRRRRRRpRRq]aB_uQhzea_q pzRRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRRBBpmih_ q ApRRRRR:RRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRuQhzBa_pRiRRRRRRRRR:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRzRmaauz_iBpRRRRRRRRRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRRmRRzzauah_ q ApRRRRRRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRR7z_maR_4RRRRRRRRR:RRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRm7_zja_RRRRRRRRRRRR:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRR_R7Q4h_RRRRRRRRRRRRRF:Rk#0R0D8_FOoHRR;
RRRRRRRRRRRRR7RR__QhjRRRRRRRRRRRRRR:FRk0#_08DHFoORRRRRRRRRRRRRRRRRR
RRRRRRRRRRRRR;R2
8CMRlOFbCFMM
0;
lOFbCFMM10RAA_t_
QmRRRRRRRRRCRoMHCsORR5u_Qha YuRRRR:HRL0C_POs0F5RR6RI8FMR0Fj
2;RRRRRRRRRRRRRRRRRRRRupzpzRuRRL:RHR0;
RRRRRRRRRRRRRRRRRRRRth _Qa)t)t RL:RHR0;
RRRRRRRRRRRRRRRRRRRR_Qm1haq77q)R#:R0MsHoRR
RRRRRRRRRRRRRRRRR;2R
RRRRRRRRbRRF5s0RR
RRRRRRRRRRRRRRqRuBtiq Q_uhRRRRRRRR:RRRFHMk#0R0D8_FOoHRR;
RRRRRRRRRRRRRpRRq]aB_uQhzea_q pzRRRR:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRpRBm_Bi AhqpR RRRRRR:RRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRuQhzBa_pRiRRRRRRRRRRRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRRmuzazBa_pRiRRRRRRRRRRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRRmRRzzauah_ q ApRRRRRRRR:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRR_R7m_za4RRRRRRRRRRRR:RRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRm7_zja_RRRRRRRRRRRRRRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRR7h_Q_R4RRRRRRRRRRRRRRF:Rk#0R0D8_FOoHRR;
RRRRRRRRRRRRR7RR__QhjRRRRRRRRRRRRRRR:kRF00R#8F_DoRHO;R
RRRRRRRRRRRRRRpRtmpAq_wAzw_ )muzaz:aRR0FkR8#0_oDFHRORRRRRRRRRRRRRRRR
RRRRRRRRRRRRR;R2
8CMRlOFbCFMM
0;
lOFbCFMM10RAm_Q_
71RRRRRRRRRCRoMHCsORR5u_Qha YuRRRR:HRL0C_POs0F5RR6RI8FMR0Fj
2;RRRRRRRRRRRRRRRRRRRRh_ tat)QtR ):HRL0
;RRRRRRRRRRRRRRRRRRRRRQ1m_a7qhqR)7:0R#soHMRR
RRRRRRRRRRRRRRRRR2
R;RRRRRRRRRFRbsR05
RRRRRRRRRRRRRRRRBuqi qt_huQRRRRRRRR:MRHFRk0#_08DHFoO
R;RRRRRRRRRRRRRRRRuiqBq_t u_QhARRRR:RRRFHMk#0R0D8_FOoHRR;
RRRRRRRRRRRRRpRRq]aB_uQhzea_q pzRRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRRBBpmih_ q ApRRRRR:RRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRuQhzBa_pRiRRRRRRRRR:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRzRmaauz_iBpRRRRRRRRRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRRmRRzzauah_ q ApRRRRRRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRR7z_maR_4RRRRRRRRR:RRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRm7_zja_RRRRRRRRRRRR:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRR_R7Q4h_RRRRRRRRRRRRRF:Rk#0R0D8_FOoHRR;
RRRRRRRRRRRRR7RR__QhjRRRRRRRRRRRRRR:FRk0#_08DHFoORRRRRRRRRRRRRRRRRR
RRRRRRRRRRRRR;R2
8CMRlOFbCFMM
0;
lOFbCFMM10RAA_t
RRRRRRRRbRRF5s0RR
RRRRRRRRRRRRRRpRtmpAq_wAzw_ )muzazRaRRRRRR:RRR0FkR8#0_oDFH;OR
RRRRRRRRRRRRRRRR z1)Q_1tphq__amtApmqAp_z ww)RR:HRMR#_08DHFoORR
RRRRRRRRRRRRR;R2
8CMRlOFbCFMM
0;
lOFbCFMM10RAp_up_cjB m)RR
RoCCMsRHO5R
RRRRRR-SS-w-RCLC8N
O	S Sw q7ABui_qSa]RRSS:0R#soHMRR:="v1Qu"p ;-R-Rs10HRMo5l#Hb,DCRD8CNR$,b#ENCM_N8C_8D,N$R0CGCNsMD
2SS S7p_qYqz7K1 avhva_m_7 w7  AiqBR:SRRs#0HRMo:"=Rw QX7R";
7SS Ypq_Kq7zv1a _hav m7_p) qeaQ RRS:0R#soHMRR:="XwQ ;7"RS
S1w]Qat) _e7Q_7vm SRS:HRL0C_POs0F584RF0IMF2RjSR:=""jj;RRS-R-Rj>--7HHP8LCR$,RcR-4->P7HHR8CL($R,RRd-7->H8PHC$RLR
6SSSRRw_7qw7  AiqBRSSS:HRL0C_POs0F58dRF0IMF2RjR=S:Rj"jj;j"R-SR-QRRMo0CC5sRj6-42
3RS7Swq _)pQqaeS RSRS:L_H0P0COFds5RI8FMR0Fj:2S=jR"j"jj;RRS-R-RQCM0oRCs54j-6R23R
RSRSRSumppz1a_ Bp aSSSR#:R0MsHo=R:R "thiBp"
;
RSRS-R--zR#C0REC#CbsN#8RE0CCRR0FbkFbDCN0RC0ERDPNkRC#LFCDIS
S7wQeSSSS:HRL0C_POs0F58nRF0IMF2Rj;-RR-CR70lCsHRMCNFRoF88RCkVNDP0RNCDk
7SSQSe)S:SSR0LH_OPC05FsdFR8IFM0R;j2R-R-R07CCHslMNCRRFoF8CR8VDNk0NRPD
kCSQS7eSTSSRS:L_H0P0COF.s5RI8FMR0FjR2;RR--7CC0sMlHCRRNo8FFRV8CN0kDRDPNkSC
SpwQa_ ))tqh SSS:HRL0C_POs0F58.RF0IMF2Rj;-RR-CR70lCsHRMCNFRoF88RCkVNDP0RNCDkRR

R-SS-q-R808HHNFMD-RBA#H0
SRRSq hA_p QtB qSa SRS:LRH0:'=Rj
';
SRRS---R#aC0FRv8uCRNlsNCs0CRR
RS Sa1va_mS7 SRS:LRH0:'=Rj
';SXS ah )q7p_Q7eQ q_wB)amSRS:HCM0oRCs:4=RRR--hRF0z8#CRRL$lCF8Dq,R888CRsVFRpupRMOFVRHot
zQRRRRR2RR;R
Rb0FsRR5
RRRRR)RR )w   hBBSpiSH:RM0R#8F_Do;HOSRSSR-RR-sR7HMPCRRL$OCFsRoDFHRO
RRRRRuRRpzpma)Bm :SSR0FkR8#0_oDFHSO;SRRRRR--uRppFbk0k00RFFROsDCRFOoH
RRRRRRRRpupmtzapqmAp:SSR0FkR8#0_oDFHSO;SRRRRR--uRppFbk0k00RFDRoFDLNR0MCI	Fs
RRRRRRRRa Xw7  AiqBSRS:H#MR0D8_FOoH;SSSRRRR-7-RsCHPM$RLRsOFCFRDo
HOSh7YqBvQ7q pY:SSRRHM#_08DHFoOC_POs0FRR5(8MFI0jFR2-;R-sR7HMPCRRL$OCFsRoDFHRO
RRRRRpRRmSBiSRS:FRk0#_08DHFoOR;SSRRRRR--mbk0kF0RVpRupR
RRRRRRYRAu1q1S:SSRRHM#_08DHFoOS;SSRRRRR--7PsHCLMR$FROsDCRFOoH
RRRRRRRR1)  SaASRS:H#MR0D8_FOoH;SSSRRRR-7-RsCHPM$RLRsOFCFRDo
HORRRRRRRRpBqa]uQhzqaepSz SH:RM0R#8F_Do;HOSRSSR-RR-BRH 0tNCHR1oDMN
SRR-a-RCR#0u#HM
SRR1S7mSRS:FRk0#_08DHFoOS;SRRRR-m-Rkk0b0VRFRpup
SRR1S7QSRS:H#MR0D8_FOoH;SSSRRRR-7-RsCHPM$RLRsOFCFRDo
HOR1RSBSpiSRS:H#MR0D8_FOoHSRSSR-RR-sR7HMPCRRL$OCFsRoDFHRO
RRRRR;R2
8CMRlOFbCFMM
0;
lOFbCFMMR0R1uA_pjpc_)Bm z_7uBpQqRa 
CSoMHCsOSR5
wSS A 7q_Biu]qaRSSS:0R#soHMRSSS:"=R1uQvp; "S-R-Rs10HRMoRH5#lCbD,CR8D,N$RNbE#NC_M88_C$DN,GRC0MCsNRD2
7SS Ypq_Kq7zv1a _hav m7_ w 7BAqi:RRRs#0HRMoS:SS=wR"Q7X "
;RS S7p_qYqz7K1 avhva_m_7 )q pa QeRRS:#H0sMSoSSR:="XwQ ;7"RS
S1w]Qat) _e7Q_7vm SRS:HRL0C_POs0F584RF0IMF2RjSR:=""jj;RRS-R-Rj>--7HHP8LCR$,RcR-4->P7HHR8CL($R,RRd-7->H8PHC$RLR
6SS7Swq _w q7ABSiRSRS:L_H0P0COFds5RI8FMR0FjS2R:"=Rjjjj"S;RRR--R0QMCsoCR-5j4362RS
Sw_7q)q pa QeRSSS:HRL0C_POs0F58dRF0IMF2RjSR:="jjjjR";S-R-RMRQ0CCosjR5-2463RRRRS
Sumppz1a_ Bp aSRSS#:R0MsHoSRSSR:="ht B"pi;
RRSQS7eS)RS:SSR0LH_OPC05FsdFR8IFM0RSj2:"=Rjjjj"S;R
7SSQRewSSSS:HRL0C_POs0F58nRF0IMF2RjR=S:Rj"jjjjjjR";
7SSQReTSSSS:HRL0C_POs0F58.RF0IMF2RjSR:="jjj"S;RSS
SwaQp ))_q htRSSS:HRL0C_POs0F58.RF0IMF2RjRRRRRRRR:"=Rj"jj;
RSShS q Ap_ QBt qaS:SSR0LHSSSS:'=Rj
';S Sa1va_mR7 S:SSR0LHSSSS:'=Rj
';SXS ah )q7p_Q7eQ q_wB)amR:SSR0HMCsoCRSSSSR:=4SRSRh--Fk0R#RC8Ll$RFD8C38Rq8RC8VRFsuRppBVFMHtoRz
Q3R2SR;S

b0FsR
S5S S)w  )hBB pSiSSH:RM0R#8F_DoRHO;SRS-7-RsCHPM$RLRsOFCFRDo
HOSpSupamzB m)S:SSR0FkR8#0_oDFHRO;S-S-RpupR0FkbRk00OFRFRsCDHFoORR5LM$RFNslDFRskM0Ho
2RSpSupamztApmqRpSRSRS:kRF00R#8F_Do;HOR-SS-pRupkRF00bkRR0FOCFsRoDFHROR5RL$oLDFNMDRCF0Is
	2SXS a w 7BAqiSRRSRS:H#MR0D8_FOoH;SSS-7-RsCHPM$RLRsOFCFRDo
HOSYS7hQqvBp7 qSYSSH:RM0R#8F_Do_HOP0COF5sR(FR8IFM0R;j2SR--7PsHCLMR$FROsDCRFOoH
pSSmSBiS:SSR0FkR8#0_oDFHRO;S-S-R0mkbRk0FuVRpSp
SuAYqS11S:SSRRHM#_08DHFoOS;RSR--7PsHCLMR$FROsDCRFOoH
)SS a1 ASSSSH:RM0R#8F_Do;HOR-SS-sR7HMPCRRL$OCFsRoDFHSO
SQ17SSSS:MRHR8#0_oDFHRO;S-S-RH7sPRCMLO$RFRsCDHFoOa3RCR#0u
HMS7S1mSSSSF:Rk#0R0D8_FOoH;-SS-kRm00bkRR0F)pARFOoHRDaHCa3RCR#0u
HMSBS1pSiSSRS:H#MR0D8_FOoH;SRS-7-RsCHPM$RLRsOFCFRDo3HOR#aC0HRuMS
SpBqa]uQhzqaepRz SRS:H#MR0D8_FOoHRSSS-H-RBN t0#CRHNoMDSS
RRRRR2RR;CR
MO8RFFlbM0CM;SSS
F
OlMbFCRM01uA_pjpc_7uq
R
RoCCMsRHO5R
RS-S--CRwCN8LOS	
S w 7BAqiq_uaR]SS:SRRs#0HRMo:"=R1uQvp; "RR--1H0sM5oR#bHlDRC,8NCD$b,RECN#_8NM_D8CNR$,CCG0sDMN2SS
Sp7 qqY_71Kzahv am_v7w _ A 7qRBiSRR:#H0sM:oR=wR"Q7X "
;RS S7p_qYqz7K1 avhva_m_7 )q pa QeR:SRRs#0HRMo:"=Rw QX7R";
1SS]aQw)_ t7_Qev m7R:SSR0LH_OPC05Fs4FR8IFM0RSj2:"=Rj;j"R-SR-jRR-7->H8PHC$RLRRc,4>--7HHP8LCR$,R(R-dR-H>7PCH8RRL$6S
Sw_7qw7  AiqBRSSS:HRL0C_POs0F58dRF0IMF2RjR=S:Rj"jj;j"R-SR-QRRMo0CC5sRj6-42
3RS7Swq _)pQqaeS RSRS:L_H0P0COFds5RI8FMR0Fj:2S=jR"j"jj;RRS-R-RQCM0oRCs54j-6R23RRRSRR
RSpSupamz_p1  SBaS:SRRs#0HRMo:"=RtB hp;i"
R
RS-S--#RzCER0CbR#s8CNRC#EC00RFFRbbNkD00CREPCRNCDk#CRLD
FISQS7eSwSSRS:L_H0P0COFns5RI8FMR0FjR2;RR--7CC0sMlHCRRNo8FFRV8CN0kDRDPNkSC
Se7Q)SSSSL:RHP0_CFO0sR5d8MFI0jFR2R;R-7-RCs0ClCHMRoNRFRF88NCVkRD0PkNDCS
S7TQeSSSS:HRL0C_POs0F58.RF0IMF2Rj;-RR-CR70lCsHRMCNFRoF88RCkVNDP0RNCDk
wSSQ pa)q_)hSt SRS:L_H0P0COF.s5RI8FMR0FjR2;RR--7CC0sMlHCRRNo8FFRV8CN0kDRDPNk
CR
SRRS---R8q8HF0HMRNDBH-A0R#
R SShpqA B_Q atq SSS:HRL0=R:R''j;R

R-SS-a-RCR#0vCF8RsuNN0lCC
sRRSRSaa 1_7vm SSS:HRL0=R:R''j;S
S  Xa)phq_e7QQ_7 waqBmS)S:MRH0CCos=R:R-4R-FRh0#RzCL8R$FRl8,CDR8q8CV8RFusRpOpRFHMVozRtQR
RRRRRR
2;RFRbs50RRR
RRRRRRqRuBtiq huQSRS:HkMF00R#8F_Do;HOSRSRRRR
RRRRRuRRpzpma)Bm :SSR0FkR8#0_oDFHSO;SRRRRR--uRppFbk0k00RFFROsDCRFOoH
RRRRRRRRpupmtzapqmAp:SSR0FkR8#0_oDFHSO;SRRRRR--uRppFbk0k00RFDRoFDLNR0MCI	Fs
RRRRRRRRa Xw7  AiqBSRS:H#MR0D8_FOoH;SSSRRRR-7-RsCHPM$RLRsOFCFRDo
HOSh7YqBvQ7q pY:SSRRHM#_08DHFoOC_POs0FRR5(8MFI0jFR2-;R-sR7HMPCRRL$OCFsRoDFHRO
RRRRRpRRmSBiSRS:FRk0#_08DHFoOS;SRRRR-m-Rkk0b0VRFRpup
RRRRRRRRuAYqS11SRS:H#MR0D8_FOoH;SSSRRRR-7-RsCHPM$RLRsOFCFRDo
HORRRRRRRR)  1aSASSH:RM0R#8F_Do;HOSRSSR-RR-sR7HMPCRRL$OCFsRoDFHRO
RRRRRpRRq]aBQzhuapeqzS S:MRHR8#0_oDFHSO;SRSRR-R-R HBtCN0Ro1HM
NDR-RS-CRa#u0RH
M#R1RS7SmSSF:Rk#0R0D8_FOoH;RSSR-RR-kRm00bkRRFVu
ppR1RS7SQSSH:RM0R#8F_Do;HOSRSSR-RR-sR7HMPCRRL$OCFsRoDFHRO
RBS1pSiSSH:RM0R#8F_DoSHOSRSRR-R-RH7sPRCMLO$RFRsCDHFoOR
RRRRRR
2;RCR
MO8RFFlbM0CM;


ObFlFMMC0AR1_pupc.j__7uq
R
RoCCMsRHO5R
RS-S--CRwCN8LOS	
S w 7BAqiq_uaR]SS:SRRs#0HRMo:"=R1uQvp; "RR--1H0sM5oR#bHlDRC,8NCD$b,RECN#_8NM_D8CNR$,CCG0sDMN2SS
Sp7 qqY_71Kzahv am_v7w _ A 7qRBiSRR:#H0sM:oR=wR"Q7X "
;RS S7p_qYqz7K1 avhva_m_7 )q pa QeR:SRRs#0HRMo:"=Rw QX7R";
1SS]aQw)_ t7_Qev m7R:SSR0LH_OPC05Fs4FR8IFM0RSj2:"=Rj;j"R-SR-jRR-7->H8PHC$RLRRc,4>--7HHP8LCR$,R(R-dR-H>7PCH8RRL$6S
Sw_7qw7  AiqBRSSS:HRL0C_POs0F58dRF0IMF2RjR=S:Rj"jj;j"R-SR-QRRMo0CC5sRj6-42
3RS7Swq _)pQqaeS RSRS:L_H0P0COFds5RI8FMR0Fj:2S=jR"j"jj;RRS-R-RQCM0oRCs54j-6R23RRRSRR
RSpSupamz_p1  _Bauam)ARSS:0R#soHMRR:="ht B"pi;R

R-SS-z-R#0CRE#CRbNsC8ER#CRC00bFRFDbkNR0C0RECPkNDCL#RCIDF
7SSQSewS:SSR0LH_OPC05FsnFR8IFM0R;j2R-R-R07CCHslMNCRRFoF8CR8VDNk0NRPD
kCSQS7eS)SSRS:L_H0P0COFds5RI8FMR0FjR2;RR--7CC0sMlHCRRNo8FFRV8CN0kDRDPNkSC
Se7QTSSSSL:RHP0_CFO0sR5.8MFI0jFR2R;R-7-RCs0ClCHMRoNRFRF88NCVkRD0PkNDCS
SwaQp ))_q htS:SSR0LH_OPC05Fs.FR8IFM0R;j2R-R-R07CCHslMNCRRFoF8CR8VDNk0NRPDRkC
R
RS-S--8Rq8HH0FDMNRAB-H
0#RSRS AhqpQ _Bq tau _mq)aSRS:LRH0:'=Rj
';RSRS AhqpQ _Bq tau _mA)aSRS:LRH0:'=Rj
';
SRRS---R#aC0FRv8uCRNlsNCs0CRR
RS Sa1va_mS7 SRS:LRH0:'=Rj
';SXS ah )q7p_Q7eQ q_wB)amSRS:HCM0oRCs:4=RRR--hRF0z8#CRRL$lCF8Dq,R888CRsVFRpupRMOFVRHot
zQRRRRR2RR;R
Rb0FsR
5RRRRRRRRRuiqBqut QShS:MRHFRk0#_08DHFoOS;SRRRR
RRRRRRRRpupmBzamq) SRS:FRk0#_08DHFoOS;SRRRR-u-RpFpRkk0b0FR0RsOFCFRDo
HORRRRRRRRumppzpatmpAqq:SSR0FkR8#0_oDFHSO;SRRRRR--uRppFbk0k00RFDRoFDLNR0MCI	Fs
RRRRRRRRpupmBzamA) SRS:FRk0#_08DHFoOS;SRRRR-u-RpFpRkk0b0FR0RsOFCFRDo
HORRRRRRRRumppzpatmpAqA:SSR0FkR8#0_oDFHSO;SRRRRR--uRppFbk0k00RFDRoFDLNR0MCI	Fs
RRRRRRRRa Xw7  AiqBSRS:H#MR0D8_FOoH;SSSRRRR-7-RsCHPM$RLRsOFCFRDo
HOSh7YqBvQ7q pY:SSRRHM#_08DHFoOC_POs0FRR5(8MFI0jFR2-;R-sR7HMPCRRL$OCFsRoDFHRO
RRRRRpRRmSBiSRS:FRk0#_08DHFoOS;SRRRR-m-Rkk0b0VRFRpup
RRRRRRRRuAYqS11SRS:H#MR0D8_FOoH;SSSRRRR-7-RsCHPM$RLRsOFCFRDo
HORRRRRRRR)  1aSASSH:RM0R#8F_Do;HOSRSSR-RR-sR7HMPCRRL$OCFsRoDFHRO
RRRRRpRRq]aBQzhuapeqzS S:MRHR8#0_oDFHSO;SRSRR-R-R HBtCN0Ro1HM
NDR-RS-CRa#u0RH
M#R1RS7SmSSF:Rk#0R0D8_FOoH;RSSR-RR-kRm00bkRRFVu
ppR1RS7SQSSH:RM0R#8F_Do;HOSRSSR-RR-sR7HMPCRRL$OCFsRoDFHRO
RBS1pSiSSH:RM0R#8F_DoSHOSRSRR-R-RH7sPRCMLO$RFRsCDHFoOR
RRRRRR
2;RCR
MO8RFFlbM0CM;O

FFlbM0CMR_1Aucppjw_._)Bm R

RMoCCOsHRR5
R-SS-w-RCLC8N
O	S Sw q7ABui_qSa]RRSS:0R#soHMRR:="v1Qu"p ;-R-Rs10HRMo5l#Hb,DCRD8CNR$,b#ENCM_N8C_8D,N$R0CGCNsMD
2SS S7p_qYqz7K1 avhva_m_7 w7  AiqBR:SRRs#0HRMo:"=Rw QX7R";
7SS Ypq_Kq7zv1a _hav m7_p) qeaQ RRS:0R#soHMRR:="XwQ ;7"RS
S1w]Qat) _e7Q_7vm SRS:HRL0C_POs0F584RF0IMF2RjSR:=""jj;RRS-R-Rj>--7HHP8LCR$,RcR-4->P7HHR8CL($R,RRd-7->H8PHC$RLRS6
Sqw7_ w 7BAqiSRSSL:RHP0_CFO0sR5d8MFI0jFR2:RS=jR"j"jj;RRS-R-RQCM0oRCs54j-6R23
wSS7)q_ apqQRe S:SSR0LH_OPC05FsdFR8IFM0RSj2:"=Rjjjj"S;RRR--R0QMCsoCR-5j4362RRRR
SRRSpupm_za1  pBua_mq)aS:SRRs#0HRMo:"=RtB hp;i"
SRRSpupm_za1  pBua_mA)aS:SRRs#0HRMo:"=RtB hp;i"
R
RS-S--#RzCER0CbR#s8CNRC#EC00RFFRbbNkD00CREPCRNCDk#CRLD
FISQS7eSwSSRS:L_H0P0COFns5RI8FMR0FjR2;RR--7CC0sMlHCRRNo8FFRV8CN0kDRDPNkSC
Se7Q)SSSSL:RHP0_CFO0sR5d8MFI0jFR2R;R-7-RCs0ClCHMRoNRFRF88NCVkRD0PkNDCS
S7TQeSSSS:HRL0C_POs0F58.RF0IMF2Rj;-RR-CR70lCsHRMCNFRoF88RCkVNDP0RNCDk
wSSQ pa)q_)hSt SRS:L_H0P0COF.s5RI8FMR0FjR2;RR--7CC0sMlHCRRNo8FFRV8CN0kDRDPNk
CR
SRRS---R8q8HF0HMRNDBH-A0R#
R SShpqA B_Q atq m_u)SaqSL:RH:0R=jR''R;
R SShpqA B_Q atq m_u)SaASL:RH:0R=jR''
;
RSRS-R--a0C#R8vFCNRusCNl0RCs
SRRS1a am_v7S SSL:RH:0R=jR''S;
Sa X q)hpQ_7e Q7_BwqaSm)SH:RMo0CC:sR=RR4-h-RFz0R#RC8Ll$RFD8C,8Rq8RC8VRFsuRppOVFMHtoRzRQ
RRRRR;R2
bRRFRs05RR
RRRRR)RR )w   hBBSpiSH:RM0R#8F_Do;HOSRSRRRRSR-RR-sR7HMPCRRL$OCFsRoDFHRO
RRRRRuRRpzpma)Bm SqS:kRF00R#8F_Do;HOSRSRR-R-RpupR0FkbRk00OFRFRsCDHFoOR
RRRRRRpRupamztApmqSpqSF:Rk#0R0D8_FOoH;RSSR-RR-pRupkRF00bkRR0FoLDFNMDRCF0IsR	
RRRRRuRRpzpma)Bm SAS:kRF00R#8F_Do;HOSRSRR-R-RpupR0FkbRk00OFRFRsCDHFoOR
RRRRRRpRupamztApmqSpASF:Rk#0R0D8_FOoH;RSSR-RR-pRupkRF00bkRR0FoLDFNMDRCF0IsR	
RRRRR RRX aw q7ABSiS:MRHR8#0_oDFHSO;SRSRR-R-RH7sPRCMLO$RFRsCDHFoO7
SYvhqQ B7pSqYSH:RM0R#8F_Do_HOP0COF5sR(FR8IFM0R;j2RR--7PsHCLMR$FROsDCRFOoH
RRRRRRRRBpmiSSS:kRF00R#8F_Do;HOSRSRR-R-R0mkbRk0FuVRpRp
RRRRRARRY1uq1SSS:MRHR8#0_oDFHSO;SRSRR-R-RH7sPRCMLO$RFRsCDHFoOR
RRRRRR R)1A aS:SSRRHM#_08DHFoOS;SSRRRRR--7PsHCLMR$FROsDCRFOoH
RRRRRRRRapqBh]Quezaq pzSRS:H#MR0D8_FOoH;SSSRRRR-H-RBN t01CRHNoMDR
RSR--a0C#RMuH#R
RSm17S:SSR0FkR8#0_oDFHSO;SRRRRR--mbk0kF0RVpRupR
RSQ17S:SSRRHM#_08DHFoOS;SSRRRRR--7PsHCLMR$FROsDCRFOoH
SRR1iBpS:SSRRHM#_08DHFoOSSSRRRR-7-RsCHPM$RLRsOFCFRDo
HORRRRR2RR;R
R
8CMRlOFbCFMM
0;
lOFbCFMM10RAp_up_cj.uw_q
7
RCRoMHCsO
R5RSRS-R--w8CCL	NO
wSS A 7q_Biu]qaSSRSR#:R0MsHo=R:RQ"1v up"-;R-0R1soHMRH5#lCbD,CR8D,N$RNbE#NC_M88_C$DN,GRC0MCsNSD2
7SS Ypq_Kq7zv1a _hav m7_ w 7BAqiRRS:0R#soHMRR:="XwQ ;7"RS
S7q pY7_qKaz1va h_7vm  _)pQqaeS RR#:R0MsHo=R:RQ"wX" 7;SR
SQ1]w a)tQ_7em_v7S RSL:RHP0_CFO0sR548MFI0jFR2=S:Rj"j"S;RRR--R-j->P7HHR8CLc$R,-R4-H>7PCH8RRL$(d,RR>--7HHP8LCR$
R6S7Swq _w q7ABSiRSRS:L_H0P0COFds5RI8FMR0FjS2R:"=Rjjjj"S;RRR--R0QMCsoCR-5j4362RS
Sw_7q)q pa QeRSSS:HRL0C_POs0F58dRF0IMF2RjSR:="jjjjR";S-R-RMRQ0CCosjR5-2463RRRRR
RSpSupamz_p1  _Bauam)qRSS:0R#soHMRR:="ht B"pi;R
RSpSupamz_p1  _Bauam)ARSS:0R#soHMRR:="ht B"pi;R

R-SS-z-R#0CRE#CRbNsC8ER#CRC00bFRFDbkNR0C0RECPkNDCL#RCIDF
7SSQSewS:SSR0LH_OPC05FsnFR8IFM0R;j2R-R-R07CCHslMNCRRFoF8CR8VDNk0NRPD
kCSQS7eS)SSRS:L_H0P0COFds5RI8FMR0FjR2;RR--7CC0sMlHCRRNo8FFRV8CN0kDRDPNkSC
Se7QTSSSSL:RHP0_CFO0sR5.8MFI0jFR2R;R-7-RCs0ClCHMRoNRFRF88NCVkRD0PkNDCS
SwaQp ))_q htS:SSR0LH_OPC05Fs.FR8IFM0R;j2R-R-R07CCHslMNCRRFoF8CR8VDNk0NRPDRkC
R
RS-S--8Rq8HH0FDMNRAB-H
0#RSRS AhqpQ _Bq tau _mq)aSRS:LRH0:'=Rj
';RSRS AhqpQ _Bq tau _mA)aSRS:LRH0:'=Rj
';
SRRS---R#aC0FRv8uCRNlsNCs0CRR
RS Sa1va_mS7 SRS:LRH0:'=Rj
';SXS ah )q7p_Q7eQ q_wB)amSRS:HCM0oRCs:4=RRR--hRF0z8#CRRL$lCF8Dq,R888CRsVFRpupRMOFVRHot
zQRRRRR2RR;R
Rb0FsR
5RRRRRRRRRuiqBqut QShS:MRHFRk0#_08DHFoOR;SRSRRRRRR
RRRRRRRRpupmBzamq) SRS:FRk0#_08DHFoOS;SRRRR-u-RpFpRkk0b0FR0RsOFCFRDo
HORRRRRRRRumppzpatmpAqq:SSR0FkR8#0_oDFHSO;SRRRRR--uRppFbk0k00RFDRoFDLNR0MCI	Fs
RRRRRRRRpupmBzamA) SRS:FRk0#_08DHFoOS;SRRRR-u-RpFpRkk0b0FR0RsOFCFRDo
HORRRRRRRRumppzpatmpAqA:SSR0FkR8#0_oDFHSO;SRRRRR--uRppFbk0k00RFDRoFDLNR0MCI	Fs
RRRRRRRRa Xw7  AiqBSRS:H#MR0D8_FOoH;SSSRRRR-7-RsCHPM$RLRsOFCFRDo
HOSh7YqBvQ7q pY:SSRRHM#_08DHFoOC_POs0FRR5(8MFI0jFR2-;R-sR7HMPCRRL$OCFsRoDFHRO
RRRRRpRRmSBiSRS:FRk0#_08DHFoOS;SRRRR-m-Rkk0b0VRFRpup
RRRRRRRRuAYqS11SRS:H#MR0D8_FOoH;SSSRRRR-7-RsCHPM$RLRsOFCFRDo
HORRRRRRRR)  1aSASSH:RM0R#8F_Do;HOSRSSR-RR-sR7HMPCRRL$OCFsRoDFHRO
RRRRRpRRq]aBQzhuapeqzS S:MRHR8#0_oDFHSO;SRSRR-R-R HBtCN0Ro1HM
NDR-RS-CRa#u0RH
M#R1RS7SmSSF:Rk#0R0D8_FOoH;RSSR-RR-kRm00bkRRFVu
ppR1RS7SQSSH:RM0R#8F_Do;HOSRSSR-RR-sR7HMPCRRL$OCFsRoDFHRO
RBS1pSiSSH:RM0R#8F_DoSHOSRSRR-R-RH7sPRCMLO$RFRsCDHFoOR
RRRRRR
2;RCR
MO8RFFlbM0CM;-

--------------------------------------------------------------------------------------------------
-RSSSS1SRAp_up_cju_q77S1RSSSS---
-------------------------------------------------------------------------------------------------O

FFlbM0CMRAR1_pupcuj_q77_1
RRSMoCCOsHR
5SS Sw q7ABui_qRa]S:SSRs#0HRMoS:SS=1R"Qpvu S";RR--1H0sMRoR5l#Hb,DCRD8CNR$,b#ENCM_N8C_8D,N$R0CGCNsMD
2RS S7p_qYqz7K1 avhva_m_7 w7  AiqBRRR:#H0sMSoRS=S:RQ"wX" 7;SR
Sp7 qqY_71Kzahv am_v7) _ apqQRe S#:R0MsHoSSS:"=Rw QX7R";
1SS]aQw)_ t7_Qev m7R:SSR0LH_OPC05Fs4FR8IFM0RSj2:"=Rj;j"R-SR-jRR-7->H8PHC$RLRRc,4>--7HHP8LCR$,R(R-dR-H>7PCH8RRL$6SS
Sqw7_ w 7BAqiSRSSL:RHP0_CFO0sR5d8MFI0jFR2:RS=jR"j"jj;RRS-R-RQCM0oRCs54j-6R23
wSS7)q_ apqQRe S:SSR0LH_OPC05FsdFR8IFM0RSj2:"=Rjjjj"S;RRR--R0QMCsoCR-5j4362RRRR
uSSpzpma _1pa BRSSS:0R#soHMRSSS:"=RtB hp;i"RSR
Se7Q)SRSSRS:L_H0P0COFds5RI8FMR0Fj:2S=jR"j"jj;
RSSQS7eSwRS:SSR0LH_OPC05FsnFR8IFM0RRj2SR:="jjjjjjj"
;RSQS7eSTRS:SSR0LH_OPC05Fs.FR8IFM0RSj2:"=Rj"jj;SRS
wSSQ pa)q_)hRt S:SSR0LH_OPC05Fs.FR8IFM0RRj2RRRRR:RR=jR"j;j"RSS
Sq hA_p QtB qSa SRS:LSH0S:SS=jR''S;
S1a am_v7S RSRS:LSH0S:SS=jR''S;
Sa X q)hpQ_7e Q7_BwqaRm)SRS:HCM0oRCsS:SS=RR4S-SR-0hFRCk#8$RLR8lFCRD3qC888FRVspRupFRBMoVHRQtz3S
RR
2;
FSbsS0R5R
SRRRRRuRSqqBitQ uhSSS:MRHFRk0#_08DHFoORR;S-S-RV)CCMsCOOCRD5	Ru#2RHNoMDER0soFkENRuOo	NCMuH3RRR
RSRRRRRRqSuBtiq huQASSS:MRHFRk0#_08DHFoORR;S-S-RV)CCMsCOOCRD5	Rh#2RHNoMDER0soFkENRuOo	NCMuHAR3RRS
SumppzmaB)S SSF:Rk#0R0D8_FOoH;SRS-u-RpFpRkk0b0FR0RsOFCFRDoRHO5RL$MlFsNsDRFHk0M
o2SpSupamztApmqRpSRSRS:kRF00R#8F_Do;HOR-SS-pRupkRF00bkRR0FOCFsRoDFH5ORLo$RDNFLDCRM0sIF	S2
Sa Xw7  AiqBRSRSSH:RM0R#8F_Do;HOS-SS-sR7HMPCRRL$OCFsRoDFHSO
Sh7YqBvQ7q pYSSS:MRHR8#0_oDFHPO_CFO0s(R5RI8FMR0FjS2;-7-RsCHPM$RLRsOFCFRDo
HOSmSpBSiSSRS:FRk0#_08DHFoOS;RSR--mbk0kF0RVpRupS
SAqYu1S1SSRS:H#MR0D8_FOoH;SRS-7-RsCHPM$RLRsOFCFRDo
HOS S)1A aSSSS:MRHR8#0_oDFHRO;S-S-RH7sPRCMLO$RFRsCDHFoOS
S1S7QS:SSRRHM#_08DHFoOS;RSR--7PsHCLMR$FROsDCRFOoH3CRa#u0RHSM
Sm17SSSS:kRF00R#8F_Do;HOS-S-R0mkbRk00)FRAFRpoRHOaCHD3CRa#u0RHSM
Sp1BiSSSSH:RM0R#8F_Do;HOR-SS-sR7HMPCRRL$OCFsRoDFHRO3a0C#RMuH
pSSq]aBQzhuapeqzS RSH:RM0R#8F_DoRHOS-SS-BRH 0tNCHR#oDMNSR
SRRRRR;R2RM
C8FROlMbFC;M0R
S
---------------------------------------------------------------------------------------------------
-SRSSRSS1uA_pjpc__.wu_q77S1RSSSS---
-------------------------------------------------------------------------------------------------O

FFlbM0CMRAR1_pupc.j_wq_u71_7RSR
oCCMsRHO5SS
S w 7BAqiq_uaS]RSRS:#H0sMSoRS=S:RQ"1v up"R;S-1-R0MsHo5RR#bHlDRC,8NCD$b,RECN#_8NM_D8CNR$,CCG0sDMN2SR
Sp7 qqY_71Kzahv am_v7w _ A 7qRBiR#:R0MsHoSRSSR:="XwQ ;7"RS
S7q pY7_qKaz1va h_7vm  _)pQqaeS R:0R#soHMS:SS=wR"Q7X "
;RS]S1Q)wa 7t_Qve_mR7 SRS:L_H0P0COF4s5RI8FMR0Fj:2S=jR"jR";S-R-R-Rj-H>7PCH8RRL$c4,R-7->H8PHC$RLRR(,d-R->P7HHR8CL6$RSS
Sw_7qw7  AiqBRSSS:HRL0C_POs0F58dRF0IMF2RjR=S:Rj"jj;j"R-SR-QRRMo0CC5sRj6-42
3RS7Swq _)pQqaeS RSRS:L_H0P0COFds5RI8FMR0Fj:2S=jR"j"jj;RRS-R-RQCM0oRCs54j-6R23RSR
Spupm_za1  pBua_mq)aSRS:#H0sMSoRS=S:R "thiBp"R;R
uSSpzpma _1pa B_)umaSAS:0R#soHMRSSS:"=RtB hp;i"RSR
Se7Q)SRSSRS:L_H0P0COFds5RI8FMR0Fj:2S=jR"j"jj;
RSSQS7eSwRS:SSR0LH_OPC05FsnFR8IFM0RRj2SR:="jjjjjjj"
;RSQS7eSTRS:SSR0LH_OPC05Fs.FR8IFM0RSj2:"=Rj"jj;SRS
wSSQ pa)q_)hRt S:SSR0LH_OPC05Fs.FR8IFM0RRj2RRRRR:RR=jR"j;j"RSS
Sq hA_p QtB q_a uam)q:SSR0LHSSSS:'=Rj
';ShS q Ap_ QBt qa_)umaSAS:HRL0SSSSR:=';j'
aSS _1av m7RSSS:HRL0SSSSR:=';j'
 SSX)a h_qp7QQe7w _qmBa)SRS:MRH0CCosSSS:4=RRRSS-F-h0#RkCL8R$FRl83CDR8q8CV8RFusRpBpRFHMVozRtQR3
S;R2
b
SFRs0SS5
RRRRRSRRuiqBqut QShSSH:RM0FkR8#0_oDFH;ORR-SS-CR)VCCsMROCORD	5Ru2#MHoN0DREksFouERNNO	oHCuMR3RRR
SRRRRRuRSqqBitQ uhSASSH:RM0FkR8#0_oDFH;ORR-SS-CR)VCCsMROCORD	5Rh2#MHoN0DREksFouERNNO	oHCuMRA3RSR
SpupmBzamq) S:SSR0FkR8#0_oDFHRO;S-S-RpupRbqRFRs0Fbk0k00RFFROsDCRFOoHR$5LRsMFlRNDs0FkH2Mo
uSSpzpmamtpAqqpSRRRSRS:FRk0#_08DHFoOS;RSR--uRppqFRbsF0Rkk0b0FR0RsOFCFRDoRHO5RL$oLDFNsDRFHk0M
o2SRRRRRRRRpupmBzamA) S:SSR0FkR8#0_oDFHRO;S-S-RpupRbARFRs0Fbk0k00RFFROsDCRFOoHR$5LRsMFlRNDs0FkH2Mo
uSSpzpmamtpAAqpSRRRSRS:FRk0#_08DHFoOS;RSR--uRppAFRbsF0Rkk0b0FR0RsOFCFRDoRHO5RL$oLDFNsDRFHk0M
o2SXS a w 7BAqiSRRSRS:H#MR0D8_FOoH;SSS-7-RsCHPM$RLRsOFCFRDo
HOSYS7hQqvBp7 qSYSSH:RM0R#8F_Do_HOP0COF5sR(FR8IFM0R;j2SR--7PsHCLMR$FROsDCRFOoH
pSSmSBiS:SSR0FkR8#0_oDFHRO;S-S-R0mkbRk0FuVRpSp
SuAYqS11S:SSRRHM#_08DHFoOS;RSR--7PsHCLMR$FROsDCRFOoH
)SS a1 ASSSSH:RM0R#8F_Do;HOR-SS-sR7HMPCRRL$OCFsRoDFHSO
SQ17SSSS:MRHR8#0_oDFHRO;S-S-RH7sPRCMLO$RFRsCDHFoOa3RCR#0u
HMS7S1mSSSSF:Rk#0R0D8_FOoH;-SS-kRm00bkRR0F)pARFOoHRDaHCa3RCR#0u
HMSBS1pSiSSRS:H#MR0D8_FOoH;SRS-7-RsCHPM$RLRsOFCFRDo3HOR#aC0HRuMS
SpBqa]uQhzqaepRz SRS:H#MR0D8_FOoHRSSS-H-RBN t0#CRHNoMDSS
RRRRR2RR;CR
MO8RFFlbM0CM;
RS
R--HcB jQRvuuQRsHHl0CHPR-R
--------------------------------------------------------------------------------------------------
-RSSSSAS1_uvQQX_)_q.phS SS-SS--
-------------------------------------------------------------------------------------------------
F
OlMbFCRM01vA_Q_uQ).X_p qhRSR
b0FsRS5
Su h7  1)SRRSH:RM0R#8F_Do;HORRSRS-S-RlBFlRFMQCM0sOVNCHRuM
#RRSRSuSzSSH:RM0R#8F_Do;HORRSR
7SSuSjSSH:RM0R#8F_Do;HORRSRS-S-RP7CHROCuRHM
7SShSjSSH:RM0R#8F_Do;HORRSRSRRRRRRRRR--7HCPOuCRH
MRSjS7)1X] ShS:MRHR8#0_oDFHRO;SRRRS-S-R07NNQjRMs0CVCNORMuH#SR
S77jauXpu:SSRRHM#_08DHFoOS;RR
RRSjS77paXuShS:MRHR8#0_oDFHRO;S
RRSjS7auXp ShS:MRHR8#0_oDFHRO;SRRRSS
S7)j7XupuSRS:FRk0#_08DHFoOS;RR
RRSjS77p)XuShS:kRF00R#8F_Do;HORSR
S)7jX puh:SSRRHM#_08DHFoOS;RRSR
S77jBS7uSRS:FRk0#_08DHFoOR;RSSR
S77jBR7hS:SSR0FkR8#0_oDFHRO;R
SRSjS7Bh7 S:SSRRHM#_08DHFoO
;RSjS7] 171  )h:SSRRHM#_08DHFoO
;RSjS7]X1)7qqaSRS:FRk0#_08DHFoOC_POs0F58(RF0IMF2Rj;RR
SjS7]Y1Aap BiS7S:kRF00R#8F_Do;HORSS
S17jYShBSRS:FRk0#_08DHFoOR;R
7SSj) )1BYhSRS:FRk0#_08DHFoO
;RSjS7hYm1hSBS:kRF00R#8F_Do;HORS
S7Su4SRS:H#MR0D8_FOoH;SRRS-S-RP7CHROCuRHM
7SShS4SSH:RM0R#8F_Do;HORSSS-7-RCOPHCHRuMSR
S)74X ]1h:SSRRHM#_08DHFoOS;RS-S-R07NNQ4RMs0CVCNORMuH#SR
S774)uXpu:SSR0FkR8#0_oDFHRO;
7SS4X7)pSuhSF:Rk#0R0D8_FOoH;
RSS4S7)uXp ShS:MRHR8#0_oDFHRO;
7SS47]1 )1  ShS:MRHR8#0_oDFHRO;
7SS4)]1Xa7qq:SSR0FkR8#0_oDFHPO_CFO0sR5(8MFI0jFR2
;RS4S71BYhS:SSR0FkR8#0_oDFHRO;
7SS4) )1BYhSRS:FRk0#_08DHFoO
;RS4S7hYm1hSBS:kRF00R#8F_Do;HORS
SBSiuSRS:H#MR0D8_FOoH;RRRRRRRRSRRSR--7HCPOuCRHRMRRS
SBSihSRS:H#MR0D8_FOoH;SSSSR--7HCPOuCRH
MRSpSBi])X1S hSH:RM0R#8F_Do;HORSSRSR--BRD	HCM0sOVNCHRuMR#R
BSSp)i7XupuSRS:FRk0#_08DHFoOS;R
BSSp)i7XhpuSRS:FRk0#_08DHFoOS;R
BSSpXi)phu SRS:H#MR0D8_FOoH;
RSSpSBiA]1YSa SF:Rk#0R0D8_FOoHRR
RRRRRSRRRR;R2RM
C8FROlMbFC;M0R-

-BRH Rcj]Q7vRHuslHH0PRCR
------------------------------------------------------------------------------------------------
---S-RSSSS1aA_v_718CC#sDHNHsxCSSSSS
---------------------------------------------------------------------------------------------------
-
ObFlFMMC0AR1_7av1C_8#HCsNxDHCRsR
CSoMHCsO
R5S Sw q7ABui_qRa]S:SSRs#0HRMoS:SS=uR"] q1_7qh_p7 q;Y"SSR
Sp7 qqY_71Kzahv am_v7w _ A 7qRBiR#:R0MsHoSRSSR:="XwQ ;7"RS
S7q pY7_qKaz1va h_7vm  _)pQqaeS R:0R#soHMS:SS=wR"Q7X "
;RS]S1Q)wa 7t_Qve_mR7 SRS:L_H0P0COF4s5RI8FMR0Fj:2S=4R"4R";S-R-RHR7PCH8RRL$6FRl8SCR
wSS7wq_ A 7qRBiS:SSR0LH_OPC05FsdFR8IFM0RRj2SR:="jjjjR";S-R-RMRQ0CCosjR5-2463SR
Sqw7_p) qeaQ SRSSL:RHP0_CFO0sR5d8MFI0jFR2=S:Rj"jj;j"R-SR-QRRMo0CC5sRj6-42R3RRS
Sumppz1a_ Bp am_u)SaqS#:R0MsHoSRSSR:="ht B"pi;RRS-R-RBGD	6S
Sumppz1a_ Bp am_u)SaAS#:R0MsHoSRSSR:="Q1]w a)t8_jC;o"R-R-R	BDGR4R
7SSQRe)SSSS:HRL0C_POs0F58dRF0IMF2RjSR:="jjjjR";SRRRRR--VRFsa1v7R	ODRRN0cEjvxSRR
7SSQRewSSSS:HRL0C_POs0F58nRF0IMF2RjR=S:Rj"jjjjjjR";
7SSQReTSSSS:HRL0C_POs0F58.RF0IMF2RjSR:="jj4"S;RSS
SwaQp ))_q htRSSS:HRL0C_POs0F58.RF0IMF2RjRRRRRRRR:"=Rj"44;
RSShS q Ap_ QBt qa_)umaSqS:HRL0SSSSR:=';j'
 SShpqA B_Q atq m_u)SaASL:RHS0SS=S:R''j;S
Saa 1_7vm SRSSL:RHS0SS=S:R''j;S
S  Xa)phq_e7QQ_7 waqBmS)RSH:RMo0CCSsSSR:=4SRSRh--Fk0R#RC8Ll$RFD8C38Rq8RC8VRFsuRppBVFMHtoRz
Q3
SSR2
;RSsbF05RS
aSSvO71ERjbS:SSRRHM#_08DHFoOS;SRSRRRRRRR-S-a1v7RROEjHR8VsVCCHM0NHDRM0bkR#bF
aSSvO71ESjMSRS:H#MR0D8_FOoH;RRRRRRRRSRS-v-a7O1RERRj8VHVCMsC0DHNRbHMkM0RCSo
S7av14OEbSSS:MRHR8#0_oDFHRO;RRRRRRRRRRRRR-SS-7av1EROR84RHCVVs0CMHRNDHkMb0FRb#S
Sa1v7OME4S:SSRRHM#_08DHFoOR;RRRRRRRRRRRRRS-S-a1v7RROE4HR8VsVCCHM0NHDRM0bkRoMC
aSSvO71ES.bSRS:H#MR0D8_FOoH;RRRRRRRRRRRRSRRSa--vR71O.ERRV8HVCCsMN0HDMRHbRk0b
F#SvSa7E1O.SMSSH:RM0R#8F_Do;HORRRRRRRRRRRRRSRS-v-a7O1RERR.8VHVCMsC0DHNRbHMkM0RCSo
S7av1	ODbSSS:MRHR8#0_oDFHRO;RRRRRRRRRRRRR-SS-7av1DROFRO	8VHVCMsC0DHNRbHMkb0RFS#
S7av1	ODMSSS:MRHR8#0_oDFHRO;RRRRRRRRRRRRR-SS-7av1DROFRO	8VHVCMsC0DHNRbHMkM0RCSo
SSSSSRSSRRRRRRRRRRRRRRRRRRRRR-RR-O)CCCHPsFROMF0sDsDCR0HMCNsVOSC
Sa)1h#8CCSsSSH:RM0R#8F_Do;HOSSSS-C-)#RC08CC#sDNHxsHCRoDFH-O#R0NOHRPCD
FIS1S)aDhbDSSSSH:RM0R#8F_Do;HORRRRRRRRRRRRRRRRS-S-)CC#0CR8#HCsNxDHCusRpRp-NHO0PDCRFSI
SS hS:SSRRHM#_08DHFoOR;RRRRRRRRRRRRRRRRRRRRRS --MDNLCCR8#HCsNxDHCRs-NHO0PECRH
oES]Suqp1 OREjS:SSRRHM#_08DHFoOC_POs0F58dRF0IMF2Rj;RRRR-RR-FBDOb	RECN#RD8CNO$RFClbM0#NHRFM#CCDOV0RFOsRE
RjS]Suqp1 ORE4S:SSRRHM#_08DHFoOC_POs0F58dRF0IMF2Rj;RRRR-RR-FBDOb	RECN#RD8CNO$RFClbM0#NHRFM#CCDOV0RFOsRE
R4S]Suqp1 ORE.S:SSRRHM#_08DHFoOC_POs0F58dRF0IMF2Rj;RRRR-RR-FBDOb	RECN#RD8CNO$RFClbM0#NHRFM#CCDOV0RFOsRE
R.SpSupODF	SSSSF:Rk#0R0D8_FOoH;RRRRRRRRRRRRRRRS-S-RpupRODF	HR#oDMN-ORN0CHPRoEHES
SSSSSSSSSSR--uRppFbk0kR0R
uSSpzpma)Bm 	ODGR4RSRS:FRk0#_08DHFoOS;RS-S-RpupRR4GFbk0kF0RMFROsMCRCF0IsR	R
uSSpzpmamtpAOqpD4	GR:SSR0FkR8#0_oDFH;ORRSSS-u-Rp4pRGkRF00bkRRFMoLDFNMDRCF0IsS	R
uSSpzpma)Bm 	ODGS6SSF:Rk#0R0D8_FOoHRS;RS-S-RpupRR6GFbk0kF0RMFROsMCRCF0Is
	RSpSupamztApmqDpO	RG6SRS:FRk0#_08DHFoORR;S-SS-pRupGR6R0FkbRk0FoMRDNFLDCRM0sIF	
RRSqS)Wa7qqjOERSRSSF:Rk#0R0D8_FOoH_OPC05FsgFR8IFM0R;j2R-S-RO)CFsPCCO8RERRj4Lj-H80RNR0N
)SSqqW7aEqO4SRRSRS:FRk0#_08DHFoOC_POs0F58gRF0IMF2Rj;-RS-CR)OCFPsRC8O4ERR-4jLRH08NN0
)SSqqW7aEqO.RRRS:SSR0FkR8#0_oDFHPO_CFO0sR5g8MFI0jFR2S;R-)-RCPOFC8sCRROE.jR4-0LHR08NNS
S wXa A 7qSBiRSRRSH:RM0R#8F_DoRHO;SRSSR--7PsHCLMR$FROsDCRFOoH3FRh0CRsJskHC]8R7RvQlCF83S
S7qYhv7QB YpqRSSS:MRHR8#0_oDFHPO_CFO0sR5(8MFI0jFR2R;RSR--7PsHCLMR$FROsDCRFOoH3FRh0CRsJskHCV8RF]sR7RvQlCF83S
SAqYu1S1SSRS:H#MR0D8_FOoHRS;RS-S-RH7sPRCMLO$RFRsCDHFoOh3RFs0RCHJksRC8VRFs]Q7vR8lFCS3
SapqBh]Quezaq pzR:SSRRHM#_08DHFoORR;S-SS-BRH 0tNCHR#oDMN3FRh0CRsJskHCV8RF]sR7RvQlCF8
SSSSSSSSSSS-a-RCR#0u#HMRSS
Sm17SSSS:kRF00R#8F_Do;HORSRSSR--a0C#Ro1HM3NDR0mkbRk0FuVRp
p3S7S1QSSSSH:RM0R#8F_DoRHO;SRSSR--a0C#Ro#HM3NDRH7sPRCMLO$RFRsCDHFoOS
S1iBpSSSS:MRHR8#0_oDFHRORS-SS-CRa#B0RD1	RHNoMD73RsCHPM$RLRsOFCFRDo
HORRRRRSRRSR2;
8CMRlOFbCFMM
0;
---------------------------------------------
-RQu)vYRauR R:vRRzQpau pQ)
1R-7-R BeQ RRRRRR:R QBc1jRq)hwh1BQB7mR BeQ -1
-------------------------------------------
-----------------------------------------
---S-RS_1Avazp_UUGR-
------------------------------------------O-
FFlbM0CMR_1Avazp_UUG
CSoMHCsORR5
7SSqqaq_t) SL:RHR0RSR:=';j'SS
S7qqaA _)t:RSR0LHSR:=';j'SS
S7qqam_za)R tSL:RHS0R:'=Rj
';SqS7a_qq1hQt S7R:HRL0SRR:'=Rj
';SqS7a_qA1hQt S7R:HRL0SRR:'=Rj
';S Sht)_aQ tt)SRR:HRL0:RS=jR''RR
RRRRRRRRRRRRR;R2Rb
SFRs0R
R5SqS7aRqqRRR:H#MR0D8_FOoH_OPC05FsR8(RF0IMF2Rj;SR
Sa7qqRARRH:RM0R#8F_Do_HOP0COFRs5(FR8IFM0R;j2RS
SBRpiRRRR:MRHR8#0_oDFHRO;RS
SBR RRRRR:MRHR8#0_oDFHRO;RS
S)  1aRRR:MRHR8#0_oDFHRO;RRRRRRRRRRRRRRRRRRRRR-R-R$q#MsOEFkMF#CR)#
C0R7SSqmaqz:aRR0FkR8#0_oDFHPO_CFO0s654RI8FMR0FjS2
2S;R
8CMRlOFbCFMMR0;S-

--------------------------------------------
R--SAS1_pvzan_4GR4n
--------------------------------------------O-
FFlbM0CMR_1Avazp_G4n4Sn
oCCMsRHO5SR
Sa7qq)q_ :tSR0LHR:RS=jR''
;SSqS7a_qA)R tSL:RH:0S=jR''S;
SuuQ hpQ  _)tRS:LSH0:'=Rj
';SqS7azqma _)t:RSR0LHR=S:R''j;S
S7qqaqQ_1t7h RRS:LRH0R=S:R''j;S
S7qqaAQ_1t7h RRS:LRH0R=S:R''j;S
Sh_ tat)QtR )RRS:LRH0SR:='Rj'
RRRRRRRRRRRRRRR2
;RSsbF0RRR5S
S7qqaqRRR:MRHR8#0_oDFHPO_CFO0s45R6FR8IFM0R;j2RS
S7qqaARRR:MRHR8#0_oDFHPO_CFO0s45R6FR8IFM0R;j2RS
SBRpiRRRR:MRHR8#0_oDFHRO;
BSS RRRR:RRRRHM#_08DHFoOR;R
)SS a1 R:RRRRHM#_08DHFoOR;RRRRRRRRRRRRRRRRRRRRRRR--qM#$OFEsM#FkR#)CC
0RR7SSqmaqz:aRR0FkR8#0_oDFHPO_CFO0s45dRI8FMR0FjS2
2S;R
8CMRlOFbCFMM
0;ObFlFMMC0AR1_v)qc4j_n
iRRCRoMHCsORR5
RSRRQW)av _mR7 :MRH0CCos=R:RRj;
RSRRq) 7m_v7R R:MRH0CCos=R:RRj;
R
SRhRQQja_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRhRQQ4a_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRhRQQ.a_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRhRQQda_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRhRQQca_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRhRQQ6a_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRhRQQna_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRhRQQ(a_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRhRQQUa_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRhRQQga_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRhRQQqa_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRhRQQAa_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRhRQQBa_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRhRQQ7a_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRhRQQ a_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRhRQQwa_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;
R
RRRRRRRRRQRRh_Qa4:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjR";
R
RRRRRRRRRRQQhaj_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha4_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha._.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhad_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhac_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha6_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhan_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha(_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaU_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhag_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaq_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaA_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaB_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha7_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha _.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaw_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;
R
RRRRRRRRRQRRh_Qad:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
"RSRRRR;2R
RSRb0Fs5SR
Sq)7a:qRR0FkR8#0_oDFHPO_CFO0s45R68RRF0IMF2RjRS;
Sp)Bi:RRRRHMR8#0_oDFH;OR
)SSB piRH:RM#RR0D8_FOoHRR:=';]'
)SS RRRRH:RM#RR0D8_FOoHRR:=';]'
)SSq)77RH:RM#RR0D8_FOoH_OPC05FsRR4.RI8FMR0Fj;2R
WSSBRpiRH:RM#RR0D8_FOoHRS;
SpWBi: RRRHMR8#0_oDFH:OR=]R''S;
SRW R:RRRRHMR8#0_oDFH:OR=]R''S;
S7Wq7:)RRRHMR8#0_oDFHPO_CFO0s45R.8RRF0IMF2RjRS;
S1vqi:RRRRHMR8#0_oDFHPO_CFO0s45R68RRF0IMF2RjRS;
SqW7a:qRRRHMR8#0_oDFHPO_CFO0s45R68RRF0IMF2Rj
RSRRRRRR
2;S
RRCRM8ObFlFMMC0
;
ObFlFMMC0AR1_v)qc4j_n)ihR
H#RCRoMHCsORR5
RSRRQW)av _mR7 :MRH0CCos=R:RRj;
RRRRRRRRRRR)7 q_7vm :RRR0HMCsoCRR:=j
;R
RSRRQQhaR_j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRQQhaR_4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRQQhaR_.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRQQhaR_d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRQQhaR_c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRQQhaR_6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRQQhaR_n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRQQhaR_(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRQQhaR_U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRQQhaR_g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRQQhaR_q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRQQhaR_A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRQQhaR_B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRQQhaR_7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRQQhaR_ :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRQQhaR_w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"RR

RRRRRRRRRhRQQ4a_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
RRRRRRRRRQRRh_Qa.:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa.:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa.:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa.:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa.:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa.:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa.:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa.:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa.:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa.:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa.:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa.:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa.:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa.:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa.: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa.:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RRRRRRRRRRRQahQ_Rdj:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_Rd4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_Rd.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_Rdd:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_Rdc:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_Rd6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_Rdn:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_Rd(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_RdU:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_Rdg:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_Rdq:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_RdA:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_RdB:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_Rd7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_Rd :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_Rdw:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjRj"
RSRRRR2;R
SRsbF0
5RS7S)qRaq:kRF00R#8F_Do_HOP0COFRs54R6R8MFI0jFR2
R;SBS)pRih:MRHR0R#8F_DoRHO;S
S)iBp RR:HRMR#_08DHFoO=R:R''];S
S)R RRRR:HRMR#_08DHFoO=R:R''];S
S)7q7)RR:HRMR#_08DHFoOC_POs0F5.R4RFR8IFM0RRj2;S
SWiBpRRR:HRMR#_08DHFoO
R;SBSWpRi :MRHR0R#8F_DoRHO:'=R]
';S SWRRRR:MRHR0R#8F_DoRHO:'=R]
';SqSW7R7):MRHR0R#8F_Do_HOP0COFRs54R.R8MFI0jFR2
R;SqSv1RiR:MRHR0R#8F_Do_HOP0COFRs54R6R8MFI0jFR2
R;S7SWqRaq:MRHR0R#8F_Do_HOP0COFRs54R6R8MFI0jFR2R
SRRRRR;R2
8CMRlOFbCFMM
0;
lOFbCFMM10RAq_)v_cj4hniW#RH
oRRCsMCH5ORRR
SR)RWQ_a v m7RH:RMo0CC:sR=;RjRR
SR R)qv7_mR7 RH:RMo0CC:sR=;RjRS

RQRRh_QajRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_Qa4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_Qa.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_QadRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_QacRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_Qa6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_QanRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_Qa(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_QaURR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_QagRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_QaqRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_QaARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_QaBRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_Qa7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_Qa RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_QawRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
RRRRRRRRRQRRh_Qa4:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RRRRRRRRRRRQahQ_R.j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R..:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R. :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
RRRRRRRRRRQQhaj_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha4_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha._dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhad_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhac_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha6_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhan_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha(_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaU_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhag_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaq_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaA_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaB_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha7_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha _dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaw_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jjRR
SR2RRRS;
RFRbsR05
)SS7qqaRF:Rk#0R0D8_FOoH_OPC05FsRR46RI8FMR0Fj;2R
)SSBRpiRH:RM#RR0D8_FOoHRS;
Sp)Bi: RRRHMR8#0_oDFH:OR=]R''S;
SR) R:RRRRHMR8#0_oDFH:OR=]R''S;
S7)q7:)RRRHMR8#0_oDFHPO_CFO0s45R.8RRF0IMF2RjRS;
SpWBi:hRRRHMR8#0_oDFH;OR
WSSB piRH:RM#RR0D8_FOoHRR:=';]'
WSS RRRRH:RM#RR0D8_FOoHRR:=';]'
WSSq)77RH:RM#RR0D8_FOoH_OPC05FsRR4.RI8FMR0Fj;2R
vSSqR1iRH:RM#RR0D8_FOoH_OPC05FsRR46RI8FMR0Fj;2R
WSS7qqaRH:RM#RR0D8_FOoH_OPC05FsRR46RI8FMR0FjS2
RRRRR2RR;M
C8FROlMbFC;M0
F
OlMbFCRM01)A_qjvc_i4nhW)hR
H#RCRoMHCsORR5
RSRRQW)av _mR7 :MRH0CCos=R:RRj;
RRRRRRRRRRR)7 q_7vm :RRR0HMCsoCRR:=j
;R
RSRRQQhaR_j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRQQhaR_4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRQQhaR_.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRQQhaR_d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRQQhaR_c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRQQhaR_6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRQQhaR_n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRQQhaR_(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRQQhaR_U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRQQhaR_g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRQQhaR_q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRQQhaR_A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRQQhaR_B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRQQhaR_7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRQQhaR_ :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRQQhaR_w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
RRRRRRRRRRQQhaj_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha4_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha._4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhad_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhac_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha6_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhan_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha(_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaU_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhag_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaq_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaA_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaB_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha7_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha _4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaw_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R

RRRRRRRRRhRQQ.a_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
RRRRRRRRRQRRh_Qad:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
"RRRRRRRRRR2RRRS;
RFRbsR05
)SS7qqaRF:Rk#0R0D8_FOoH_OPC05FsRR46RI8FMR0Fj;2R
)SSBhpiRH:RM#RR0D8_FOoHRS;
Sp)Bi: RRRHMR8#0_oDFH:OR=]R''S;
SR) R:RRRRHMR8#0_oDFH:OR=]R''S;
S7)q7:)RRRHMR8#0_oDFHPO_CFO0s45R.8RRF0IMF2RjRS;
SpWBi:hRRRHMR8#0_oDFH;OR
WSSB piRH:RM#RR0D8_FOoHRR:=';]'
WSS RRRRH:RM#RR0D8_FOoHRR:=';]'
WSSq)77RH:RM#RR0D8_FOoH_OPC05FsRR4.RI8FMR0Fj;2R
vSSqR1iRH:RM#RR0D8_FOoH_OPC05FsRR46RI8FMR0Fj;2R
WSS7qqaRH:RM#RR0D8_FOoH_OPC05FsRR46RI8FMR0FjS2
RRRRR2RR;M
C8FROlMbFC;M0
F
OlMbFCRM01)A_qjv4.4cGnRR
RMoCCOsHR
5RSRRRQahQ_:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RRRRRRRRRRRQahQ_R4j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R44:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R46:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R47:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4 :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
RRRRRRRRRRQQhaj_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha4_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha._.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhad_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhac_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha6_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhan_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha(_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaU_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhag_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaq_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaA_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaB_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha7_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha _.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaw_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R

RRRRRRRRRhRQQda_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"SR
RRRR2
R;SbRRF5s0RS
S)a7qqRR:FRk0#_08DHFoOC_POs0F56R4RFR8IFM0RRj2;S
S)iBpRRR:HRMR#_08DHFoO
R;SBS)pRi :MRHR0R#8F_DoRHO:'=R]
';S S)RRRR:MRHR0R#8F_DoRHO:'=R]
';SqS)7R7):MRHR0R#8F_Do_HOP0COFRs5g8RRF0IMF2RjRS;
SpWBi:RRRRHMR8#0_oDFH;OR
WSSB piRH:RM#RR0D8_FOoHRR:=';]'
WSS RRRRH:RM#RR0D8_FOoHRR:=';]'
WSSq)77RH:RM#RR0D8_FOoH_OPC05FsRRgR8MFI0jFR2
R;SqSv1RiR:MRHR0R#8F_Do_HOP0COFRs54R6R8MFI0jFR2
R;S7SWqRaq:MRHR0R#8F_Do_HOP0COFRs54R6R8MFI0jFR2R
SRRRRR;R2
RSR
8CMRlOFbCFMM
0;
lOFbCFMM10RAq_)v.4jcnG4hH)R#R
RoCCMsRHO5SR
RQRRh_QajRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_Qa4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_Qa.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_QadRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_QacRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_Qa6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_QanRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_Qa(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_QaURR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_QagRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_QaqRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_QaARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_QaBRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_Qa7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_Qa RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_QawRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
RRRRRRRRRQRRh_Qa4:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RRRRRRRRRRRQahQ_R.j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R..:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R. :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
RRRRRRRRRRQQhaj_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha4_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha._dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhad_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhac_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha6_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhan_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha(_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaU_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhag_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaq_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaA_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaB_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha7_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha _dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaw_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jjRR
SR2RRRS;
RFRbsR05
)SS7qqaRF:Rk#0R0D8_FOoH_OPC05FsRR46RI8FMR0Fj;2R
)SSBhpiRH:RM#RR0D8_FOoHRS;
Sp)Bi: RRRHMR8#0_oDFH:OR=]R''S;
SR) R:RRRRHMR8#0_oDFH:OR=]R''S;
S7)q7:)RRRHMR8#0_oDFHPO_CFO0sg5RRFR8IFM0RRj2;S
SWiBpRRR:HRMR#_08DHFoO
R;SBSWpRi :MRHR0R#8F_DoRHO:'=R]
';S SWRRRR:MRHR0R#8F_DoRHO:'=R]
';SqSW7R7):MRHR0R#8F_Do_HOP0COFRs5g8RRF0IMF2RjRS;
S1vqi:RRRRHMR8#0_oDFHPO_CFO0s45R68RRF0IMF2RjRS;
SqW7a:qRRRHMR8#0_oDFHPO_CFO0s45R68RRF0IMF2Rj
RSRRRRRR
2;CRM8ObFlFMMC0
;
ObFlFMMC0AR1_v)q4cj.Gh4nW#RH
oRRCsMCH5ORRR
SRhRQQja_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRhRQQ4a_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRhRQQ.a_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRhRQQda_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRhRQQca_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRhRQQ6a_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRhRQQna_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRhRQQ(a_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRhRQQUa_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRhRQQga_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRhRQQqa_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRhRQQAa_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRhRQQBa_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRhRQQ7a_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRhRQQ a_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRhRQQwa_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R

RRRRRRRRRhRQQ4a_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
RRRRRRRRRQRRh_Qa.:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa.:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa.:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa.:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa.:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa.:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa.:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa.:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa.:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa.:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa.:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa.:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa.:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa.:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa.: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa.:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RRRRRRRRRRRQahQ_Rdj:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_Rd4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_Rd.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_Rdd:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_Rdc:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_Rd6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_Rdn:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_Rd(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_RdU:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_Rdg:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_Rdq:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_RdA:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_RdB:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_Rd7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_Rd :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_Rdw:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjRj"
RSRRRR2;R
SRsbF0
5RS7S)qRaq:kRF00R#8F_Do_HOP0COFRs54R6R8MFI0jFR2
R;SBS)pRiR:MRHR0R#8F_DoRHO;S
S)iBp RR:HRMR#_08DHFoO=R:R''];S
S)R RRRR:HRMR#_08DHFoO=R:R''];S
S)7q7)RR:HRMR#_08DHFoOC_POs0F5RRgRI8FMR0Fj;2R
WSSBhpiRH:RM#RR0D8_FOoHRS;
SpWBi: RRRHMR8#0_oDFH:OR=]R''S;
SRW R:RRRRHMR8#0_oDFH:OR=]R''S;
S7Wq7:)RRRHMR8#0_oDFHPO_CFO0sg5RRFR8IFM0RRj2;S
Sviq1RRR:HRMR#_08DHFoOC_POs0F56R4RFR8IFM0RRj2;S
SWa7qqRR:HRMR#_08DHFoOC_POs0F56R4RFR8IFM0R
j2SRRRRRRR2C;
MO8RFFlbM0CM;O

FFlbM0CMR_1A)4qvjG.c4)nhhHWR#R
RoCCMsRHO5SR
RQRRh_QajRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_Qa4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_Qa.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_QadRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_QacRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_Qa6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_QanRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_Qa(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_QaURR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_QagRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_QaqRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_QaARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_QaBRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_Qa7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_Qa RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_QawRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
RRRRRRRRRQRRh_Qa4:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RRRRRRRRRRRQahQ_R.j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R..:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R. :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
RRRRRRRRRRQQhaj_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha4_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha._dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhad_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhac_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha6_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhan_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha(_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaU_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhag_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaq_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaA_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaB_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha7_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha _dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaw_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jjRR
SR2RRRS;
RFRbsR05
)SS7qqaRF:Rk#0R0D8_FOoH_OPC05FsRR46RI8FMR0Fj;2R
)SSBhpiRH:RM#RR0D8_FOoHRS;
Sp)Bi: RRRHMR8#0_oDFH:OR=]R''S;
SR) R:RRRRHMR8#0_oDFH:OR=]R''S;
S7)q7:)RRRHMR8#0_oDFHPO_CFO0sg5RRFR8IFM0RRj2;S
SWiBphRR:HRMR#_08DHFoO
R;SBSWpRi :MRHR0R#8F_DoRHO:'=R]
';S SWRRRR:MRHR0R#8F_DoRHO:'=R]
';SqSW7R7):MRHR0R#8F_Do_HOP0COFRs5g8RRF0IMF2RjRS;
S1vqi:RRRRHMR8#0_oDFHPO_CFO0s45R68RRF0IMF2RjRS;
SqW7a:qRRRHMR8#0_oDFHPO_CFO0s45R68RRF0IMF2Rj
RSRRRRRR
2;CRM8ObFlFMMC0
;
ObFlFMMC0AR1_v)q.UjcGHUR#R
RoCCMsRHO5SR
RQRRh_QajRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_Qa4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_Qa.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_QadRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_QacRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_Qa6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_QanRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_Qa(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_QaURR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_QagRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_QaqRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_QaARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_QaBRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_Qa7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_Qa RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_QawRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
RRRRRRRRRQRRh_Qa4:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RRRRRRRRRRRQahQ_R.j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R..:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R. :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
RRRRRRRRRRQQhaj_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha4_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha._dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhad_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhac_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha6_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhan_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha(_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaU_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhag_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaq_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaA_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaB_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha7_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha _dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaw_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jjRR
SR2RRRS;
RFRbsR05
)SS7qqaRF:Rk#0R0D8_FOoH_OPC05FsRR(R8MFI0jFR2
R;SBS)pRiR:MRHR0R#8F_DoRHO;S
S)iBp RR:HRMR#_08DHFoO=R:R''];S
S)R RRRR:HRMR#_08DHFoO=R:R''];S
S)7q7)RR:HRMR#_08DHFoOC_POs0F5jR4RFR8IFM0RRj2;S
SWiBpRRR:HRMR#_08DHFoO
R;SBSWpRi :MRHR0R#8F_DoRHO:'=R]
';S SWRRRR:MRHR0R#8F_DoRHO:'=R]
';SqSW7R7):MRHR0R#8F_Do_HOP0COFRs54RjR8MFI0jFR2
R;S7SWqRaq:MRHR0R#8F_Do_HOP0COFRs5(8RRF0IMF2Rj
RSRRRRRR
2;CRM8ObFlFMMC0
;
ObFlFMMC0AR1_v)q.UjcG)UhR
H#RCRoMHCsORR5
RSRRQQhaR_j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRQQhaR_4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRQQhaR_.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRQQhaR_d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRQQhaR_c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRQQhaR_6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRQQhaR_n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRQQhaR_(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRQQhaR_U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRQQhaR_g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRQQhaR_q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRQQhaR_A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRQQhaR_B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRQQhaR_7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRQQhaR_ :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRQQhaR_w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
RRRRRRRRRRQQhaj_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha4_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha._4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhad_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhac_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha6_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhan_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha(_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaU_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhag_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaq_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaA_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaB_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha7_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha _4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaw_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R

RRRRRRRRRhRQQ.a_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
RRRRRRRRRQRRh_Qad:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
"RSRRRR;2R
RSRb0Fs5SR
Sq)7a:qRR0FkR8#0_oDFHPO_CFO0s(5RRFR8IFM0RRj2;S
S)iBphRR:HRMR#_08DHFoO
R;SBS)pRi :MRHR0R#8F_DoRHO:'=R]
';S S)RRRR:MRHR0R#8F_DoRHO:'=R]
';SqS)7R7):MRHR0R#8F_Do_HOP0COFRs54RjR8MFI0jFR2
R;SBSWpRiR:MRHR0R#8F_DoRHO;S
SWiBp RR:HRMR#_08DHFoO=R:R''];S
SWR RRRR:HRMR#_08DHFoO=R:R''];S
SW7q7)RR:HRMR#_08DHFoOC_POs0F5jR4RFR8IFM0RRj2;S
SWa7qqRR:HRMR#_08DHFoOC_POs0F5RR(RI8FMR0FjS2
RRRRR2RR;M
C8FROlMbFC;M0
F
OlMbFCRM01)A_qjv.cUUGhHWR#R
RoCCMsRHO5SR
RQRRh_QajRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_Qa4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_Qa.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_QadRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_QacRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_Qa6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_QanRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_Qa(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_QaURR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_QagRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_QaqRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_QaARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_QaBRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_Qa7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_Qa RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_QawRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
RRRRRRRRRQRRh_Qa4:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RRRRRRRRRRRQahQ_R.j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R..:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R. :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
RRRRRRRRRRQQhaj_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha4_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha._dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhad_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhac_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha6_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhan_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha(_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaU_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhag_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaq_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaA_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaB_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha7_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha _dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaw_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jjRR
SR2RRRS;
RFRbsR05
)SS7qqaRF:Rk#0R0D8_FOoH_OPC05FsRR(R8MFI0jFR2
R;SBS)pRiR:MRHR0R#8F_DoRHO;S
S)iBp RR:HRMR#_08DHFoO=R:R''];S
S)R RRRR:HRMR#_08DHFoO=R:R''];S
S)7q7)RR:HRMR#_08DHFoOC_POs0F5jR4RFR8IFM0RRj2;S
SWiBphRR:HRMR#_08DHFoO
R;SBSWpRi :MRHR0R#8F_DoRHO:'=R]
';S SWRRRR:MRHR0R#8F_DoRHO:'=R]
';SqSW7R7):MRHR0R#8F_Do_HOP0COFRs54RjR8MFI0jFR2
R;S7SWqRaq:MRHR0R#8F_Do_HOP0COFRs5(8RRF0IMF2Rj
RSRRRRRR
2;CRM8ObFlFMMC0
;
ObFlFMMC0AR1_v)q.UjcG)Uhh
WRRCRoMHCsORR5
RSRRQQhaR_j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRQQhaR_4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRQQhaR_.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRQQhaR_d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRQQhaR_c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRQQhaR_6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRQQhaR_n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRQQhaR_(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRQQhaR_U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRQQhaR_g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRQQhaR_q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRQQhaR_A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRQQhaR_B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRQQhaR_7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRQQhaR_ :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRQQhaR_w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
RRRRRRRRRRQQhaj_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha4_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha._4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhad_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhac_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha6_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhan_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha(_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaU_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhag_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaq_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaA_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaB_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha7_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha _4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaw_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R

RRRRRRRRRhRQQ.a_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
RRRRRRRRRQRRh_Qad:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
"RSRRRR;2R
RSRb0Fs5SR
Sq)7a:qRR0FkR8#0_oDFHPO_CFO0s(5RRFR8IFM0RRj2;S
S)iBphRR:HRMR#_08DHFoO
R;SBS)pRi :MRHR0R#8F_DoRHO:'=R]
';S S)RRRR:MRHR0R#8F_DoRHO:'=R]
';SqS)7R7):MRHR0R#8F_Do_HOP0COFRs54RjR8MFI0jFR2
R;SBSWpRih:MRHR0R#8F_DoRHO;S
SWiBp RR:HRMR#_08DHFoO=R:R''];S
SWR RRRR:HRMR#_08DHFoO=R:R''];S
SW7q7)RR:HRMR#_08DHFoOC_POs0F5jR4RFR8IFM0RRj2;S
SWa7qqRR:HRMR#_08DHFoOC_POs0F5RR(RI8FMR0FjS2
RRRRR2RR;M
C8FROlMbFC;M0
F
OlMbFCRM01)A_qjvcgcnGRR
RoCCMsRHO5SR
RQRRh_QajRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_Qa4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_Qa.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_QadRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_QacRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_Qa6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_QanRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_Qa(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_QaURR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_QagRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_QaqRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_QaARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_QaBRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_Qa7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_Qa RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_QawRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
RRRRRRRRRQRRh_Qa4:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RRRRRRRRRRRQahQ_R.j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R..:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R. :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
RRRRRRRRRRQQhaj_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha4_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha._dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhad_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhac_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha6_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhan_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha(_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaU_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhag_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaq_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaA_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaB_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha7_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha _dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaw_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jjRR
SR2RRRS;
RFRbsR05
)SS7qqaRF:Rk#0R0D8_FOoH_OPC05FsRRdR8MFI0jFR2
R;SBS)pRiR:MRHR0R#8F_DoRHO;S
S)iBp RR:HRMR#_08DHFoO=R:R''];S
S)R RRRR:HRMR#_08DHFoO=R:R''];S
S)7q7)RR:HRMR#_08DHFoOC_POs0F54R4RFR8IFM0RRj2;S
SWiBpRRR:HRMR#_08DHFoO
R;SBSWpRi :MRHR0R#8F_DoRHO:'=R]
';S SWRRRR:MRHR0R#8F_DoRHO:'=R]
';SqSW7R7):MRHR0R#8F_Do_HOP0COFRs54R4R8MFI0jFR2
R;S7SWqRaq:MRHR0R#8F_Do_HOP0COFRs5d8RRF0IMF2Rj
RSRRRRRR
2;CRM8ObFlFMMC0
;
ObFlFMMC0AR1_v)qcnjgG)chR
H#RCRoMHCsORR5
RSRRQQhaR_j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRQQhaR_4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRQQhaR_.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRQQhaR_d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRQQhaR_c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRQQhaR_6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRQQhaR_n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRQQhaR_(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRQQhaR_U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRQQhaR_g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRQQhaR_q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRQQhaR_A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRQQhaR_B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRQQhaR_7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRQQhaR_ :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRQQhaR_w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
RRRRRRRRRRQQhaj_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha4_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha._4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhad_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhac_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha6_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhan_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha(_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaU_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhag_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaq_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaA_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaB_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha7_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha _4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaw_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R

RRRRRRRRRhRQQ.a_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
RRRRRRRRRQRRh_Qad:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qad:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
"RSRRRR;2R
RSRb0Fs5SR
Sq)7a:qRR0FkR8#0_oDFHPO_CFO0sd5RRFR8IFM0RRj2;S
S)iBphRR:HRMR#_08DHFoO
R;SBS)pRi :MRHR0R#8F_DoRHO:'=R]
';S S)RRRR:MRHR0R#8F_DoRHO:'=R]
';SqS)7R7):MRHR0R#8F_Do_HOP0COFRs54R4R8MFI0jFR2
R;SBSWpRiR:MRHR0R#8F_DoRHO;S
SWiBp RR:HRMR#_08DHFoO=R:R''];S
SWR RRRR:HRMR#_08DHFoO=R:R''];S
SW7q7)RR:HRMR#_08DHFoOC_POs0F54R4RFR8IFM0RRj2;S
SWa7qqRR:HRMR#_08DHFoOC_POs0F5RRdRI8FMR0FjS2
RRRRR2RR;M
C8FROlMbFC;M0
F
OlMbFCRM01)A_qjvcgcnGhHWR#R
RoCCMsRHO5SR
RQRRh_QajRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_Qa4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_Qa.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_QadRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_QacRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_Qa6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_QanRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_Qa(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_QaURR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_QagRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_QaqRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_QaARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_QaBRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_Qa7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_Qa RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQRRh_QawRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
RRRRRRRRRQRRh_Qa4:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RRRRRRRRRRRQahQ_R.j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R..:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R. :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R.w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
RRRRRRRRRRQQhaj_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha4_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha._dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhad_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhac_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha6_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhan_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha(_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaU_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhag_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaq_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaA_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaB_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha7_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha _dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaw_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jjRR
SR2RRRS;
RFRbsR05
)SS7qqaRF:Rk#0R0D8_FOoH_OPC05FsRRdR8MFI0jFR2
R;SBS)pRiR:MRHR0R#8F_DoRHO;S
S)iBp RR:HRMR#_08DHFoO=R:R''];S
S)R RRRR:HRMR#_08DHFoO=R:R''];S
S)7q7)RR:HRMR#_08DHFoOC_POs0F54R4RFR8IFM0RRj2;S
SWiBphRR:HRMR#_08DHFoO
R;SBSWpRi :MRHR0R#8F_DoRHO:'=R]
';S SWRRRR:MRHR0R#8F_DoRHO:'=R]
';SqSW7R7):MRHR0R#8F_Do_HOP0COFRs54R4R8MFI0jFR2
R;S7SWqRaq:MRHR0R#8F_Do_HOP0COFRs5d8RRF0IMF2Rj
RSRRRRRR
2;CRM8ObFlFMMC0
;

lOFbCFMM10RAq_)vgcjnhGc)RhWHR#
RMoCCOsHR
5RSRRRQahQ_:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RRRRRRRRRRRQahQ_R4j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R44:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R46:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R47:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4 :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
RRRRRRRRRRQQhaj_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha4_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha._.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhad_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhac_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha6_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhan_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha(_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaU_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhag_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaq_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaA_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaB_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha7_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha _.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaw_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R

RRRRRRRRRhRQQda_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"SR
RRRR2
R;SbRRF5s0RS
S)a7qqRR:FRk0#_08DHFoOC_POs0F5RRdRI8FMR0Fj;2R
)SSBhpiRH:RM#RR0D8_FOoHRS;
Sp)Bi: RRRHMR8#0_oDFH:OR=]R''S;
SR) R:RRRRHMR8#0_oDFH:OR=]R''S;
S7)q7:)RRRHMR8#0_oDFHPO_CFO0s45R48RRF0IMF2RjRS;
SpWBi:hRRRHMR8#0_oDFH;OR
WSSB piRH:RM#RR0D8_FOoHRR:=';]'
WSS RRRRH:RM#RR0D8_FOoHRR:=';]'
WSSq)77RH:RM#RR0D8_FOoH_OPC05FsRR44RI8FMR0Fj;2R
WSS7qqaRH:RM#RR0D8_FOoH_OPC05FsRRdR8MFI0jFR2R
SRRRRR;R2
8CMRlOFbCFMM
0;
lOFbCFMM10RAq_)vgU4.RG.HR#
RMoCCOsHR
5RSRRRQahQ_:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RRRRRRRRRRRQahQ_R4j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R44:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R46:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R47:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4 :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
RRRRRRRRRRQQhaj_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha4_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha._.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhad_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhac_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha6_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhan_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha(_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaU_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhag_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaq_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaA_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaB_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha7_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha _.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaw_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R

RRRRRRRRRhRQQda_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"SR
RRRR2
R;SbRRF5s0RR
RRRSRRRRRR7R)qRaq:kRF00R#8F_Do_HOP0COFRs548RRF0IMF2RjRS;
Sp)Bi:RRRRHMR8#0_oDFH;OR
)SSB piRH:RM#RR0D8_FOoHRR:=';]'
)SS RRRRH:RM#RR0D8_FOoHRR:=';]'
)SSq)77RH:RM#RR0D8_FOoH_OPC05FsRR4.RI8FMR0Fj;2R
WSSBRpiRH:RM#RR0D8_FOoHRS;
SpWBi: RRRHMR8#0_oDFH:OR=]R''S;
SRW R:RRRRHMR8#0_oDFH:OR=]R''S;
S7Wq7:)RRRHMR8#0_oDFHPO_CFO0s45R.8RRF0IMF2RjRS;
SqW7a:qRRRHMR8#0_oDFHPO_CFO0s45RRFR8IFM0R
j2SRRRRRRR2C;
MO8RFFlbM0CM;O

FFlbM0CMR_1A)Uqv4Gg..Rh)HR#
RMoCCOsHR
5RSRRRQahQ_:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RRRRRRRRRRRQahQ_R4j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R44:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R46:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R47:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4 :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
RRRRRRRRRRQQhaj_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha4_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha._.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhad_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhac_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha6_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhan_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha(_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaU_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhag_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaq_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaA_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaB_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha7_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha _.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaw_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R

RRRRRRRRRhRQQda_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"SR
RRRR2
R;SbRRF5s0RS
S)a7qqRR:FRk0#_08DHFoOC_POs0F5RR4RI8FMR0Fj;2R
)SSBhpiRH:RM#RR0D8_FOoHRS;
Sp)Bi: RRRHMR8#0_oDFH:OR=]R''S;
SR) R:RRRRHMR8#0_oDFH:OR=]R''S;
S7)q7:)RRRHMR8#0_oDFHPO_CFO0s45R.8RRF0IMF2RjRS;
SpWBi:RRRRHMR8#0_oDFH;OR
WSSB piRH:RM#RR0D8_FOoHRR:=';]'
WSS RRRRH:RM#RR0D8_FOoHRR:=';]'
WSSq)77RH:RM#RR0D8_FOoH_OPC05FsRR4.RI8FMR0Fj;2R
WSS7qqaRH:RM#RR0D8_FOoH_OPC05FsRR4R8MFI0jFR2R
SRRRRR;R2
8CMRlOFbCFMM
0;
lOFbCFMM10RAq_)vgU4.hG.WRR
RMoCCOsHR
5RSRRRQahQ_:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RRRRRRRRRRRQahQ_R4j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R44:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R46:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R47:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4 :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
RRRRRRRRRRQQhaj_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha4_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha._.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhad_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhac_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha6_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhan_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha(_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaU_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhag_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaq_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaA_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaB_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha7_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha _.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaw_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R

RRRRRRRRRhRQQda_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"SR
RRRR2
R;SbRRF5s0RS
S)a7qqRR:FRk0#_08DHFoOC_POs0F5RR4RI8FMR0Fj;2R
)SSBRpiRH:RM#RR0D8_FOoHRS;
Sp)Bi: RRRHMR8#0_oDFH:OR=]R''S;
SR) R:RRRRHMR8#0_oDFH:OR=]R''S;
S7)q7:)RRRHMR8#0_oDFHPO_CFO0s45R.8RRF0IMF2RjRS;
SpWBi:hRRRHMR8#0_oDFH;OR
WSSB piRH:RM#RR0D8_FOoHRR:=';]'
WSS RRRRH:RM#RR0D8_FOoHRR:=';]'
WSSq)77RH:RM#RR0D8_FOoH_OPC05FsRR4.RI8FMR0Fj;2R
WSS7qqaRH:RM#RR0D8_FOoH_OPC05FsRR4R8MFI0jFR2R
SRRRRR;R2
8CMRlOFbCFMM
0;
lOFbCFMM10RAq_)vgU4.hG.)RhWHR#
RMoCCOsHR
5RSRRRQahQ_:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRQahQ_:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RRRRRRRRRRRQahQ_R4j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R44:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R46:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R47:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4 :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_R4w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
RRRRRRRRRRQQhaj_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha4_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha._.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhad_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhac_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha6_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhan_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha(_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaU_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhag_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaq_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaA_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaB_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha7_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQha _.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaw_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R

RRRRRRRRRhRQQda_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"SR
RRRR2
R;SbRRF5s0RS
S)a7qqRR:FRk0#_08DHFoOC_POs0F5RR4RI8FMR0Fj;2R
)SSBhpiRH:RM#RR0D8_FOoHRS;
Sp)Bi: RRRHMR8#0_oDFH:OR=]R''S;
SR) R:RRRRHMR8#0_oDFH:OR=]R''S;
S7)q7:)RRRHMR8#0_oDFHPO_CFO0s45R.8RRF0IMF2RjRS;
SpWBi:hRRRHMR8#0_oDFH;OR
WSSB piRH:RM#RR0D8_FOoHRR:=';]'
WSS RRRRH:RM#RR0D8_FOoHRR:=';]'
WSSq)77RH:RM#RR0D8_FOoH_OPC05FsRR4.RI8FMR0Fj;2R
WSS7qqaRH:RM#RR0D8_FOoH_OPC05FsRR4R8MFI0jFR2R
SRRRRR;R2
8CMRlOFbCFMM
0;
lOFbCFMM10RAq_vBR4nHR#
SMoCCOsHR
5RShSR at_)tQt S)RSRS:LRH0S=S:';j'RS
SR)B_ StSSRS:LRH0S=S:';j'R-SS-jRB
RSSq _)tSSSSL:RHS0RS':=jR';SRRRR-S-RRB4
RSSA _)tSSSSL:RHS0RS':=jS';SR--BS.
S_R7)R tSSSS:HRL0SRS:j=''S;S-B-RdS
SRuam_UUG_pvza _)t:SSR0LHR:SS=''j;RRSR-RS-cRB
RSSA_maU_GUvazp_t) SRS:LRH0S=S:';j'SRRRSR--BS6
SQRuuQ ph4 _nnG4_pvza _)t:4SR0LHR:SS=''j;-SS-nRB
RSSu Qup Qh_G4n4vn_z_pa). tSL:RHS0RS':=jS';SR--B
(
SaSRmzumaauz_p1  RBaRRRRR:SSR0LH_OPC05Fs4FR8IFM0RRj2:"=RjRj";-S-RvBmAq,RBvBz_t) ,zRvpUa_GRU,vazp_G4n4/nR/g{B,}BUR=RRR,jjR,j4R,4jR
44SaSRm7uq7A1z_Wpm h)QuRzaR:SSR0LH_OPC05Fs4FR8IFM0RRj2:"=RjRj";-RS-qR7aRq,vazp_UUG,zRvp4a_nnG4,QR1tXh aRRS/B/{4B4,4Rj}=jRj,4Rj,jR4,4R4
RSSaqmu7z71Au_zuQ )hauzRSRS:HRL0SRSS=R:R''jRRR;SR--qzBBv _)t7,RqBaqRRSSS/R/R.B4Rj=R,
R4SaSRm7uq7A1z_)Bq) Y1pa BR:SSR0LH_OPC05Fs4FR8IFM0RRj2:"=RjRj";-RS-mRptjQB,tpmQ,B4qzBBv,BQt  h) qa7q_B)R)Y/B/{4Rc,B}4dRj=j,4Rj,jR4,4R4
S
SRaAmmuzaz1a_ Bp a:SSR0LH_OPC05Fs4FR8IFM0RRj2:"=RjRj";-RS-vBmAq,RBvBz_t) ,zRvpUa_GRU,vazp_G4n4RnR/{/RB,4nB}46Rj=j,4Rj,jR4,4R4
RSSAqma7z71Am_pWQ )hauzR:SSR0LH_OPC05Fs4FR8IFM0RRj2:"=RjRj";-RS-a7qqv,Rz_paU,GURpvzan_4G,4nRt1Qha XQ/hR/{RRB,4UB}4(Rj=j,4Rj,jR4,4R4
RSSAqma7z71Au_zuQ )hauzR:SSR0LHRSSSRR:='Rj'RR;RSq--BvBz_t) ,qR7aRq7RSRSSR//RgB4Rj=R,
R4SASRm7aq7A1z_)Bq) Y1pa BR:SSR0LH_OPC05Fs4FR8IFM0RRj2:"=RjRj";-RS-tpmQ,BjRtpmQ,B4RBqBzQvB,QRBRSRS/R/R{4B.,.RBjj}=j4,j,,4j4S4
SmRv7U _GSURSRS:LRH0SRSS:'=Rj;'RR-S-R.B.RS

S_Rq1hQt S7RSRS:LRH0SRSS:'=Rj;'RR-RS-.RBdS
SR1A_Q th7SRSSL:RHS0RS:SR=jR''RRRSR--B
.cS
2;SsbF0
S5
qSSSRS:HSMR#_08DHFoOC_POs0F5R468MFI0jFR2RR;RS
SA:SSRRHMR#RR0D8_FOoH_OPC05Fs486RF0IMF2RjRS;R
BSSSRS:HSMR#_08DHFoOC_POs0F5R468MFI0jFR2RR;
7SSSRS:HSMR#_08DHFoOC_POs0F5R468MFI0jFR2RR;
mSSSRS:FRk0S8#0_oDFHPO_CFO0s45dRI8FMR0Fj;2R
BSSpSiS:MRHR0S#8F_DoRHO;SR
SSB SH:RM#RS0D8_FOoHR
;RS)SQ1maau:RSRRHMS8#0_oDFH;ORRR
SRSRRQa)1ARmaSH:RM#RS0D8_FOoHR
;RS)Sm1maau:RSRRHMS8#0_oDFH;ORRS
Sma)1ARmaSH:RM#RS0D8_FOoHR
;RS]SqmRp7SRS:H#MS0D8_FOoHR
;RS]SAmSp7SH:RM#RS0D8_FOoHR
;RS]SBmSp7SH:RM#RS0D8_FOoHR
;RS]S7mSp7SH:RM#RS0D8_FOoHR
;RS]Smmap7m:uSRRHMS8#0_oDFH;ORRS
Smp]m7aAmSH:RM#RS0D8_FOoHR
;RSpSmmaq7m:uSRSHM#_08DHFoORR;
mSSp7mqASma:MRHR0S#8F_DoRHO;SR
S7q71azAm:uSRRHMS8#0_oDFH;ORRS
Sq177zmAAaRS:HSMR#_08DHFoO
R;SmSBSRS:FRk0S8#0_oDFH;OR
BSSQ:SSRRHMS8#0_oDFH;ORRSR
SBqBzQvBSRS:HSMR#_08DHFoORR;
qSSBvBzBRmRRRRRR:RSR0FkR0S#8F_DoRHO;S
S1hQt QXahRS:H#MS0D8_FOoHR
;RSQS1tXh aamzRRRRRRR:FRk0S8#0_oDFHRORSSSS
;S2RC

MO8RFFlbM0CM;O

FFlbM0CMR_1AQ7m_pHYR#SR
oCCMsSHO5S

Sth _Qa)t)t R:SSR0LHSSSS:j=''S;
ShuQ_uaY :SSR0LH_OPC0RFs586RF0IMF2RjS":=jjjjj;j"
uSSzzppuSSS:HRL0SSSS':=j
';SmSQ_q1ah)7q7:SSRs#0HSMoS=S:"_1ApveBm;1"
QSShp7 qeY_qSpS:HRL0C_POs0FRR568MFI0jFR2:RS=j"jjjjj"S;
Samz7q pYq_epSRS:HRL0C_POs0FRR568MFI0jFR2:RS=j"jjjjj"2
S;SS
b0FsR
S5SqSuBtiq Q_uhSRS:MRHFRk0#_08koDFHRO;
pSSq]aB_uQhzea_q pzRRS:HSMR#_08DHFoO
;RSpSBm_Bi AhqpS S:MRHR0S#8F_Do;HORS
SQzhuap_Bi:SSRRHMS8#0_oDFHRO;
mSSzzauap_Bi:SSRRHMS8#0_oDFHRO;
mSSzzauah_ q ApSRS:HSMR#_08DHFoO=R:';]'RS
S7z_maS_4SRS:HSMR#_08DHFoOR;RRS
S7z_maS_jSRS:HSMR#_08DHFoOR;R
7SS__Qh4SSS:kRF0#RS0D8_FOoH;SR
SQ7_hS_jSRS:FRk0S8#0_oDFHRO;
1SSBSpiSRS:HSMR#_08DHFoOS;R
1SS7SQSSH:RM#RS0D8_FOoH;
RSS_SB) _1pSSS:MRHR0S#8F_Do;HORSR
Sm17S:SSR0FkR0S#8F_DoRHO
2SR;


CRM8ObFlFMMC0
;RRF
OlMbFCRM01vA_Q_uQacX_p qhRSR
oCCMsSHO5SRS
7SSQRe)S:SSR0LH_OPC05FsR8cRF0IMF2RjR:RS=4R"4444"RR;RRRRR-S-RV)CR	BDRP8HHs8C
7SSQRewS:SSR0LH_OPC05FsR8(RF0IMF2RjR:RS=4R"4j44j"jj;SRS-w-RCLC8NRO	8HHP8
CsSQS7eSTRSRS:L_H0P0COFRs54FR8IFM0RRj2R=S:Rj"j"R;RRRRRR-SS-BRemHR8PCH8sS
Saa 1_7vm SRS:HRL0SRSS=S:R''j;S
Saa 1_aAQ1SRS:HRL0C_POs0F5RRd8MFI0jFR2:RS=4R"j"j4
;S2Rb
SFRs0S
5RS-SS-lBFlRFMQCM0sOVNCHRuMS#
SSuzSRS:HSMR#_08DHFoORR;
pSSAS hSRS:HSMR#_08DHFoORR;
SRS)amzBSqpSRS:HSMR#_08DHFoOC_POs0F584RF0IMF2RjR
;RR SSh u71S )SH:RM0S#8F_DoRHO;
RSSRRRRRRRSBu7iStSSH:RM0S#8F_DoRHO;SR
S-S-Ra7qqQjRMs0CVCNORMbH#S
S7SujSRS:HkMF00S#8D_kFOoHRS;R
7SShSjSSH:RM0FkR8#0_FkDoRHO;RR
SjS7mmuv7S S:MRHS8#0_oDFH;ORRRR
SjS77paXuSuS:MRHS8#0_oDFH;ORRS
RS77jauXph:SSRRHMS8#0_oDFH;ORRS
RSa7jX puh:SSRSHM#_08DHFoORR;RRS
SjS77p)XuSuS:kRF00S#8F_DoRHO;SR
R7RSjX7)pSuhSF:RkS0R#_08DHFoORR;
SRS7Xj)phu SRS:HSMR#_08DHFoORR;
SRS7Bj77SuSSF:RkS0R#_08DHFoORR;
7SSj77BhSSS:kRF0#RS0D8_FOoHR
;RR7SSj B7hSSS:MRHS8#0_oDFH;ORR
SSRSRS7Xja]71uSRS:H#MS0D8_FOoHR
;RR7SSj]aX1S hSH:RM#RS0D8_FOoHR
;RRSRRS]7j17aXqSaqSH:RM#RS0D8_FOoH_OPC05FsR8(RF0IMF2RjR
;RRSRS71j]1  )h:SSRSHM#_08DHFoORR;SRR
SjS7)1X] ShS:MRHS8#0_oDFH;ORRR
RSjS7] 171  )h:SSRRHMS8#0_oDFH;ORRRS
S7RSj)]1Xa7qq:SSR0FkR0S#8F_Do_HOP0COFRs5(FR8IFM0RRj2;RR
SjS7]Y1Aap BiS7S:kRF0#RS0D8_FOoHR
;RR7SSjh1YBSSS:kRF0#RS0D8_FOoHR
;RR7SSj) )1BYhSRS:FRk0S8#0_oDFH;ORRR
SRRRRRjS7]Y1Aap Bim1h1BYhSF:RkS0R#_08DHFoORR;
SSS-7-Rq4aqR0QMCNsVObCRH
M#SuS74SSS:MRHFRk0#_08koDFH;ORRS
S7Sh4SRS:HkMF00R#8D_kFOoHRR;R
SRS7a47XupuSRS:HSMR#_08DHFoORR;
SRS7a47XhpuSRS:H#MS0D8_FOoHR
;RRSRS7X4aphu SRS:HSMR#_08DHFoORR;
SRS7)47XupuSRS:FRk0S8#0_oDFH;OR
RSRS774)uXph:SSR0FkR0S#8F_DoRHO;RR
S4S7)uXp ShS:MRHS8#0_oDFH;OR
SRS7B477SuSSF:RkS0R#_08DHFoORR;
7SS477BhSSS:kRF0SRR#_08DHFoORR;
SRS774B ShSSH:RM0S#8F_DoRHO;RR
R7SS4]aX1Su7SH:RM#RS0D8_FOoHR
;RR7SS4]aX1S hSH:RM0S#8F_DoRHO;
RRS4S7]X1a7qqaSRS:HSMR#_08DHFoOC_POs0F5RR(8MFI0jFR2RR;
SRRS]741)1  ShS:MRHS8#0_oDFH;ORRS
RS)74X ]1h:SSRRHMS8#0_oDFH;OR
SRRS]74117  h) SRS:HSMR#_08DHFoORR;
SSR714])qX7aSqS:kRF0RRR#_08DHFoOC_POs0F5RR(8MFI0jFR2RR;
SRS7Y41hSBSSF:RkS0R#_08DHFoORR;
SRS7)4 )h1YB:SSR0FkR0S#8F_DoRHO;RR
S4S7hYm1hSBS:kRF0#RS0D8_FOoHR
;RS-SS-qR7aRq.QCM0sOVNCHRbMS#
S.7uS:SSRFHMk#0R0k8_DHFoO
R;ShS7.SSS:MRHFRk0#_08koDFH;ORRS
RS77.auXpu:SSRSHM#_08DHFoORR;
SRS7a.7XhpuSRS:HSMR#_08DHFoORR;
SRRSa7.X puh:SSRRHMS8#0_oDFH;ORRS
RS77.)uXpu:SSR0FkR0S#8F_DoRHO;SR
R7RS.X7)pSuhSF:RkS0R#_08DHFoORR;
SRS7X.)phu SRS:HSMR#_08DHFoORR;
SRS7B.77SuSSF:RkS0R#_08DHFoORR;
7SS.77BhSSS:kRF0#RS0D8_FOoHR
;RR7SS. B7hSSS:MRHS8#0_oDFH;OR
SRRSa7.Xu]17:SSRSHM#_08DHFoORR;
SRS7X.a]h1 SRS:H#MS0D8_FOoHRS;RSRR
RSRRR.S7]X1a7qqaSRS:H#MS0D8_FOoH_OPC05FsR8(RF0IMF2RjR
;RRSRS71.]1  )h:SSRSHM#_08DHFoORR;
SRS7X.)]h1 SRS:H#MS0D8_FOoHR
;RRSRS71.]7  1)S hSH:RM0S#8F_DoRHO;RR
S7RS.)]1Xa7qq:SSR0FkR0S#8F_Do_HOP0COFRs5(FR8IFM0RRj2;RR
S.S71BYhS:SSR0FkR0S#8F_DoRHO;RR
S.S7 1))YShBSF:RkS0R#_08DHFoO
R;R7SS.1hmYShBSF:RkS0R#_08DHFoORR;
SSS-7-RqdaqR0QMCNsVObCRH
M#SuS7dSSS:MRHFRk0#_08koDFH;ORRS
S7ShdSRS:HkMF00R#8D_kFOoHRR;
SdS77paXuSuS:MRHR0S#8F_DoRHO;RR
SdS77paXuShS:MRHS8#0_oDFH;ORRR
RSdS7auXp ShS:MRHR0S#8F_DoRHO;RR
SdS77p)XuSuS:kRF0#RS0D8_FOoHR
;RSSRR7)d7XhpuSRS:FRk0S8#0_oDFH;OR
SRS7Xd)phu SRS:H#MS0D8_FOoHR
;RR7SSd77BuSSS:kRF0#RS0D8_FOoHR
;RSdS77hB7S:SSR0FkR0S#8F_DoRHO;RR
SdS7Bh7 S:SSRSHM#_08DHFoORR;
SRRSa7dXu]17:SSRSHM#_08DHFoORR;
SRS7Xda]h1 SRS:H#MS0D8_FOoHRR;R
SRRRdS7]X1a7qqaSRS:HSMR#_08DHFoOC_POs0F5RR(8MFI0jFR2RR;
SRRS]7d1)1  ShS:MRHS8#0_oDFH;ORRS
RS)7dX ]1h:SSRSHM#_08DHFoORR;
SRRS]7d117  h) SRS:H#MS0D8_FOoHR
;RRSSR71d])qX7aSqS:kRF0#RS0D8_FOoH_OPC05FsR8(RF0IMF2RjR
;RR7SSdh1YBSSS:kRF0#RS0D8_FOoHR
;SR7SSd) )1BYhSRS:FSk0#_08DHFoORR;
SRS7mdh1BYhSRS:FRk0S8#0_oDFH;ORRS
SSR--BBpmiMRQ0VCsNROCb#HM
BSSiSuSSH:RM0FkR8#0_FkDoRHO;
RRSiSBhSSS:MRHFRk0#_08koDFH;ORRS
RSiBp7paXuSuS:MRHR0S#8F_DoRHO;RR
SpSBiX7apSuhSH:RM0S#8F_DoRHO;RR
RBSSpXiaphu SRS:HSMR#_08DHFoORR;
RSRSiBp7p)XuSuS:kRF0#RS0D8_FOoHR
;RSSRRB7pi)uXph:SSR0FkR0S#8F_DoRHO;RR
RBSSpXi)phu SRS:H#MS0D8_FOoHR
;RRSRSBapiXu]17:SSRSHM#_08DHFoORR;
SRSBapiX ]1h:SSRSHM#_08DHFoORR;
RSRRRRRRpSBi]aX1atq :SSRSHM#_08DHFoORR;
SRRSiBp)1X] ShS:MRHS8#0_oDFH;ORRR
SRRRRSiBp]Y1AaS S:kRF0#RS0D8_FOoHR
;RS-SS-MRzHsPC#RNDvQQuRpupR0QMCNsVObCRH
M#RuSSpzpuS:SSRRHMS8#0_oDFH;ORRS
RSpup)S wSRS:H#MS0D8_FOoHR
;RRuSSpmppBSiSSF:RkS0R#_08DHFoORR;
SSS-z-RMCHPsD#NRuvQQpRupCR1sDHNRMBFVkHosHN0F)MRC#oH0RCsQCM0sOVNCHRbMR#
SpSuptBw1Q)7SRS:H#MS0D8_FOoHR
;RRuSSpwpBt)1) a1 SRS:H#MS0D8_FOoHR
;RRuSSpwpBtB1)pSiS:MRHS8#0_oDFH;ORRS
RSpupB1wt)S7mSF:RkS0R#_08DHFoOSR
2
;
CRM8ObFlFMMC0
;R
vBmu mhh1aRA._QBR
RRht  B)QRR5
RRRRRR--BMENM#CDR8NMRNTk8q#R0
0sRRRRQ_.B1epq h_QQqa_7R7):0R1soHMRR:=RL"j44444jjjj;4"
RRRR1Az_7q7)R(cRRR:1H0sM:oR=jR"L4j4j2"R;m
u)5aR
SRS1pABiSQSSH:RM#RS0D8_FOoHR
;RR1SSAQ)WS:SSRRHMS8#0_oDFH;ORRS
RS11AaSAQSRS:HSMR#_08DHFoORR;
SRS17Aq)SQ(SRS:HSMR#_08DHFoORR;
SRS17Aq)SQnSRS:HSMR#_08DHFoORR;
SRS17Aq)SQ6SRS:HSMR#_08DHFoORR;
SRS17Aq)SQcSRS:HSMR#_08DHFoORR;
SRS17Aq)SQdSRS:HSMR#_08DHFoORR;
SRS17Aq)SQ.SRS:HSMR#_08DHFoORR;
SRS17Aq)SQ4SRS:HSMR#_08DHFoORR;
SRS17Aq)SQjSRS:HSMR#_08DHFoORR;
SRS1qA7aSQ(SRS:HSMR#_08DHFoORR;
SRS1qA7aSQnSRS:HSMR#_08DHFoORR;
SRS1qA7aSQ6SRS:HSMR#_08DHFoORR;
SRS1qA7aSQcSRS:HSMR#_08DHFoORR;
SRS1qA7aSQdSRS:HSMR#_08DHFoORR;
SRS1qA7aSQ.SRS:HSMR#_08DHFoORR;
SRS1qA7aSQ4SRS:HSMR#_08DHFoORR;
SRS1qA7aSQjSRS:HSMR#_08DHFoORR;
SRS1QBpS:SSRRHMS8#0_oDFH;ORRS
RSq17QSSS:MRHR0S#8F_DoRHO;
R
R1SSAa7qmS(SSF:RkS0R#_08DHFoORR;
SRS1qA7aSmnSRS:FRk0S8#0_oDFH;ORRS
RS71Aq6amS:SSR0FkR0S#8F_DoRHO;RR
SAS17mqacSSS:kRF0#RS0D8_FOoHR
;RR1SSAa7qmSdSSF:RkS0R#_08DHFoORR;
SRS1qA7aSm.SRS:FRk0S8#0_oDFH;ORRS
RS71Aq4amS:SSR0FkR0S#8F_DoRHO;RR
SAS17mqajSSS:kRF0#RS0D8_FOoHR
;RR1SSAiqBmSSS:kRF0#RS0D8_FOoHR
;RRQSS.)BQTSSS:kRF0#RS0D8_FOoHRR;
S.SQBzWiuSSS:kRF0#RS0D8_FOoH;S
RSp1BmSSS:kRF0#RS0D8_FOoHR
;RR1SSB pmS:SSR0FkR0S#8F_DoRHO;RR
S7S1qSmSSF:RkS0R#_08DHFoORR;
SRS1m7q SSS:kRF0#RS0D8_FOoHR
R
RRRRRRRR2 ;
hB7Rmmvuha h;B

mmvuha hR_1A1
uQRtRR )h Q5BR
RRRR-RR-ERBNCMMDN#RMT8Rk#N8R0q0sR
RRzRA17_q7c)(R:RRRs10HRMo:"=Rj4LjjR4"2u;
mR)a5R
RRRRRRRRRRRRRRAR1BQpiRRRRRRRRRRRRRRRRRRR:HRMRR0R#8F_DoRHO;R
RRRRRRRRRRRRRRAR1)RWQRRRRRRRRRRRRRRRRRRR:HRMRR0R#8F_DoRHO;R
RRRRRRRRRRRRRRAR11QaARRRRRRRRRRRRRRRRRRR:HRMRR0R#8F_DoRHO;R
RRRRRRRRRRRRRRAR1qQ7)(RRRRRRRRRRRRRRRRRR:HRMRR0R#8F_DoRHO;R
RRRRRRRRRRRRRRAR1qQ7)nRRRRRRRRRRRRRRRRRR:HRMRR0R#8F_DoRHO;R
RRRRRRRRRRRRRRAR1qQ7)6RRRRRRRRRRRRRRRRRR:HRMRR0R#8F_DoRHO;R
RRRRRRRRRRRRRRAR1qQ7)cRRRRRRRRRRRRRRRRRR:HRMRR0R#8F_DoRHO;R
RRRRRRRRRRRRRRAR1qQ7)dRRRRRRRRRRRRRRRRRR:HRMRR0R#8F_DoRHO;R
RRRRRRRRRRRRRRAR1qQ7).RRRRRRRRRRRRRRRRRR:HRMRR0R#8F_DoRHO;R
RRRRRRRRRRRRRRAR1qQ7)4RRRRRRRRRRRRRRRRRR:HRMRR0R#8F_DoRHO;R
RRRRRRRRRRRRRRAR1qQ7)jRRRRRRRRRRRRRRRRRR:HRMRR0R#8F_DoRHO;R
RRRRRRRRRRRRRRAR17Qqa(RRRRRRRRRRRRRRRRRR:HRMRR0R#8F_DoRHO;R
RRRRRRRRRRRRRRAR17QqanRRRRRRRRRRRRRRRRRR:HRMRR0R#8F_DoRHO;R
RRRRRRRRRRRRRRAR17Qqa6RRRRRRRRRRRRRRRRRR:HRMRR0R#8F_DoRHO;R
RRRRRRRRRRRRRRAR17QqacRRRRRRRRRRRRRRRRRR:HRMRR0R#8F_DoRHO;R
RRRRRRRRRRRRRRAR17QqadRRRRRRRRRRRRRRRRRR:HRMRR0R#8F_DoRHO;R
RRRRRRRRRRRRRRAR17Qqa.RRRRRRRRRRRRRRRRRR:HRMRR0R#8F_DoRHO;R
RRRRRRRRRRRRRRAR17Qqa4RRRRRRRRRRRRRRRRRR:HRMRR0R#8F_DoRHO;R
RRRRRRRRRRRRRRAR17QqajRRRRRRRRRRRRRRRRRR:HRMRR0R#8F_DoRHO;R
RRRRRRRRRRRRRRQRvRRRRRRRRRRRRRRRRRRRRRRR:HRMRR0R#8F_DoRHO;R
RRRRRRRRRRRRRRQR1RRRRRRRRRRRRRRRRRRRRRRR:HRMRR0R#8F_DoRHO;R
RRRRRRRRRRRRRRBR1iRQRRRRRRRRRRRRRRRRRRRR:HRMRR0R#8F_DoRHO;R
RRRRRRRRRRRRRRBR11RhQRRRRRRRRRRRRRRRRRRR:HRMRR0R#8F_DoRHO;R

RRRRRRRRRRRRR1RRAa7qmR(RRRRRRRRRRRRRR:RRR0FkR#RR0D8_FOoHRR;
RRRRRRRRRRRRR1RRAa7qmRnRRRRRRRRRRRRRR:RRR0FkR#RR0D8_FOoHRR;
RRRRRRRRRRRRR1RRAa7qmR6RRRRRRRRRRRRRR:RRR0FkR#RR0D8_FOoHRR;
RRRRRRRRRRRRR1RRAa7qmRcRRRRRRRRRRRRRR:RRR0FkR#RR0D8_FOoHRR;
RRRRRRRRRRRRR1RRAa7qmRdRRRRRRRRRRRRRR:RRR0FkR#RR0D8_FOoHRR;
RRRRRRRRRRRRR1RRAa7qmR.RRRRRRRRRRRRRR:RRR0FkR#RR0D8_FOoHRR;
RRRRRRRRRRRRR1RRAa7qmR4RRRRRRRRRRRRRR:RRR0FkR#RR0D8_FOoHRR;
RRRRRRRRRRRRR1RRAa7qmRjRRRRRRRRRRRRRR:RRR0FkR#RR0D8_FOoHRR;
RRRRRRRRRRRRR1RRAiqBmRRRRRRRRRRRRRRRR:RRR0FkR#RR0D8_FOoHRR;
RRRRRRRRRRRRR1RRu)QQTRRRRRRRRRRRRRRRR:RRR0FkR#RR0D8_FOoHRS;
S1SSuiQWzSuSSF:RkR0R#_08DHFoOR;
RRRRRRRRRRRRR1RRmRRRRRRRRRRRRRRRRRRRR:RRR0FkR#RR0D8_FOoHRR;
RRRRRRRRRRRRR1RRmR RRRRRRRRRRRRRRRRRR:RRR0FkR#RR0D8_FOoHRR;
RRRRRRRRRRRRRvRRmRRRRRRRRRRRRRRRRRRRR:RRR0FkR#RR0D8_FOoHRR;
RRRRRRRRRRRRRvRRmR RRRRRRRRRRRRRRRRRR:RRR0FkR#RR0D8_FOoHRR;
RRRRRRRRRRRRR1RRBRimRRRRRRRRRRRRRRRRR:RRR0FkR#RR0D8_FOoHRR;
RRRRRRRRRRRRR1RRB imRRRRRRRRRRRRRRRRR:RRR0FkR#RR0D8_FOoHRR;
RRRRRRRRRRRRRvRRBm1hdRRRRRRRRRRRRRRRR:RRR0FkR#RR0D8_FOoHRR;
RRRRRRRRRRRRRvRRBm1h.RRRRRRRRRRRRRRRR:RRR0FkR#RR0D8_FOoHRR;
RRRRRRRRRRRRRvRRBm1h4RRRRRRRRRRRRRRRR:RRR0FkR#RR0D8_FOoHRR;
RRRRRRRRRRRRRvRRBm1hjRRRRRRRRRRRRRRRR:RRR0FkR#RR0D8_FOoHRR;
RRRRRRRRRRRRRvRRBm1h RdRRRRRRRRRRRRRR:RRR0FkR#RR0D8_FOoHRR;
RRRRRRRRRRRRRvRRBm1h R.RRRRRRRRRRRRRR:RRR0FkR#RR0D8_FOoHRR;
RRRRRRRRRRRRRvRRBm1h R4RRRRRRRRRRRRRR:RRR0FkR#RR0D8_FOoHRR;
RRRRRRRRRRRRRvRRBm1h RjRRRRRRRRRRRRRR:RRR0FkR#RR0D8_FOoHRR
RR;R2
7 hRvBmu mhh
a;
vBmu mhh1aRA1_]m
1BRRRRRRRRRFRbs
05RRRRRRRRRRRRRRRRBvpiRF:Rk#0R0D8_FOoHR
R;RRRRRRRRRRRRRRRR BhqpRiv:MRHR0R#8F_DoRHO
RRRRRRRRRRRRRRR2 ;
hB7Rmmvuha h;B

mmvuha hR_1Ap11mBR
RRRRRRRRRb0Fs5R
RRRRRRRRRRRRRRpRBi:iRR0FkR8#0_oDFHROR;R
RRRRRRRRRRRRRRhR qiBpiRR:HRMR#_08DHFoOR
RRRRRRRRRRRRRR
2; Rh7Bumvmhh a
;

vBmu mhhRaR1]A_wBm1R
RRSMoCCOsH5SR
B]piwQ_7e#:R0MsHo":=jjLj";R2RS
SSsbF0S5
SSSSB]piwRR:FRk0#_08DHFoOS;
SSSSB]piwR hRM:HR8#0_oDFH
O;SSSSSiBp]zwuRH:RM0R#8F_Do
HORRRR2C;
MB8Rmmvuha hR
;

vBmu mhhRaR1pA_wBm1R
RRSbSSF5s0
SSSBppiwRR:FRk0#_08DHFoOS;
SpSBi pwh:RRH#MR0D8_FOoH;S
SSiBppzwuRH:RM0R#8F_Do
HOSSSS2C;
MB8Rmmvuha h;


Bumvmhh a1RRAt_)A)_7e
RRSMoCCOsH5)
St_AjB)z) :haRs#0H:Mo=L"jjjjjj;j"R)
St_A4B)z) :haRs#0H:Mo=L"jjjjjj;j"
tS)AB._z ))hRa:#H0sM=o:"jjLjjjjj;"2R
RRSbSSF5s0
SSSSA)tjF:Rk#0R0D8_FOoH;
RRSSSS)4tA:kRF00R#8F_Do;HO
SSSSA)t.F:Rk#0R0D8_FOoH;S
SStS)A7p  RhR:RHM#_08DHFoOS;
S)SStuAjWRvR:RHM#_08DHFoOS;
S)SStuA4WHv:M0R#8F_Do;HO
SSSSA)t.vuWRM:HR8#0_oDFH
O;SSSS)utAzRR:H#MR0D8_FOoH
SSSS
2;CRM8Bumvmhh a
R;
m
Bvhum Rha1QA_))_7eRRR
CSoMHCsOS5
QB)_z ))hRa:#H0sM=o:"jjLjjjjjjjjj2"R;SR
SFSbs
05SSSSQ )p7RR:FRk0#_08DHFoOS;
SQSS)7p  RhR:RHM#_08DHFoOS;
SQSS)RuzRM:HR8#0_oDFHSO;SSSSSSR
SQSS)vuWRH:RM0R#8F_Do
HORRRR2C;
MB8Rmmvuha hR
;
Bumvmhh aAR1_7p 7u_QR
RRSbSSF5s0
SSSumWvzRaj:kRF00R#8F_Do;HOSS
SSvuWm4zaRF:Rk#0R0D8_FOoH;S
SSvuWm.zaRF:Rk#0R0D8_FOoH;S
SS7p 7Rmh:kRF00R#8F_Do;HORS
SS7p 7:B1H#MR0D8_FOoH;S
SS7p 7iBp:RHM#_08DHFoOS;
S Sp7q77aH(:M0R#8F_Do;HO
SSSp7 77nqa:RHM#_08DHFoOS;
S Sp7q77aH6:M0R#8F_Do;HO
SSSp7 77cqa:RHM#_08DHFoOS;
S Sp7q77aHd:M0R#8F_Do;HO
SSSp7 77.qa:RHM#_08DHFoOS;
S Sp7q77aH4:M0R#8F_Do;HO
SSSp7 77jqa:RHM#_08DHFoOS;
S Sp777q7:)dH#MR0D8_FOoH;S
SS7p 77q7)H.:M0R#8F_Do;HO
SSSp7 7q)774M:HR8#0_oDFH
O;SpSS q777j7):RHM#_08DHFoOS;
S Sp7 77hM:HR8#0_oDFH
O;SpSS  77XH :M0R#8F_Do;HO
SSSp7 7):1aH#MR0D8_FOoH
SSSS
2;CRM8Bumvmhh a
R;
lOFbCFMM10RAm_Q_
m7RRRRRRRRRCRoMHCsORR5u_Qha YuRRRR:HRL0C_POs0F5RR6RI8FMR0Fj
2;RRRRRRRRRRRRRRRRRRRR-z-upupzR:RRR0LH;RR
RRRRRRRRRRRRRRRRRhRR at_)tQt :)RR0LHRR
RRRRRRRRRRRRRRRRRR-R-Q1m_a7qhqR)7:0R#soHMRR
RRRRRRRRRRRRRRRRR2
R;RRRRRRRRRFRbsR05
RRRRRRRRRRRRRRR7amz4SRSRRRR:MRHR8#0_oDFH
O;SSSS7amzjSRSRRRR:MRHR8#0_oDFH
O;SSSSBBpmiq hASp SH:RM0R#8F_Do;HO
SSSSapqBh]Quezaq pzSH:RM0R#8F_Do;HO
SSSSuQhzpaBiSSS:MRHR8#0_oDFH
O;SSSS74QhSSSS:kRF00R#8F_Do;HO
SSSSh7QjSSSSF:Rk#0R0D8_FOoH;S
SSzSmaauz AhqpS S:MRHR8#0_oDFH:OS=''];S
SSzSmaauzBSpiSRS:H#MR0D8_FOoH;S
SSqSuBtiq huQS:SSRFHMk#0S0D8_FOoHRRRRRRRRRRRRRRRRRR
RRRRRRRRRRRRRR
2;CRM8ObFlFMMC0
;

vBmu mhh1aRA _p7)_7ez_B)SR
SFSus50RRS
SShS RH:RM1RRap7_mBtQ;S
SS Sp7Ruz:kRF01RRap7_mBtQ2C;
MB8Rmmvuha h;


Bumvmhh a1RRAt_)A7q_)ReR
CRoMHCsORR5
SSSB)z) _hav m7R0:#soHMRR:="jjL"S;
StS)ABj_z ))h:aR#H0sM:oR=jR"Ljjjj"jj;S
SRRRR)4tA_)Bz)a hR0:#soHMRR:="jjLjjjjj
";SRSRRtR)AB._z ))h:aR#H0sM:oR=jR"Ljjjj"jj

2;b0FsRR5
RRRRR)RRtuAjW:vRRRHM#_08DHFoOS;
StR)AW4uvRR:H#MR0D8_FOoH;S
SRA)t.vuWRH:RM0R#8F_Do;HO
RSSB)z) :hRRRHM#_08DHFoOS;
StR)A7p  :hRRRHM#_08DHFoOR;
RRRRR)RRtRAj:kRF00R#8F_Do;HO
RSS)4tARF:Rk#0R0D8_FOoH;S
SRA)t.RR:FRk0#_08DHFoO2
S;
SRCRM8Bumvmhh a
;
-------------------------------------------------------------------------
---R-RRNADOF	AGRR:1QA_)jcj_e7)
---------------------------------------------------------------------------
vBmu mhhRaR1QA_)jcj_e7)RRR
oCCMsRHO5SR
RBRRz ))hva_mR7 :s#0HRMo:"=Rj"Lj;R
SR)RQc_jjB)z) Rha:s#0HRMo:"=RjjLjjjjjj
j"2b;
FRs05R
RRRRRRzRB)h) RH:RM0R#8F_Do;HO
RSSQ )p7R h:MRHR8#0_oDFH
O;SQSR)vuWRH:RM0R#8F_Do;HO
RRRRRRRRpQ) :7RR0FkR8#0_oDFHSO
2R;S
8CMRvBmu mhh
a;
-
---------------------------------------------------------------------------
-RARRD	NOARFG:AR1_)AqB m7_e7)
---------------------------------------------------------------------------
vBmu mhhRaR1AA_qm)B77 _)ReR
CRoMHCsORR5
BSSz ))hva_mR7 :s#0HRMo:"=Rj"Lj;S
SABq)m_7 B)z) Rha:s#0HRMo:"=RjjLjj
j"2b;
FRs05R
RRRRRRqRA)7Bm : hRRHM#_08DHFoOS;
S)Bz): hRRHM#_08DHFoOS;
S)AqB m7uRWv:MRHR8#0_oDFH
O;RRRRRRRRABq)mR7 :kRF00R#8F_Do
HOSS2;RM
C8mRBvhum ;ha
-
--------------------------------------------------------------
---A-RpiqBRXAmRQ:R)RQu5a)GG
2R-----------------------------------------------------------------
-RBumvmhh a1RRA)_Q_RQuRF
bs50R
RRRRRRRR7Rq):QdRRHM#_08DHFoOS;
S7Rq):Q.RRHM#_08DHFoOS;
S7Rq):Q4RRHM#_08DHFoOS;
S7Rq)RQj:MRHR8#0_oDFH
O;SBSRp:iQRRHM#_08DHFoOS;
S1RBQH:RM0R#8F_Do;HO
RSS7Q h:MRHR8#0_oDFH
O;SWSR :QRRRHM#_08DHFoOS;
SXR  H:RM0R#8F_Do;HO
RSSp) qhRR:H#MR0D8_FOoH;S
SRa)1:MRHR8#0_oDFH
O;SQSR)RQh:MRHR8#0_oDFH
O;SWSR7qqa(H:RM0R#8F_Do;HO
RSSWa7qqRn:H#MR0D8_FOoH;S
SRqW7a:q6RRHM#_08DHFoOS;
S7RWqcaq:MRHR8#0_oDFH
O;SWSR7qqadH:RM0R#8F_Do;HO
RSSWa7qqR.:H#MR0D8_FOoH;S
SRqW7a:q4RRHM#_08DHFoO
;SSWSR7qqajRR:H#MR0D8_FOoH;R
RRRRRRARRz:1YFRk0#_08DHFoOS;
S)R77FY:k#0R0D8_FOoH;S
SR) )RF:Rk#0R0D8_FOoH;S
SRmQ)z:aRR0FkR8#0_oDFH
O;S)SR7qqa(F:Rk#0R0D8_FOoH;SS
S7R)qnaq:kRF00R#8F_Do;HO
RSS)a7qqR6:FRk0#_08DHFoOS;
S7R)qcaq:kRF00R#8F_Do;HO
RSS)a7qqRd:FRk0#_08DHFoOS;
S7R)q.aq:kRF00R#8F_Do;HO
RSS)a7qqR4:FRk0#_08DHFoOS;
S7R)qjaqRF:Rk#0R0D8_FOoH
;S2SCR
MB8Rmmvuha h;-

--------------------------------------------------R
-pRAqABim:XRS_1AQ_.BwmQwR-R
-------------------------------------------------
-RBumvmhh a1RRA._QBQ_wwRmR
CRoMHCsORR5
RSRRBQ._q1peq _7R7):s#0HRMo:"=Rj4L44j44j4jj";
2
sbF0
R5RRRRRRRRRiBpQH:RM0R#8F_Do;HO
RSSB:1QRRHM#_08DHFoOS;
SaR1ARQ:H#MR0D8_FOoH;S
SRQW :MRHR8#0_oDFH
O;SqSR7d)Q:MRHR8#0_oDFH
O;SqSR7.)Q:MRHR8#0_oDFH
O;SqSR74)Q:MRHR8#0_oDFH
O;SqSR7j)QRH:RM0R#8F_Do;HO
RSS7QqagH:RM0R#8F_Do;HO
RSS7QqaUH:RM0R#8F_Do;HO
RSS7Qqa(H:RM0R#8F_Do;HO
RSS7QqanH:RM0R#8F_Do;HO
RSS7Qqa6H:RM0R#8F_Do;HO
RSS7QqacH:RM0R#8F_Do;HO
RSS7QqadH:RM0R#8F_Do;HO
RSS7Qqa.H:RM0R#8F_Do;HO
RSS7Qqa4H:RM0R#8F_Do;HO
RSS7QqajRR:H#MR0D8_FOoH;S
SRwwQma)1RH:RM0R#8F_Do;HO
RSS1QBpRH:RM0R#8F_Do;HO
RSS1Q7qRH:RM0R#8F_Do;HO
RRRRRRRRBRqiRm:FRk0#_08DHFoOS;
S.RQBTQ):kRF00R#8F_Do;HO
RSSQW.Bi:zuR0FkR8#0_oDFH
O;S1SR)RWm:kRF00R#8F_Do;HO
RSS7mqagF:Rk#0R0D8_FOoH;S
SRa7qmRU:FRk0#_08DHFoOS;
SqR7a:m(R0FkR8#0_oDFH
O;S7SRqnam:kRF00R#8F_Do;HO
RSS7mqa6F:Rk#0R0D8_FOoH;S
SRa7qmRc:FRk0#_08DHFoOS;
SqR7a:mdR0FkR8#0_oDFH
O;S7SRq.am:kRF00R#8F_Do;HO
RSS7mqa4F:Rk#0R0D8_FOoH;S
SRa7qm:jRR0FkR8#0_oDFH
O;S1SRB:pmR0FkR8#0_oDFH
O;S1SRB pmRF:Rk#0R0D8_FOoH;S
SRq17mF:Rk#0R0D8_FOoH;S
SRq17m: RR0FkR8#0_oDFH
O;SaSRXwwQmvq uRaY:kRF00R#8F_Do;HO
RSSaQXwwvm u:aYR0FkR8#0_oDFH
O;SaSRXwwQmpwzpF:Rk#0R0D8_FOoH;S
SRw)XQqwmwpzp:kRF00R#8F_Do;HO
RSS)QXwwzmwpRp:FRk0#_08DHFoOS;
SXR)wmQw avuYF:Rk#0R0D8_FOoH;S
SR7v)BpvuRF:Rk#0R0D8_FOoH
;S2SCR
MB8Rmmvuha h;B

mmvuha hR_1Ap7 7qu_QR
RRSbSSF5s0
SSSumWvzRaj:kRF00R#8F_Do;HOSS
SSvuWm4zaRF:Rk#0R0D8_FOoH;S
SSvuWm.zaRF:Rk#0R0D8_FOoH;S
SS7p 7Rmh:kRF00R#8F_Do;HORS
SS7p 7:B1H#MR0D8_FOoH;S
SS7p 7iBp:RHM#_08DHFoOS;
S Sp7q77aH(:M0R#8F_Do;HO
SSSp7 77nqa:RHM#_08DHFoOS;
S Sp7q77aH6:M0R#8F_Do;HO
SSSp7 77cqa:RHM#_08DHFoOS;
S Sp7q77aHd:M0R#8F_Do;HO
SSSp7 77.qa:RHM#_08DHFoOS;
S Sp7q77aH4:M0R#8F_Do;HO
SSSp7 77jqa:RHM#_08DHFoOS;
S Sp777q7:)dH#MR0D8_FOoH;S
SS7p 77q7)H.:M0R#8F_Do;HO
SSSp7 7q)774M:HR8#0_oDFH
O;SpSS q777j7):RHM#_08DHFoOS;
S Sp7 77hM:HR8#0_oDFH
O;SpSS  77XH :M0R#8F_Do;HO
SSSp7 7):1aH#MR0D8_FOoH
SSSS
2;CRM8Bumvmhh a
R;
vBmu mhhRaR1QA_)j6j_e7)
ht  B)QRS5
RBRRz ))hva_mR7 :s#0HRMo:"=Rj"Lj;R
SR)RQ6_jjB)z) Rha:s#0HRMo:"=RjjLjjjjjjjjjj
j"2b;
FRs05)
Qp  7hH:RM0R#8F_Do;HO
uQ)WRv:H#MR0D8_FOoH;z
B)h) :MRHR8#0_oDFH
O;Q )p7R4:FRk0#_08DHFoOQ;
)7p .F:Rk#0R0D8_FOoH
2RR;M
C8FROlMbFC;M0
B

mmvuha hRAR1_A)t_
Qub0FsRB5
pRi:H#MR0D8_FOoH;1
)aH:RM0R#8F_Do;HO
)uqqmv1iH:RM0R#8F_Do;HO
A)tBmmp)H:RM0R#8F_Do_HOP0COF5sRdFR8IFM0R;j2R)
AQat]h1 1:MRHR8#0_oDFHPO_CFO0sdR5RI8FMR0FjR2;
 A)q)a]q:vuRRHM#_08DHFoOC_POs0FRR5d8MFI0jFR2
;RAhpQia)q H:RM0R#8F_Do_HOP0COF5sRdFR8IFM0R;j2R 
)7vuW:kRF00R#8F_Do;HO
 t) Whuvk:F00R#8F_Do;HO
zAp vuW:0FkR8#0_oDFHRO
R
2;CRM8ObFlFMMC0
;
ObFlFMMC0AR1__QmQ
dBRRRRRRRRRCRoMHCsORR5u_Qha YuRRRR:HRL0C_POs0F5RR6RI8FMR0Fj
2;RRRRRRRRRRRRRRRRRRRRupzpzRuRRL:RH:0R=jR''
;RSRSRR RWqui_zzppuRR:LRH0:'=Rj
';RRRRRRRRRRRRRRRRRRRRh_ tat)QtR ):HRL0=R:R''jR
;RRRRRRRRRRRRRRRRRRRRRQ1m_a7qhqR)7:0R#soHMR":=1pA_emBv1R"
RRRRRRRRRRRRRRRRR;2R
RRRRRRRRbRRF5s0RR
RRRRRRRRRRRRRRqRuBtiq Q_uhRRRRRRRRH:RM0FkR8#0_oDFH;OR
RRRRRRRRRRRRRRRRapqBQ]_hauz_peqzR R:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRpRBm_Bi AhqpR RRRRRRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRRQRRhauz_iBpRRRRRRRRRRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRRmuzazBa_pRiRRRRRR:RRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRamzu_za AhqpR RRRRR:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRR_R7m_za4RRRRRRRRRRRRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRR7RR_amz_RjRRRRRRRRRRRR:HRMR#_08DHFoO
R;SSRRu z_hSASR:RRRRHMR8#0_oDFH;OR
RSRSqW iz_u_A hSRRR:MRHR0R#8F_DoRHO;RR
RRRRRRRRRRRRR7RR__Qh4RRRRRRRRRRRRRR:FRk0#_08DHFoO
R;RRRRRRRRRRRRRRRR7h_Q_RjRRRRRRRRRR:RRR0FkR8#0_oDFHRORRRRRRRRRRRRRR
RRRRRRRRRRRRRRR2RR;M
C8FROlMbFC;M0RO

FFlbM0CMR_1A1qu)vn.6ibq
FRs05q
S7 7)1:1RRRHMR8#0_oDFHPO_CFO0s4R5dFR8IFM0R;j2
qS7ahqQRH:RM0R#8F_Do_HOP0COF5sR486RF0IMF2Rj;v
SqW1i)R h:MRHR8#0_oDFHPO_CFO0sR5d8MFI0jFR2S;
Wh) ,QB]up1  ,BaBBpmia,1qAh7Yp,1 , uu mW)wmwRH:RM0R#8F_Do;HO
qS7azqmaRR:FRk0R8#0_oDFHPO_CFO0s654RI8FMR0Fj22
;M
C8FROlMbFC;M0
m
Bvhum RhaR_1A7q pYj_6hb1
FRs05 
7pQqYhRR:H#MR0D8_FOoH; 
7pmqYz:aRR0FkR8#0_oDFH2O
;M
C8FROlMbFC;M0
m
Bvhum RhaR_1AwaQp 6)_j
h1b0FsRw5
Q pa)RQh:MRHR8#0_oDFH
O;waQp z)maRR:FRk0#_08DHFoO;
2
8CMRlOFbCFMM
0;
vBmu mhheaRBbB
FRs05R
Y:kRF00R#8F_Do
HO2C;
MO8RFFlbM0CM;B

mmvuha hR7th
sbF0
R5YRR:FRk0#_08DHFoO;
2
8CMRlOFbCFMM
0;
0
N0LsHkR0C#_$MLODN	F_LGVRFRDNDRO:RFFlbM0CMRRH#0Csk;0
N0LsHkR0C#_$MD_HLODCDRRFVNRDD:FROlMbFCRM0H0#Rs;kC
0N0skHL0LCRD	NO_GLF_8bN_MbHRRFV1QA_mp_7YRR:ObFlFMMC0#RHRq"uBtiq Q_uh
";Ns00H0LkCDRLN_O	L_FGb_N8bRHMF1VRAm_Q_BQdRO:RFFlbM0CMRRH#"Buqi qt_huQ"N;
0H0sLCk0RNLDOL	_FbG_Nb8_HFMRVAR1_uvQQX_a_qcph: RRlOFbCFMMH0R#7R"u7d,h7d,u7.,h7.,u74,h74,u7j,hBj,iBu,i;h"
0N0skHL0LCRD	NO_GLF_8bN_MbHRRFV1QA_m7_mRO:RFFlbM0CMRRH#"Buqi qtu"Qh;0
N0LsHkR0CLODN	F_LGN_b8H_bMVRFR_1A)_tA7R)e:FROlMbFCRM0H"#R)jtA,A)t4t,)A;."
0N0skHL0LCRD	NO_GLF_8bN_MbHRRFV1QA_))_7eRR:ObFlFMMC0#RHR)"Qp" 7;0
N0LsHkR0C)amz ]_a)tmz]q_wAB)QRRFV1pA_wBm1RO:RFFlbM0CMRRH#0Csk;0
N0LsHkR0C)amz ]_a)tmz]q_wAB)QRRFV1]A_wBm1RO:RFFlbM0CMRRH#0Csk;0
N0LsHkR0C1_7qQzhua _7p qY7VRFR_1AQR.B:FROlMbFCRM0H0#Rs;kC
0N0skHL01CR7mq_zzaua _7p qY7VRFR_1AQR.B:FROlMbFCRM0HV#RNCD#;0
N0LsHkR0C1_BpQzhuaQ_wp)a  F7RVAR1_BQ.RO:RFFlbM0CMRRH#V#NDCN;
0H0sLCk0RNLDOL	_FbG_Nb8_HFMRVAR1_)AqB m7_e7)RO:RFFlbM0CMRRH#")AqB m7"N;
0H0sLCk0RNLDOL	_FbG_Nb8_HFMRVAR1_A)tq)_7eRR:ObFlFMMC0#RHRt")A)j,t,A4).tA"N;
0H0sLCk0RNLDOL	_FbG_Nb8_HFMRVAR1_cQ)j7j_):eRRlOFbCFMMH0R#QR")7p "N;
0H0sLCk0RNLDOL	_FbG_Nb8_HFMRVAR1_6Q)j7j_):eRRlOFbCFMMH0R#QR")7p 4),Qp. 7"N;
0H0sLCk0Rq17_uQhz7a_ Ypq F7RVAR1_BQ._wwQmRR:ObFlFMMC0#RHRk0sCN;
0H0sLCk0Rq17_amzu_za7q pYR 7F1VRA._QBQ_ww:mRRlOFbCFMMH0R#NRVD;#C
0N0skHL0QCR.BB_p7i_Q7eQ F)RVAR1_BQ._wwQmRR:ObFlFMMC0#RHR
j;Ns00H0LkC.RQBQ_ww m_hFARVAR1_BQ._wwQmRR:ObFlFMMC0#RHRh" q Ap7
";Ns00H0LkC Ra11a_uv)qRRFV11A_uv)q.i6nqRR:ObFlFMMC0#RHR;""
8CMRvBmu mhh;a1








