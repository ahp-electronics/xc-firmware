-- $Header: //synplicity/maplat2018q2p1/mappers/att/lib/gen_orca5g/seq_srl.vhd#1 $
@ELDHs$NsR Q  k;
#QCR 3  #_08DHFoO4_4nNc3D
D;kR#CQ   38#0_oDFHkO_Mo#HM3C8N;DD
Ck#R Q  03#8F_Do_HON0sHED3NDD;
HNLssF$RsdON;#
kCsRFO3NdFNsOObFl3DND;C

M00H$ R1T)_1p#RH
oRRCsMCH
O5RRRRR8RN8Is_HE80RH:RMo0CC:sR=;R(
RRRRNRR8_8s#CHxRH:RMo0CC:sR=6Rn;R
RRRRR8H_I8R0E:MRH0CCos=R:R
U;RRRRRCRMoD_O	RR:LDFFCRNM:0=Rs;kC
RRRRHRR#M_HbRk0:FRLFNDCM=R:Rk0sCR;
RRRRR_H#Fbk0k:0RRFLFDMCNRR:=0Csk2R;
RsbF0R5
RRRRR7)q7:)RRRHM#_08DHFoOC_POs0F58N8sH_I8-0E4FR8IFM0R;j2
RRRR7RRqRaqR:RRRRHM#_08DHFoOC_POs0F5I8_HE80-84RF0IMF2Rj;R
RRRRRWR RRH:RM0R#8F_Do;HO
RRRRBRRpRiR:MRHR8#0_oDFH
O;RRRRR_Rq)R1aRH:RM0R#8F_Do;HO
RRRR1RR_a)1RRR:H#MR0D8_FOoH;R
RRRRR7amzRRRR:kRF00R#8F_Do_HOP0COF8s5_8IH04E-RI8FMR0Fj;22
8CMRT1 _p1);N

sHOE00COkRsCsHCo#s0C#VRFRT1 _p1)R
H#0C$bRD#s_sNsNH$R#sRNsRN$50jRF_R8I0H8E2-4RRFV#_08DHFoOC_POs0F58N8sH_#x4C-RI8FMR0Fj
2;#MHoNJDR_0HMR#:RsND_s$sN;C
Lo
HM
zRRjRR:HNV58_8s#CHxR4>R2CRoMNCs0RC
RzRR4RR:VRFsHMRHR0jRF_R8I0H8E4R-RMoCC0sNCR
RRRRRbOsFC5##B2pi
RRRRLRRCMoH
RSRRVRHRH5s#oHM_oC8Cp5BiR220MEC
RSRRHRRVWR5 RR='24'RC0EMS
SR_RJH5M0H<2R=JR5_0HM55H2Ns88_x#HCR-.8MFI0jFR2RR&7qqa52H2;R
SRRRRCRM8H
V;SRRRR8CMR;HV
RSRCRM8bOsFC;##
RSR7amz5RH2<J=R_0HM55H2OPFM_0HMCsoC57)q72)2;R
RRMRC8CRoMNCs0zCR4R;
R8CMRMoCC0sNCjRz;R

RRz.:VRH58N8sH_#x=CRRR42oCCMsCN0
RRRRRzd:FRVsRRHHjMRRR0F8H_I8R0E-o4RCsMCN
0CRRRRRsRbF#OC#p5BiR2
RRRRRoLCHRM
RRRRRHRRVsR5HM#Ho8_CoBC5p2i2RC0EMR
RRRRRRHRRVWR5 RR='24'RC0EMR
RRRRRRRRR7amz5RH2<7=Rq5aqH
2;RRRRRRRRR8CMR;HV
RRRRRRRR8CMR;HV
RRRRCRRMb8RsCFO#
#;RRRRCRM8oCCMsCN0R;zd
CRRMo8RCsMCNR0Cz
.;
8CMRosCHC#0s
#;
ONsECH0Os0kC0R#NO0H_D#sRRFV1_ T1R)pHV#
k0MOHRFMM_klODCD5:MRR0HMCsoC;#RH_bHMkR0,HF#_kk0b0RR:LDFFC2NMskC0sHMRMo0CCHsR#RRRRPR
NNsHLRDCPkNDCRR:HCM0o;Cs
sPNHDNLCkRMlC_so:#RR0HMCsoC;C
Lo
HMRkRMlC_so:#R=;Rj
HRRV#5H_bHMkR020MECRR
RRRRRM_kls#CoRR:=M_kls#CoR4+R;R
RCRM8H
V;RVRH5_H#Fbk0kR020MECRR
RRRRRRlMk_osC#=R:RlMk_osC#RR+4R;
R8CMR;HV
PRRNCDkRR:=5-MRRlMk_osC#42/nR;
R0sCkRsMPkNDCC;
MM8RkOl_C;DD
k
VMHO0FsMRCHlNMoHM_osC5RM:HCM0o;CsR_H#HkMb0H,R#k_F00bkRL:RFCFDNsM2Cs0kMMRH0CCos#RHRRRRRN
PsLHNDPCRNCDkRH:RMo0CC
s;PHNsNCLDRlMk_osC#RR:HCM0o;Cs
oLCHRM
RlMk_osC#=R:R
j;RNRPDRkC:j=R;R
RHHV5#M_Hb2k0RC0EMRR
RRRRRlMk_osC#=R:RlMk_osC#RR+4R;
R8CMR;HV
HRRV#5H_0Fkb2k0RC0EMRR
RRRRRkRMlC_so:#R=kRMlC_so+#RR
4;RMRC8VRH;R
RPkNDC=R:RR5M-kRMlC_soR#2sRCl4
n;RCRs0MksRDPNk
C;CRM8sNClHMMHoC_so
;
VOkM0MHFRN#0sM0HoC_so#5H_bHMk:0RRFLFDMCN2CRs0MksR0HMCsoCR
H#LHCoMR
RHHV5#M_Hb2k0RC0EMR
RRRRRskC0s4MR;R
RCRM8H
V;RCRs0MksR
j;CRM8#s0N0oHM_osC;V

k0MOHRFMbVsCHoG_CHM5#k_F00bkRL:RFCFDNRM2skC0s#MR0MsHo#RH
oLCHRM
R5HVHF#_kk0b002RE
CMRRRRRCRs0MksRa"pa
";RMRC8VRH;R
RskC0s"MRp"wa;M
C8sRbCGVH_MoC;O

F0M#NRM0M_kl#_sDODCD#RR:HCM0oRCs:M=RkOl_C5DDNs88_x#HCH,R#M_Hb,k0R_H#Fbk0k;02
MOF#M0N0kRMl	_#Hsb_CRo#:MRH0CCos=R:RlsCNHHMMso_CNo58_8s#CHx,#RH_bHMkR0,HF#_kk0b0
2;O#FM00NMRlMk_N#0ss0_C:oRR0HMCsoCRR:=#s0N0oHM_osC5_H#HkMb0
2;O#FM00NMRD#s_CbsVRHG:0R#soHMRR:=bVsCHoG_CHM5#k_F00bk2
;
#MHoNDDR#:LRR8#0_oDFHPO_CFO0sR5d8MFI0jFR2=R:Rj"jj;j"
b0$C#RRs0D_lNb_s$sNRRH#NNss$jR5RR0F5lMk_D#s_DOCD+#RR242RRFV#_08DHFoOC_POs0F5I8_HE80R4-RRI8FMR0Fj
2;
o#HMRND0_lbNNss$RR:#_sD0_lbNNss$#;
HNoMDlR0b8_N8:sRR8#0_oDFHPO_CFO0s85N8Is_HE80-84RF0IMF2Rj;H
#oDMNRb0l_0Fk_8N8sRR:#_08DHFoOC_POs0F5I8_HE80-84RF0IMF2Rj;N

0H0sLCk0R#\3sFD_VCV#0:\RRs#0H;Mo
C
Lo
HM
Rzj:VRHR_H#HkMb0CRoMNCs0
CRRsRbF#OC#p5BiR2
RoLCHRM
RHRRVsR5HM#Ho8_CoBC5p2i2RC0EMR
RRRRRH5VRW= RR''42ER0CRM
RRRRR0RRlNb_s$sN5Rj2<7=Rq;aq
RRRRCRRMH8RVR;
RCRRMH8RVR;
R8CMRFbsO#C#;CR
Mo8RCsMCN;0C
j
z4RR:HMVRFH05#M_Hb2k0RMoCC0sNCRR
RRRRR0RRlNb_s$sN5Rj2<7=Rq;aq
8CMRMoCC0sNC
;

4
z:VRHR8N8sH_I8R0E<c=RRMoCC0sNCR
RRCRLo
HMS#SDL=R<RhBmea_17m_pt_QBea BmM)5k#l_	_Hbs#CoR4-R,2Rc;R
RRRRRR4Rz4RR:VRFsHMRHR0jRF8R5_8IH0-ER4o2RCsMCN
0CSNSS0H0sLCk0R#\3sFD_VCV#0F\RV4Rz4:4RRLDNCHDR#sR#Ds_bCGVHRH&RMo0CCHs'lCNo5I8_HE802RR&"R7"&MRH0CCosl'HN5oCM_kl#s0N0C_so&2RR""WRH&RMo0CCHs'lCNo5RH2& R""RR&HCM0o'CsHolNCk5Ml0_#N_s0sRCo+kRMl	_#Hsb_C2o#R"&RX&"RR0HMCsoC'NHloHC5R4+R2S;
SCSLo
HMRRRRRRRRRRRRz444:]R1Q4wanR
RRRRRRRRRRFRbsl0RN
b5RRRRRRRRRRRRRRRRqR7j=D>R#jL52R,
RRRRRRRRRRRRRqRR7=4R>#RDL254,R
RRRRRRRRRRRRRR7Rq.>R=RLD#5,.2
RRRRRRRRRRRRRRRRdq7RR=>D5#Ld
2,RRRRRRRRRRRRRRRRB= R> RW,R
RRRRRRRRRRRRRRpRBi>R=RiBp,R
RRRRRRRRRRRRRR)R1Q>R=Rb0l_sNsNj$5225H,R
RRRRRRRRRRRRRRmR7RR=>0_lbNNss$2545
H2RRRRRRRRRRRR2R;
RRRRRCRRMo8RCsMCNR0Cz;44
RRRRRRRR.z4RH:RV#RH_0FkbRk0oCCMsCN0RR
RRRRRRsRbF#OC#D5O	R2
RRRRRRRRRLRRCMoH
RRRRRRRRRRRRRRRRRHV5#sHH_MoCC8o5iBp202RE
CMRRRRRRRRRRRRRRRRRRRRH5VRW= RR''42ER0CRM
RRRRRRRRRRRRRRRRRRRRR7RRmRza<0=RlNb_s$sN5;42
RRRRRRRRRRRRRRRRRRRR8CMR;HV
RRRRRRRRRRRRRRRR8CMR;HV
RRRRRRRRRRRR8CMRFbsO#C#;RR
RRRRRCRRMo8RCsMCN;0C
RRRRRRRRdz4RH:RVFRM0#5H_0Fkb2k0RMoCC0sNCS
SRRRR7amzRR<=0_lbNNss$254;R
RRRRRRMRC8CRoMNCs0zCR4
d;CRM8oCCMsCN0R;z4
.
z:VRHR8N8sH_I8R0E>RRcoCCMsCN0
RRRRoLCHRM
RRRRR
RRRRRRRRRRzR..:FRVsRRHH4MRRR0F5lMk_D#s_DOCDR#2oCCMsCN0RR
RRRRRRRRRR.Rz.R4:VRFs[MRHR0jRF8R5_8IH0-ER4o2RCsMCN
0CSNSS0H0sLCk0R#\3sFD_VCV#0F\RV.Rz.:.RRLDNCHDR#pR"wRa"&MRH0CCosl'HN5oC8H_I820ER"&R7&"RR0HMCsoC'NHloMC5k#l_00Ns_osCR5+RHRR-442*n&2RR""WRH&RMo0CCHs'lCNo5R[2& R""RR&HCM0o'CsHolNCk5Ml0_#N_s0sRCo+*RH4Rn2&XR""RR&HCM0o'CsHolNCR5[+2R4;R
RRRRRRRRRRCRLo
HMRRRRRRRRRRRRRRRRz...:]R1Q4wanR
RRRRRRRRRRRRRRFRbsl0RN
b5RRRRRRRRRRRRRRRRqR7j=4>''R,
RRRRRRRRRRRRRqRR7=4R>4R''R,
RRRRRRRRRRRRRqRR7=.R>4R''R,
RRRRRRRRRRRRRqRR7=dR>4R''R,
RRRRRRRRRRRRRBRR >R=R,W 
RRRRRRRRRRRRRRRRiBpRR=>B,pi
RRRRRRRRRRRRRRRRQ1)RR=>0_lbNNss$R5H-2R45,[2
RRRRRRRRRRRRRRRRR7m=0>RlNb_s$sN55H2[R2
RRRRRRRRR2RR;S
SSR
RRRRRRRRRRRRRRRRRRRR
RRRRRRRRRCRRMo8RCsMCNR0CR.z.4S;
S6Sz:VRH5lMk_H#	bC_so=#RRRj2oCCMsCN0RS
SSlS0bk_F08_N8<sR=lR0bs_Ns5N$M_kl#_sDODCD#
2;SCSSMo8RCsMCNR0Cz
6;RRRRRRRRCRM8oCCMsCN0R.z.;R
RRRRRRRR
RRRRRzRR.R.d:VRH5lMk_H#	bC_so/#R=2RjRMoCC0sNCSR
S#SDL=R<RhBmea_17m_pt_QBea BmM)5k#l_	_Hbs#CoR4-R,2Rc;R
RRRRRRRRRR.Rz.Rc:VRFs[MRHR0jRF8R5_8IH0-ER4o2RCsMCN
0CSNSS0H0sLCk0R#\3sFD_VCV#0F\RV.Rz.:.RRLDNCHDR#sR#Ds_bCGVHRH&RMo0CCHs'lCNo5I8_HE802RR&"R7"&MRH0CCosl'HN5oCM_kl#s0N0C_soRR+M_kl#_sDODCD#n*42RR&"RW"&MRH0CCosl'HN5oC[&2RR"" RH&RMo0CCHs'lCNo5lMk_N#0ss0_C+oRRlMk_D#s_DOCD4#*nRR+M_kl#b	H_osC#&2RR""XRH&RMo0CCHs'lCNo5+[RR;42
RRRRRRRRRRRRoLCHRM
RRRRRRRRRRRRRzRR.:..RQ1]wna4
RRRRRRRRRRRRRRRRsbF0NRlbR5
RRRRRRRRRRRRRqRR7=jR>#RDL25j,R
RRRRRRRRRRRRRR7Rq4>R=RLD#5,42
RRRRRRRRRRRRRRRR.q7RR=>D5#L.
2,RRRRRRRRRRRRRRRRqR7d=D>R#dL52R,
RRRRRRRRRRRRRBRR >R=R,W 
RRRRRRRRRRRRRRRRiBpRR=>B,pi
RRRRRRRRRRRRRRRRQ1)RR=>0_lbNNss$k5Mls_#DC_OD2D#5,[2
SRRSRRRRR7m=0>RlNb_s$sN5lMk_D#s_DOCD+#RR542[R2
RRRRRRRRR2RR;S
SSR
RRRRRRRRRRMRC8CRoMNCs0RCRzc..;S
SSb0l_0Fk_8N8s=R<Rb0l_sNsNM$5k#l_sOD_C#DDR4+R2R;
RRRRRCRRMo8RCsMCNR0Czd..;R
RRRRRR.RzdRR:HHVR#k_F00bkRMoCC0sNCRR
RRRRRbRRsCFO#O#5D
	2RRRRRRRRRRRRLHCoMR
RRRRRRRRRRRRRRVRHRH5s#oHM_oC8Cp5BiR220MEC
RRRRRRRRRRRRRRRRRRRRRHV5RW =4R''02RE
CMRRRRRRRRRRRRRRRRRRRRRRRR7amzRR<=0_lbF_k0Ns88;R
RRRRRRRRRRRRRRRRRRMRC8VRH;R
RRRRRRRRRRRRRRMRC8VRH;R
RRRRRRRRRRMRC8sRbF#OC#
;RRRRRRRRRCRM8oCCMsCN0;R
RRRRRR.RzcRR:HMVRFH05#k_F00bk2CRoMNCs0SC
SRRRRz7ma=R<Rb0l_0Fk_8N8sR;
RRRRRCRRMo8RCsMCNR0Cz;.c
8CMRMoCC0sNC.Rz;C

MN8RsHOE00COkRsC#00NH#O_s
D;
s
NO0EHCkO0s#CRCODC0s_#DVRFRT1 _p1)R
H#VOkM0MHFRlMk_DOCDR5M:MRH0CCosH;R#M_Hb,k0R_H#Fbk0k:0RRFLFDMCN20sCkRsMHCM0oRCsHR#RR
RRPHNsNCLDRDPNk:CRR0HMCsoC;N
PsLHNDMCRksl_CRo#:MRH0CCosL;
CMoH
MRRksl_CRo#:M=R;R
RPkNDC=R:RlMk_osC#n/4;R
RH5VRMCRslnR4RR/=j02RE
CMRRRRPkNDC=R:RDPNk+CRR
4;RMRC8VRH;R
RskC0sPMRNCDk;M
C8kRMlC_OD
D;VOkM0MHFR0oC_8CM_b8C0#E5HRxC:MRH0CCosRR;80CbERR:HCM0o2CsR0sCkRsMHCM0oRCsHP#
NNsHLRDCl_HM#CHxRH:RMo0CC:sR=;Rj
oLCHRM
RMlH_x#HC=R:Rb8C0
E;RVRHRH5#x<CRRb8C0RE20MEC
RRRRMlH_x#HC=R:Rx#HCR;
R8CMR;HV
sRRCs0kMHRlMH_#x
C;CRM8o_C0C_M880CbE
;
O#FM00NMRlMk_D#s_DOCD:#RR0HMCsoCRR:=M_klODCD58N8sH_#xRC,HH#_M0bk,#RH_0Fkb2k0;#

HNoMD#RDLRR:#_08DHFoOC_POs0F58dRF0IMF2RjRR:="jjjj
";0C$bRsR#Dl_0bs_NsRN$HN#Rs$sNRR5j0MFRk#l_sOD_C#DDR4+R2VRFR8#0_oDFHPO_CFO0s_58I0H8ERR-4FR8IFM0R;j2
H
#oDMNRb0l_sNsN:$RRD#s_b0l_sNsN
$;#MHoN0DRl8b__sNsN:$RRD#s_b0l_sNsN
$;
0N0skHL0\CR3D#s_VFV#\C0R#:R0MsHo
;
LHCoM0

lNb_s$sN5Rj2<7=Rq;aq
4
z:VRHR8N8sH_I8R0E<c=RRMoCC0sNCR
RRCRLo
HMRRRRRRRRD5#LNs88_8IH0-ERR84RF0IMF2RjRR<=)7q7)R;
RRRRRzRR4:4RRsVFRHHRMRRj05FR8H_I8R0E-R42oCCMsCN0
SSSNs00H0LkC3R\#_sDF#VVCR0\FzVR4R44:NRDLRCDH"#R)"waRH&RMo0CCHs'lCNo5I8_HE802RR&"R7"&MRH0CCosl'HN5oCj&2RR""WRH&RMo0CCHs'lCNo5RH2& R""RR&HCM0o'CsHolNC85N8#s_H2xCR"&RX&"RR0HMCsoC'NHloHC5R4+R2S;
SCSLo
HMRRRRRRRRRRRRz444:]R1Q4wanR
RRRRRRRRRRFRbsl0RN
b5RRRRRRRRRRRRRRRRqR7j=D>R#jL52R,
RRRRRRRRRRRRRqRR7=4R>#RDL254,R
RRRRRRRRRRRRRR7Rq.>R=RLD#5,.2
RRRRRRRRRRRRRRRRdq7RR=>D5#Ld
2,RRRRRRRRRRRRRRRRB= R> RW,R
RRRRRRRRRRRRRRpRBi>R=RiBp,R
RRRRRRRRRRRRRR)R1Q>R=Rb0l_sNsNj$5225H,R
RRRRRRRRRRRRRRmR7RR=>0_lbNNss$2545
H2RRRRRRRRRRRR2R;
RRRRRCRRMo8RCsMCNR0Cz;44
7SSmRza<0=RlNb_s$sN5;42
8CMRMoCC0sNC4Rz;z

.H:RV8RN8Is_HE80Rc>RRMoCC0sNCR
RRCRLo
HMRRRRRRRRDR#L<)=Rq)7758dRF0IMF2Rj;R
RRRRRR.Rz.RR:VRFsHMRHR04RFMR5k#l_sOD_C#DD2CRoMNCs0
CRRRRRRRRRRRRRz4..:FRVsRR[HjMRRR0F5I8_HE80R2-4RMoCC0sNCS
SS0N0skHL0\CR3D#s_VFV#\C0RRFVz4..RD:RNDLCRRH#"a)w"RR&HCM0o'CsHolNC_58I0H8E&2RR""7RH&RMo0CCHs'lCNo5R5H-2R4*24nR"&RW&"RR0HMCsoC'NHlo[C52RR&"R "&MRH0CCosl'HN5oCo_C0C_M880CbE85N8#s_H,xCR4H*nR22&XR""RR&HCM0o'CsHolNCR5[+2R4;S
SS0N0skHL0\CR3D#s_VFV#\C0RRFVz...RD:RNDLCRRH#"a)w"RR&HCM0o'CsHolNC_58I0H8E&2RR""7RH&RMo0CCHs'lCNo5R5H-2R4*24nR"&RW&"RR0HMCsoC'NHlo[C52RR&"R "&MRH0CCosl'HN5oCo_C0C_M880CbE85N8#s_H,xCR4H*nR22&XR""RR&HCM0o'CsHolNCR5[+2R4;R
RRRRRRRRRRCRLo
HMRRRRRRRRRRRRRRRRz4..:]R1Q4wanR
RRRRRRRRRRRRRRFRbsl0RN
b5RRRRRRRRRRRRRRRRqR7j='>R4
',RRRRRRRRRRRRRRRRqR74='>R4
',RRRRRRRRRRRRRRRRqR7.='>R4
',RRRRRRRRRRRRRRRRqR7d='>R4
',RRRRRRRRRRRRRRRRB= R> RW,R
RRRRRRRRRRRRRRpRBi>R=RiBp,R
RRRRRRRRRRRRRR)R1Q>R=Rb0l_sNsNH$5R4-R225[,R
RRRRRRRRRRRRRRmR7RR=>0_lbNNss$25H5
[2RRRRRRRRRRRR2R;
RRRRRRRRRRRRRzRR.:..RQ1]wna4
RRRRRRRRRRRRRRRRsbF0NRlbR5
RRRRRRRRRRRRRqRR7=jR>#RDL25j,R
RRRRRRRRRRRRRR7Rq4>R=RLD#5,42
RRRRRRRRRRRRRRRR.q7RR=>D5#L.
2,RRRRRRRRRRRRRRRRqR7d=D>R#dL52R,
RRRRRRRRRRRRRBRR >R=R,W 
RRRRRRRRRRRRRRRRiBpRR=>B,pi
RRRRRRRRRRRRRRRRQ1)RR=>0_lbNNss$R5H-2R45,[2
RRRRRRRRRRRRRRRRR7m=0>Rl8b__sNsNH$5R4-R225[
RRRRRRRRRRRR
2;RRRRRRRRRRRRRRRRRRRR
RRRRRRRRRRRR8CMRMoCC0sNCzRR.;.4
RRRRRRRR8CMRMoCC0sNC.Rz.S;
Sz7ma=R<Rb0l_N8_s$sN5MOFPM_H0CCosq5)757)Ns88_8IH0-ERR84RF0IMF2Rc2
2;CRM8oCCMsCN0R;z.
M
C8sRNO0EHCkO0s#CRCODC0s_#D
;

