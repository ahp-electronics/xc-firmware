--
@ER--B$FbsEHo0OR52gR4g-cRRj.jd$R1MHbDO$H0ROQM
R--fN]C8:CsR#//$DMbH0OH$N/lb0DN.Uj4J4.b/blNb#Cs/DGHH/MGD/HLoCCMs/HOo_CMoCCMs/HOs_NlsPI3E48yR-f
-D

HNLssH$RC;CC
Ck#RCHCC03#8F_Do_HO4c4n3DND;#
kCCRHC#C30D8_FOoH_o#HM3C8N;DD
LDHs$NsRHkM#;Hl
Ck#RHkM#3HlPlOFbCFMM30#N;DD
0CMHR0$Xv)q4X.U4H1R#R
Rb0FsRR5
RRRRRmRRR:RRR0FkR8#0_FkDo;HO
R
RRRRRRjRqR:RRRRHM#_08koDFH
O;RRRRRRRRqR4RRH:RM0R#8D_kFOoH;R
RRRRRR.RqR:RRRRHM#_08koDFH
O;RRRRRRRRqRdRRH:RM0R#8D_kFOoH;R
RRRRRRcRqR:RRRRHM#_08koDFH
O;RRRRRRRRqR6RRH:RM0R#8D_kFOoH;S
SqRnRRH:RM0R#8D_kFOoH;R
RRRRRRRR7RRR:H#MR0k8_DHFoOR;
RRRRRWRRBRpi:MRHR8#0_FkDo;HO
RRRRRRRRRW RRR:H#MR0k8_DHFoOR
RRRRRR
2;CRM8Xv)q4X.U4
1;
ONsECH0Os0kCqR)vR_eFXVR)4qv.4UX1#RH
o#HMRND0Rj,0:4RR8#0_FkDo;HO
o#HMRNDI,C4R.ICR#:R0k8_DHFoOL;
CMoH
RRRRRRRRRRRR)XzqcvnR):RqcvnXR41
RRRRRRRRRRRRRRRRsbF0NRlb7R5RR=>7q,Rj>R=R,qjRRq4=q>R4q,R.>R=R,q.
RRRRRRRRRRRRRRRRRRRRRRRRqRRd>R=R,qdRRqc=q>Rcq,R6>R=R,q6
SSSSRSSRRW =I>RCR4,WiBpRR=>WiBp,RRm=0>Rj
2;RRRRRRRRRRRRX)4zqcvnR):RqcvnXR41
RRRRRRRRRRRRRRRRsbF0NRlb7R5RR=>7q,Rj>R=R,qjRRq4=q>R4q,R.>R=R,q.
RRRRRRRRRRRRRRRRRRRRRRRRqRRd>R=R,qdRRqc=q>Rcq,R6>R=R,q6
SSSSRSSRRW =I>RCR.,WiBpRR=>WiBp,RRm=0>R4
2;m=R<RR0jIMECRRqn=jR''DRC#0CR4I;
C<4R= RWR8NMR0MF52qn;C
I.=R<RRW NRM8q
n;
8CMRv)q_
e;
H
DLssN$CRHC
C;kR#CHCCC38#0_oDFH4O_43ncN;DD
Ck#RCHCC03#8F_Do_HO#MHoCN83D
D;DsHLNRs$k#MHH
l;kR#Ck#MHHPl3ObFlFMMC0N#3D
D;CHM00X$R)nqvc1X.R
H#RFRbs50R
RRRRRRRRRmjRRR:FRk0#_08koDFH
O;RRRRRRRRmR4RRF:Rk#0R0k8_DHFoO
;
RRRRRRRRqRjRRH:RM0R#8D_kFOoH;R
RRRRRR4RqR:RRRRHM#_08koDFH
O;RRRRRRRRqR.RRH:RM0R#8D_kFOoH;R
RRRRRRdRqR:RRRRHM#_08koDFH
O;RRRRRRRRqRcRRH:RM0R#8D_kFOoH;R
RRRRRR6RqR:RRRRHM#_08koDFH
O;RRRRRRRR7RjRRH:RM0R#8D_kFOoH;R
RRRRRR4R7R:RRRRHM#_08koDFH
O;RRRRRRRRWiBpRH:RM0R#8D_kFOoH;R
RRRRRR RWR:RRRRHM#_08koDFHRO
RRRRR;R2
8CMRqX)vXnc.
1;
ONsECH0Os0kCqR)vXnc.e1_RRFVXv)qn.cX1#RH
oLCHRM
RRRRRRRRRXRRzv)qn:cRRv)qn4cX1RR
RRRRRRRRRRRRRbRRFRs0lRNb5=7R>jR7,jRqRR=>qRj,q=4R>4Rq,.RqRR=>q
.,RRRRRRRRRRRRRRRRRRRRRRRRRdRqRR=>qRd,q=cR>cRq,6RqRR=>q
6,SSSSSRSRW= R> RW,BRWp=iR>BRWpRi,m>R=R2mj;R
RRRRRRRRRR4RXzv)qn:cRRv)qn4cX1RR
RRRRRRRRRRRRRbRRFRs0lRNb5=7R>4R7,jRqRR=>qRj,q=4R>4Rq,.RqRR=>q
.,RRRRRRRRRRRRRRRRRRRRRRRRRdRqRR=>qRd,q=cR>cRq,6RqRR=>q
6,SSSSSRSRW= R> RW,BRWp=iR>BRWpRi,m>R=R2m4;M
C8qR)vXnc.e1_;D

HNLssH$RC;CC
Ck#RCHCC03#8F_Do_HO4c4n3DND;#
kCCRHC#C30D8_FOoH_o#HM3C8N;DD
LDHs$NsRHkM#;Hl
Ck#RHkM#3HlPlOFbCFMM30#N;DD
0CMHR0$Xv)qdU.X1#RH
bRRFRs05S
SmRR:FRk0#_08DHFoOC_POs0F5RR(8MFI0jFR2R;
RRRRRqRRjRRR:MRHR8#0_FkDo;HO
RRRRRRRRRq4RRR:H#MR0k8_DHFoOR;
RRRRRqRR.RRR:MRHR8#0_FkDo;HO
RRRRRRRRRqdRRR:H#MR0k8_DHFoOR;
RRRRRqRRcRRR:MRHR8#0_FkDo;HO
RRRRRRRRR7RRRR:H#MR0D8_FOoH_OPC0RFs5RR(8MFI0jFR2R;
RRRRRWRRBRpi:MRHR8#0_FkDo;HO
RRRRRRRRRW RRR:H#MR0k8_DHFoOR
RRRRRR
2;CRM8Xv)qdU.X1
;
NEsOHO0C0CksRv)q_FeRV)RXq.vdXRU1HL#
CMoH
RRRRRRRRRRRR)Xzq:vRRv)qd..X1RR
RRRRRRRRRRRRRbRRFRs0lRNb5R7j=7>R5,j2R=74>5R74R2,q=jR>jRq,4RqRR=>qR4,q=.R>.Rq,R
RRRRRRRRRRRRRRRRRRRRRRRRRq=dR>dRq,cRqRR=>qRc,
SSSSRSSRRW =W>R W,RBRpi=W>RB,piRRmj=m>R5,j2RRm4=m>R5242;R
RRRRRRRRRR4RXzv)qR):Rq.vdXR.1
RRRRRRRRRRRRRRRRsbF0NRlb7R5j>R=R.7527,R4R=>725d,jRqRR=>qRj,q=4R>4Rq,.RqRR=>q
.,RRRRRRRRRRRRRRRRRRRRRRRRRdRqRR=>qRd,q=cR>cRq,S
SSSSSR RWRR=>WR ,WiBpRR=>WiBp,jRmRR=>m25.,4RmRR=>m25d2R;
RRRRRRRRRXRR.qz)vRR:)dqv.1X.RR
RRRRRRRRRRRRRRFRbsl0RN5bR7=jR>5R7cR2,7>4=R6752q,Rj>R=R,qjRRq4=q>R4q,R.>R=R,q.
RRRRRRRRRRRRRRRRRRRRRRRRqRRd>R=R,qdRRqc=q>RcS,
SSSSSWRR >R=R,W RpWBi>R=RpWBim,Rj>R=Rcm52m,R4>R=R6m52
2;RRRRRRRRRRRRX)dzq:vRRv)qd..X1RR
RRRRRRRRRRRRRbRRFRs0lRNb5R7j=7>R5,n2R=74>5R7(R2,q=jR>jRq,4RqRR=>qR4,q=.R>.Rq,R
RRRRRRRRRRRRRRRRRRRRRRRRRq=dR>dRq,cRqRR=>q
c,SSSSSRSRW= R> RW,BRWp=iR>BRWpRi,m=jR>5RmnR2,m=4R>5Rm(;22
8CMRv)q_
e;DsHLNRs$HCCC;#
kCCRHC#C30D8_FOoH_n44cD3NDk;
#HCRC3CC#_08DHFoOH_#o8MC3DND;H
DLssN$MRkHl#H;#
kCMRkHl#H3FPOlMbFC#M03DND;C

M00H$)RXq.vdXRc1HR#
RsbF0
R5RRRRSRmj:kRF00R#8D_kFOoH;R
RRmRS4RR:FRk0#_08koDFH
O;RRRRSRm.:kRF00R#8D_kFOoH;R
RRmRSdRR:FRk0#_08koDFH
O;
RRRRRRRRRqjRRR:H#MR0k8_DHFoOR;
RRRRRqRR4RRR:MRHR8#0_FkDo;HO
RRRRRRRRRq.RRR:H#MR0k8_DHFoOR;
RRRRRqRRdRRR:MRHR8#0_FkDo;HO
RRRRRRRRRqcRRR:H#MR0k8_DHFoOR;
RSRR7RjRRH:RM0R#8D_kFOoH;R
RR7RS4RRR:MRHR8#0_FkDo;HO
RRRR.S7R:RRRRHM#_08koDFH
O;RRRRSR7dRRR:H#MR0k8_DHFoOR;
RRRRRWRRBRpi:MRHR8#0_FkDo;HO
RRRRRRRRRW RRR:H#MR0k8_DHFoOR
RRRRRR
2;CRM8Xv)qdc.X1
;
NEsOHO0C0CksRv)q_FeRV)RXq.vdXRc1HL#
CMoH
RRRRRRRRRRRR)Xzq:vRRv)qd..X1RR
RRRRRRRRRRRRRbRRFRs0lRNb5R7j=7>Rj7,R4R=>7R4,q=jR>jRq,4RqRR=>qR4,q=.R>.Rq,R
RRRRRRRRRRRRRRRRRRRRRRRRRq=dR>dRq,cRqRR=>qRc,
SSSSRSSRRW =W>R W,RBRpi=W>RB,piRRmj=m>Rjm,R4>R=R2m4;R
RRRRRRRRRR4RXzv)qR):Rq.vdXR.1
RRRRRRRRRRRRRRRRsbF0NRlb7R5j>R=R,7.R=74>dR7,jRqRR=>qRj,q=4R>4Rq,.RqRR=>q
.,RRRRRRRRRRRRRRRRRRRRRRRRRdRqRR=>qRd,q=cR>cRq,S
SSSSSR RWRR=>WR ,WiBpRR=>WiBp,jRmRR=>mR.,m=4R>dRm2C;
M)8Rqev_;H
DLssN$CRHC
C;kR#CHCCC38#0_oDFH4O_43ncN;DD
Ck#RCHCC03#8F_Do_HO#MHoCN83D
D;DsHLNRs$k#MHH
l;kR#Ck#MHHPl3ObFlFMMC0N#3D
D;
0CMHR0$Xv)q4UnX1#RH
bRRFRs05S
SmRR:FRk0#_08DHFoOC_POs0FR(5RRI8FMR0Fj
2;RRRRRRRRqRjRRH:RM0R#8D_kFOoH;R
RRRRRR4RqR:RRRRHM#_08koDFH
O;RRRRRRRRqR.RRH:RM0R#8D_kFOoH;R
RRRRRRdRqR:RRRRHM#_08koDFH
O;RRRRRRRR7RRRRH:RM0R#8F_Do_HOP0COF5sRR8(RF0IMF2Rj;R
RRRRRRBRWp:iRRRHM#_08koDFH
O;RRRRRRRRWR RRH:RM0R#8D_kFOoH
RRRRRRR2C;
MX8R)4qvn1XU;N

sHOE00COkRsC)_qveVRFRqX)vX4nUH1R#C
Lo
HMRRRRRRRRRRRRXqz)vRR:)4qvn1XcRR
RRRRRRRRRRRRRRFRbsl0RN5bR7=jR>5R7jR2,7>4=R47527,R.>R=R.7527,Rd>R=Rd752
,RSSSSRRRRRRRRRjRqRR=>qRj,q=4R>4Rq,.RqRR=>qR.,q=dR>dRq,SR
SSSSSWRR >R=R,W RpWBi>R=RpWBi
,RSSSSSRSRm=jR>5RmjR2,m=4R>5Rm4R2,m=.R>5Rm.R2,m=dR>5Rmd;22
RRRRRRRRRRRRzX4)Rqv:qR)vX4nc
1RRRRRRRRRRRRRRRRRb0FsRblNRj57RR=>725c,4R7=7>R5,62RR7.=7>R5,n2RR7d=7>R5,(2RS
SSRSRRRRRRRRRq=jR>jRq,4RqRR=>qR4,q=.R>.Rq,dRqRR=>qRd,
SSSSRSSRRW =W>R W,RBRpi=W>RB,piRS
SSSSSRjRmRR=>m25c,4RmRR=>m256,.RmRR=>m25n,dRmRR=>m25(2C;
M)8Rqev_;-
-

---1-RHDlbCqR)vHRI0#ERHDMoC7Rq71) 1FRVsFRL0sERCRN8NRM8I0sHC-
-RsaNoRC0:HRXDGHM

--DsHLNRs$HCCC;#
kCCRHC#C30D8_FOoH_n44cD3NDk;
#HCRC3CC#_08DHFoOH_#o8MC3DND;H
DLssN$MRkHl#H;#
kCMRkHl#H3FPOlMbFC#M03DND;M
C0$H0Rv)q_R)WHR#
RoRRCsMCH5OR
RRRRRRRRlVNHRD$:0R#soHMRR:="MMFC
";RRRRRRRRI0H8ERR:HCM0oRCs:U=R;RR
RRRRRNRR8I8sHE80RH:RMo0CC:sR=;RURRRRRRRR-L-RHCoRMoFkEFRVsCR8b
0ERRRRRRRR80CbERR:HCM0oRCs:.=R6
n;RRRRRRRR80Fk_osCRL:RFCFDN:MR=NRVD;#CRRRRRR--ERN#Fbk0ks0RCRo
RRRRR8RRHsM_C:oRRFLFDMCNRR:=V#NDCR;RRRRR-E-RN8#RNR0NHkMb0CRsoR
RRRRRR8RN8ss_C:oRRFLFDMCNRR:=V#NDCRRRR-RR-NRE88RN8#sC#CRsoR
RRRRRR;R2
RRRRsbF0
R5RRRRRRRR7amz:kRF00R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj;R
RRRRRRQR7h:RRRRHM#_08DHFoOC_POs0F58IH04E-RI8FMR0Fj
2;RRRRRRRRq)77RH:RM0R#8F_Do_HOP0COFNs58I8sHE80-84RF0IMF2Rj;R
RRRRRR RWRRR:H#MR0D8_FOoH;RRRRRRR-I-RsCH0RNCMLRDCVRFss
NlRRRRRRRRBRpi:MRHR8#0_oDFHRO;RRRRR-R-RFODOV	RFssRNRl,Ns88,HR8MR
RRRRRRBRmp:iRRRHM#_08DHFoORRRRRRR-F-RbO0RD	FORsVFRk8F0R
RRRRRR;R2
8CMR0CMHR0$)_qv)
W;

---w-RH0s#RbHlDCClM00NHRFMl0k#RRLCODNDCN8RsjOE

--NEsOHO0C0CksRFLDOs	_NFlRVqR)vW_)R
H#
lOFbCFMMX0R)4qv.4UX1b
RFRs05R
RR:mRR0FkR8#0_oDFH
O;RqRRjRR:H#MR0D8_FOoH;R
RRRq4:MRHR8#0_oDFH
O;RqRR.RR:H#MR0D8_FOoH;R
RRRqd:MRHR8#0_oDFH
O;RqRRcRR:H#MR0D8_FOoH;R
RRRq6:MRHR8#0_oDFH
O;RqRRnRR:H#MR0D8_FOoH;R
RR:7RRRHM#_08DHFoOR;
RBRWp:iRRRHM#_08DHFoOR;
R RWRH:RM0R#8F_Do
HOR
2;CRM8ObFlFMMC0
;

lOFbCFMMX0R)nqvc1X.
FRbs50R
RRRm:jRR0FkR8#0_oDFH
O;RmRR4RR:FRk0#_08DHFoOR;
RjRqRH:RM0R#8F_Do;HO
RRRq:4RRRHM#_08DHFoOR;
R.RqRH:RM0R#8F_Do;HO
RRRq:dRRRHM#_08DHFoOR;
RcRqRH:RM0R#8F_Do;HO
RRRq:6RRRHM#_08DHFoOR;
RjR7RH:RM0R#8F_Do;HO
RRR7:4RRRHM#_08DHFoOR;
RBRWp:iRRRHM#_08DHFoOR;
R RWRH:RM0R#8F_Do
HOR
2;CRM8ObFlFMMC0
;
ObFlFMMC0)RXq.vdX
c1RsbF0
R5RmRRjRR:FRk0#_08DHFoOR;
R4RmRF:Rk#0R0D8_FOoH;R
RRRm.:kRF00R#8F_Do;HO
RRRm:dRR0FkR8#0_oDFH
O;RqRRjRR:H#MR0D8_FOoH;R
RRRq4:MRHR8#0_oDFH
O;RqRR.RR:H#MR0D8_FOoH;R
RRRqd:MRHR8#0_oDFH
O;RqRRcRR:H#MR0D8_FOoH;R
RRR7j:MRHR8#0_oDFH
O;R7RR4RR:H#MR0D8_FOoH;R
RRR7.:MRHR8#0_oDFH
O;R7RRdRR:H#MR0D8_FOoH;R
RRpWBiRR:H#MR0D8_FOoH;R
RRRW :MRHR8#0_oDFHRO
2C;
MO8RFFlbM0CM;F
OlMbFCRM0Xv)qdU.X1R

b0FsRR5
RRRm:kRF00R#8F_Do_HOP0COF(s5RI8FMR0Fj
2;RqRRjRR:H#MR0D8_FOoH;R
RRRq4:MRHR8#0_oDFH
O;RqRR.RR:H#MR0D8_FOoH;R
RRRqd:MRHR8#0_oDFH
O;RqRRcRR:H#MR0D8_FOoH;R
RR:7RRRHM#_08DHFoOC_POs0F58(RF0IMF2Rj;R
RRpWBiRR:H#MR0D8_FOoH;R
RRRW :MRHR8#0_oDFHRO
2C;
MO8RFFlbM0CM;O

FFlbM0CMRqX)vX4nUR1
b0FsRR5
RRRm:kRF00R#8F_Do_HOP0COF(s5RI8FMR0Fj
2;RqRRjRR:H#MR0D8_FOoH;R
RRRq4:MRHR8#0_oDFH
O;RqRR.RR:H#MR0D8_FOoH;R
RRRqd:MRHR8#0_oDFH
O;R7RRRH:RM0R#8F_Do_HOP0COF(s5RI8FMR0Fj
2;RWRRBRpi:MRHR8#0_oDFH
O;RWRR RR:H#MR0D8_FOoH
;R2
8CMRlOFbCFMM
0;
MVkOF0HMkRVMHO_M5H0LRR:LDFFC2NMR0sCkRsM#H0sMHoR#C
Lo
HMRVRHR25LRC0EMR
RRCRs0Mks52"";R
RCCD#
RRRR0sCk5sM"kBFDM8RFH0RlCbDl0CMRFADO)	RqRv3Q0#REsCRCRN8Ns88CR##sHCo#s0CCk8R#oHMRC0ERl#NCDROFRO	N0#RE)CRq"v?2R;
R8CMR;HV
8CMRMVkOM_HH
0;VOkM0MHFR0oC_8CM_b8C0#E5HRxC:MRH0CCosRR;80CbERR:HCM0o2CsR0sCkRsMHCM0oRCsHP#
NNsHLRDCl_HM#CHxRH:RMo0CC:sR=;Rj
oLCHRM
RMlH_x#HC=R:Rb8C0
E;RVRHRH5#x<CRRb8C0RE20MEC
RRRRMlH_x#HC=R:Rx#HCR;
R8CMR;HV
sRRCs0kMHRlMH_#x
C;CRM8o_C0C_M880CbEN;
0H0sLCk0RMoCC0sNFss_CsbF0RR:#H0sM
o;Ns00H0LkCCRoMNCs0_FssFCbsF0RVDRLF_O	sRNl:sRNO0EHCkO0sHCR#kRVMHO_M5H0Ns88_osC2-;
-CRLoRHMLODF	NRsllRHblDCCNM00MHFRo#HM#ND
b0$CMRH0s_NsRN$HN#Rs$sNRR5j06FR2VRFR0HMCsoC;F
OMN#0MI0RHE80_sNsN:$RR0HM_sNsN:$R=4R5,,R.RRc,g4,RUd,Rn
2;O#FM00NMRb8C0NE_s$sNRH:RMN0_s$sNRR:=5d4nURc,U.4g,jRcgRn,.Ujc,jR4.Rc,624.;F
OMN#0M80RH.PdRH:RMo0CC:sR=IR5HE80-/42d
n;O#FM00NMRP8H4:nRR0HMCsoCRR:=58IH04E-2U/4;F
OMN#0M80RHRPU:MRH0CCos=R:RH5I8-0E4g2/;F
OMN#0M80RHRPc:MRH0CCos=R:RH5I8-0E4c2/;F
OMN#0M80RHRP.:MRH0CCos=R:RH5I8-0E4.2/;F
OMN#0M80RHRP4:MRH0CCos=R:RH5I8-0E442/;O

F0M#NRM0LDFF4RR:LDFFCRNM:5=R84HPRj>R2O;
F0M#NRM0LDFF.RR:LDFFCRNM:5=R8.HPRj>R2O;
F0M#NRM0LDFFcRR:LDFFCRNM:5=R8cHPRj>R2O;
F0M#NRM0LDFFURR:LDFFCRNM:5=R8UHPRj>R2O;
F0M#NRM0LDFF4:nRRFLFDMCNRR:=5P8H4>nRR;j2
MOF#M0N0FRLF.DdRL:RFCFDN:MR=8R5H.PdRj>R2
;
O#FM00NMRP8H4UndcRR:HCM0oRCs:5=R80CbE2-4/d4nU
c;O#FM00NMRP8HU.4gRH:RMo0CC:sR=8R5CEb0-/42U.4g;F
OMN#0M80RHjPcg:nRR0HMCsoCRR:=5b8C04E-2j/cg
n;O#FM00NMRP8H.UjcRH:RMo0CC:sR=8R5CEb0-/42.Ujc;F
OMN#0M80RHjP4.:cRR0HMCsoCRR:=5b8C04E-2j/4.
c;O#FM00NMRP8H6R4.:MRH0CCos=R:RC58b-0E462/4
.;
MOF#M0N0FRLF4D6.RR:LDFFCRNM:5=R86HP4>.RR;j2
MOF#M0N0FRLFjD4.:cRRFLFDMCNRR:=5P8H4cj.Rj>R2O;
F0M#NRM0LDFF.UjcRL:RFCFDN:MR=8R5HjP.c>URR;j2
MOF#M0N0FRLFjDcg:nRRFLFDMCNRR:=5P8HcnjgRj>R2O;
F0M#NRM0LDFFU.4gRL:RFCFDN:MR=8R5H4PUg>.RR;j2
MOF#M0N0FRLFnD4dRUc:FRLFNDCM=R:RH58Pd4nU>cRR;j2
F
OMN#0M#0RkIl_HE80RH:RMo0CC:sR=mRAmqp hF'b#F5LF2D4RA+Rm mpqbh'FL#5F.FD2RR+Apmm 'qhb5F#LDFFc+2RRmAmph q'#bF5FLFDRU2+mRAmqp hF'b#F5LFnD42O;
F0M#NRM0#_kl80CbERR:HCM0oRCs:6=RR5-RApmm 'qhb5F#LDFF624.RA+Rm mpqbh'FL#5F4FDj2.cRA+Rm mpqbh'FL#5F.FDj2cURA+Rm mpqbh'FL#5FcFDj2gnRA+Rm mpqbh'FL#5FUFD42g.2
;
O#FM00NMROI_EOFHCH_I8R0E:MRH0CCos=R:R8IH0NE_s$sN5l#k_8IH0;E2
MOF#M0N0_RIOHEFO8C_CEb0RH:RMo0CC:sR=CR8b_0ENNss$k5#lH_I820E;F
OMN#0M80R_FOEH_OCI0H8ERR:HCM0oRCs:I=RHE80_sNsN#$5k8l_CEb02O;
F0M#NRM08E_OFCHO_b8C0:ERR0HMCsoCRR:=80CbEs_Ns5N$#_kl80CbE
2;
MOF#M0N0_RII0H8Ek_MlC_ODRD#:MRH0CCos=R:RH5I8-0E4I2/_FOEH_OCI0H8ERR+4O;
F0M#NRM0IC_8b_0EM_klODCD#RR:HCM0oRCs:5=R80CbE2-4/OI_EOFHCC_8bR0E+;R4
F
OMN#0M80R_8IH0ME_kOl_C#DDRH:RMo0CC:sR=IR5HE80-/428E_OFCHO_8IH0+ERR
4;O#FM00NMR88_CEb0_lMk_DOCD:#RR0HMCsoCRR:=5b8C04E-2_/8OHEFO8C_CEb0R4+R;O

F0M#NRM0IH_#x:CRR0HMCsoCRR:=IH_I8_0EM_klODCD#RR*IC_8b_0EM_klODCD#O;
F0M#NRM08H_#x:CRR0HMCsoCRR:=8H_I8_0EM_klODCD#RR*8C_8b_0EM_klODCD#
;
O#FM00NMRFLFDR_8:FRLFNDCM=R:R_58#CHxRI-R_x#HC=R<R;j2
MOF#M0N0FRLFID_RL:RFCFDN:MR=FRM0F5LF8D_2
;
O#FM00NMRFOEH_OCI0H8ERR:HCM0oRCs:5=RApmm 'qhb5F#LDFF_R82*_R8OHEFOIC_HE802RR+5mAmph q'#bF5FLFD2_IRI*R_FOEH_OCI0H8E
2;O#FM00NMRFOEH_OC80CbERR:HCM0oRCs:5=RApmm 'qhb5F#LDFF_R82*_R8OHEFO8C_CEb02RR+5mAmph q'#bF5FLFD2_IRI*R_FOEH_OC80CbE
2;O#FM00NMR8IH0ME_kOl_C#DDRH:RMo0CC:sR=AR5m mpqbh'FL#5F_FD8*2R58IH04E-2_/8OHEFOIC_HE802RR+5mAmph q'#bF5FLFD2_IR5*RI0H8E2-4/OI_EOFHCH_I820ER4+R;F
OMN#0M80RCEb0_lMk_DOCD:#RR0HMCsoCRR:=5mAmph q'#bF5FLFD2_8R8*5CEb0-/428E_OFCHO_b8C0RE2+AR5m mpqbh'FL#5F_FDI*2RRC58b-0E4I2/_FOEH_OC80CbE+2RR
4;-F-OMN#0MM0RkOl_C#DDRH:RMo0CC:sR=5R55b8C0-ERRR42/.Rd2RR+5855CEb0R4-R2FRl8.Rd2RR/42n2;RRR-y-RRRFV)dqv.1X4RDOCDM#RCCC88-R
-MOF#M0N0CRDVF0_PRCs:MRH0CCos=R:R55580CbERR+4R62lRF8dR.2/nR42R;RRRRRRRRRRRRRRRRRRRRRR-RR-RRyF)VRqnv4XR41M8CCCV8RFDsRCRV0FsPCRsIF80#
$RbCF_k0L4k#_b0$C#RHRsNsN5$R80CbEk_MlC_OD-D#4FR8IFM0RRj,I0H8Ek_MlC_OD-D#4FR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNR0Fk_#Lk4RR:F_k0L4k#_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFR8s_FRk05bHMk00RFsR0H0-#N#0C2$
0bFCRkL0_k_#.0C$bRRH#NNss$8R5CEb0_lMk_DOCD4#-RI8FMR0Fj.,R*8IH0ME_kOl_C#DD+84RF0IMF2RjRRFV#_08DHFoO#;
HNoMDkRF0k_L#:.RR0Fk_#Lk.$_0bRC;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RV_Rs80FkRM5HbRk000FRs#H-0CN0#02
$RbCF_k0Lck#_b0$C#RHRsNsN5$R80CbEk_MlC_OD-D#4FR8IFM0RRj,cH*I8_0EM_klODCD#R+d8MFI0jFR2VRFR8#0_oDFH
O;#MHoNFDRkL0_kR#c:kRF0k_L#0c_$;bCRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$FsVR_k8F0HR5M0bkRR0F0-sH#00NC
#20C$bR0Fk_#LkU$_0bHCR#sRNsRN$5b8C0ME_kOl_C#DD-84RF0IMF,RjRIU*HE80_lMk_DOCD(#+RI8FMR0FjF2RV0R#8F_Do;HO
o#HMRNDF_k0LUk#RF:RkL0_k_#U0C$b;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFVsF_8k50RHkMb0FR0RH0s-N#002C#
b0$CNRbs$H0_#LkU$_0bHCR#sRNsRN$5b8C0ME_kOl_C#DD-84RF0IMF,RjR8IH0ME_kOl_C#DD-84RF0IMF2RjRRFV#_08DHFoO#;
HNoMDNRbs$H0_#LkURR:bHNs0L$_k_#U0C$b;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RV_Rs80FkRM5HbRk000FRs#H-0CN0#02
$RbCF_k0L4k#n$_0bHCR#sRNsRN$5b8C0ME_kOl_C#DD-84RF0IMF,RjR*4nI0H8Ek_MlC_OD+D#486RF0IMF2RjRRFV#_08DHFoO#;
HNoMDkRF0k_L#R4n:kRF0k_L#_4n0C$b;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFVsF_8k50RHkMb0FR0RH0s-N#002C#
b0$CNRbs$H0_#Lk40n_$RbCHN#Rs$sNRC58b_0EM_klODCD#R-48MFI0jFR,*R.I0H8Ek_MlC_OD+D#4FR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNRsbNH_0$L4k#nRR:bHNs0L$_kn#4_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$FsVR_k8F0HR5M0bkRR0F0-sH#00NC
#20C$bR0Fk_#Lkd0._$RbCHN#Rs$sNRC58b_0EM_klODCD#R-48MFI0jFR,.Rd*8IH0ME_kOl_C#DD+Rd48MFI0jFR2VRFR8#0_oDFH
O;#MHoNFDRkL0_k.#dRF:RkL0_k.#d_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFR8s_FRk05bHMk00RFsR0H0-#N#0C2$
0bbCRN0sH$k_L#_d.0C$bRRH#NNss$8R5CEb0_lMk_DOCD4#-RI8FMR0Fjc,R*8IH0ME_kOl_C#DD+8dRF0IMF2RjRRFV#_08DHFoO#;
HNoMDNRbs$H0_#Lkd:.RRsbNH_0$Ldk#.$_0bRC;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFVsF_8k50RHkMb0FR0RH0s-N#002C#
o#HMRNDF_k0C:MRR8#0_oDFHPO_CFO0sC58b_0EM_klODCD#R-48MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-MRCNCLD#FRVssR0H0-#N#0C
o#HMRNDI_s0C:MRR8#0_oDFHPO_CFO0sC58b_0EM_klODCD#R-48MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-sRIHR0CCLMNDRC#VRFsCENORIsFRRFV)RqvODCD#H
#oDMNR_HMsRCo:0R#8F_Do_HOP0COFIs5HE80+Rd68MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--k8#CRR0FsHCo#s0CRh7QRH
#oDMNR0Fk_osCR#:R0D8_FOoH_OPC05FsI0H8E6+dRI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--k8#CRR0FsHCo#s0CRz7maH
#oDMNR0Fk_osC4RR:#_08DHFoOC_POs0F58IH04E-RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-k-R#RC80OFRE#FFCCRL0CICMQR7hMRN8kRF00bkRRFVAODF	qR)vH
#oDMNR_N8sRCo:0R#8F_Do_HOP0COFNs58I8sHE80-84RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-k-R#RC80sFRC#oH0RCsq)77RsVFRHIs0#C
HNoMDFRDIN_s8R8s:0R#8F_Do_HOP0COF4s5dFR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-NRs8R8sL#H0RbHMk00RFqR)vCRODRD#5LcRHR0#skCJH8sC2H
#oDMNRIDF_8IN8:sRR8#0_oDFHPO_CFO0sd54RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-R8IN8LsRHR0#HkMb0FR0Rv)qRDOCD5#RcHRL0s#RCHJks2C8
o#HMRND)7q7)l_0bRR:#_08DHFoOC_POs0F58N8s8IH04E-RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RCk#8FR0RbbHCMDHCqR)7
7)#MHoNWDRq)77_b0lR#:R0D8_FOoH_OPC05FsNs88I0H8ER-48MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--k8#CRR0FbCHbDCHMR7Wq7#)
HNoMDQR7hl_0bRR:#_08DHFoOC_POs0F58IH04E-RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-k-R#RC80bFRHDbCHRMC7
Qh#MHoNWDR l_0bRR:#_08DHFoOR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RCk#8FR0RbbHCMDHC RW
R--CRM8LODF	NRsllRHblDCCNM00MHFRo#HM#ND
-
-RoLCH#MRCODC0NRsllRHblDCCNM00MHFRo#HM#ND
b0$CCRDVP0FC0s_RRH#NNss$jR5RR0FdF2RVMRH0CCos0;
$RbCD0CVFsPC_.0_RRH#NNss$jR5RR0F4F2RVMRH0CCosV;
k0MOHRFMb5N8HRR:#_08DHFoOC_POs0F;4RI,.RIRH:RMo0CCRs2skC0s#MR0D8_FOoH_OPC0RFsHP#
NNsHLRDCPRNs:0R#8F_Do_HOP0COFIs54R-48MFI0jFR2L;
CMoH
VRRF[sRRRHMP'NssoNMCFRDFRb
RHRRV[R5RR<=IR.20MECRR
SRsPN5R[2:H=R5DH'F[I+2S;
CCD#
RSRP5Ns[:2R=jR''S;
CRM8H
V;RMRC8FRDF
b;RCRs0MksRsPN;M
C8NRb8V;
k0MOHRFMo_C0I0H8E5_UI0H8EH:RMo0CCRs2skC0sHMRMo0CCHsR#N
PsLHNDPCRN:DRR0HMCsoCRR:=jL;
CMoH
PRRN:DR=HRI8/0EUR;
RRHV5H5I8R0ElRF8U>2RRRc20MEC
RRRRDPNRR:=PRND+;R4
CRRMH8RVR;
R0sCkRsMP;ND
8CMR0oC_8IH0UE_;k
VMHO0FoMRCI0_HE80_I.5HE80:MRH0CCoss2RCs0kMMRH0CCos#RH
sPNHDNLCNRPDRR:HCM0oRCs:j=R;C
Lo
HMRNRPD=R:R8IH0.E/;R
RskC0sPMRN
D;CRM8o_C0I0H8E;_.
MVkOF0HMCRo0H_I850EI0H8ERR:HCM0o2CsR0sCkRsMD0CVFsPC_.0_R
H#PHNsNCLDRDPNRD:RCFV0P_Cs0;_.
oLCHRM
RDPN5R42:o=RCI0_HE80_I.5HE802R;
RRHV58IH0lERF.8RRj=R2ER0CRM
RPRRNjD52=R:R
j;RDRC#RC
RPRRNjD52=R:R
4;RMRC8VRH;R
RskC0sPMRN
D;CRM8o_C0I0H8EV;
k0MOHRFMo_C0I0H8EH5I8R0E:MRH0CCoss2RCs0kMCRDVP0FC0s_R
H#PHNsNCLDRDPNRD:RCFV0P_Cs0=R:R,5jRRj,jj,R2L;
CMoH
PRRNdD52=R:R0oC_8IH0UE_58IH0;E2
ORRNR#C58IH0lERFU8R2#RH
IRRERCMcRR|d>R=RDPN5R.2:4=R;R
RIMECR=.R>NRPD254RR:=4R;
RCIEMRR4=P>RNjD52=R:R
4;RERICFMR0sEC#>R=RDMkDR;
R8CMR#ONCR;
R0sCkRsMP;ND
8CMR0oC_8IH0
E;O#FM00NMRI#_HE80_sNsN:$RRVDC0CFPsR_0:o=RCI0_HE8058IH0;E2
MOF#M0N0_R#I0H8Es_Ns_N$n:cRRVDC0CFPs__0.=R:R0oC_8IH0IE5HE802V;
k0MOHRFMo_C0M_kl45.U80CbEH:RMo0CCRs2skC0sHMRMo0CCHsR#N
PsLHNDPCRN:DRR0HMCsoCRR:=jL;
CMoH
PRRN:DR=CR8b/0E4;.U
HRRV5R580CbEFRl8.R4U>2RR.442ER0CRM
RPRRN:DR=NRPDRR+4R;
R8CMR;HV
sRRCs0kMNRPDC;
Mo8RCM0_k4l_.
U;VOkM0MHFR0oC_VDC0CFPsc_n5b8C0:ERR0HMCsoC2CRs0MksR0HMCsoCR
H#LHCoMR
RskC0s8M5CEb0R8lFRU4.2C;
Mo8RCD0_CFV0P_Csn
c;VOkM0MHFR0oC_lMk_5nc80CbERR:HCM0o2CsR0sCkRsMHCM0oRCsHP#
NNsHLRDCPRND:MRH0CCos=R:R
j;LHCoMR
RRRHV5b8C0<ER=4R4.MRN8CR8bR0E>URc2ER0CRM
RRRRPRND:4=R;R
RCRM8H
V;RCRs0MksRDPN;M
C8CRo0k_Mlc_n;k
VMHO0FoMRCD0_CFV0P5Cs80CbERR:HCM0o;CsRGlNRH:RMo0CCRs2skC0sHMRMo0CCHsR#N
PsLHNDPCRN:DRR0HMCsoCRR:=jL;
CMoH
HRRV8R5CEb0Rl-RN>GR=2RjRC0EMR
RRNRPD=R:Rb8C0-ERRGlN;R
RCCD#
RRRRDPNRR:=80CbER;
R8CMR;HV
sRRCs0kMN5PD
2;CRM8o_C0D0CVFsPC;k
VMHO0FoMRCM0_kdl_.C58bR0E:MRH0CCoss2RCs0kMMRH0CCos#RH
sPNHDNLCNRPDRR:HCM0oRCs:j=R;C
Lo
HMRVRHRC58bR0E<c=RUMRN8CR8bR0E>nR42ER0CRM
RRRRPRND:4=R;R
RCRM8H
V;RCRs0MksRDPN;M
C8CRo0k_Ml._d;k
VMHO0FoMRCM0_k4l_nC58bR0E:MRH0CCoss2RCs0kMMRH0CCos#RH
sPNHDNLCNRPDRR:HCM0oRCs:j=R;C
Lo
HMRVRHRC58bR0E<4=RnMRN8CR8bR0E>2RjRC0EMR
RRPRRN:DR=;R4
CRRMH8RVR;
R0sCkRsMP;ND
8CMR0oC_lMk_;4n
O--F0M#NRM0M_klODCD#RR:HCM0oRCs:5=R5C58bR0E-2R4Rd/R.+2RR55580CbERR-4l2RFd8R./2RR24n2R;RRR--yVRFRv)qd4.X1CRODRD#M8CCC
8RO#FM00NMRlMk_DOCD._4URR:HCM0oRCs:o=RCM0_k4l_.8U5CEb02O;
F0M#NRM0D0CVFsPC_Rnc:MRH0CCos=R:R0oC_VDC0CFPsc_n5b8C0;E2
MOF#M0N0kRMlC_ODnD_cRR:HCM0oRCs:o=RCM0_knl_cC5DVP0FCns_c
2;O#FM00NMRVDC0CFPs._dRH:RMo0CC:sR=CRo0C_DVP0FCDs5CFV0P_CsnRc,n;c2
MOF#M0N0kRMlC_ODdD_.RR:HCM0oRCs:o=RCM0_kdl_.C5DVP0FCds_.
2;O#FM00NMRVDC0CFPsn_4RH:RMo0CC:sR=CRo0C_DVP0FCDs5CFV0P_CsdR.,d;.2
MOF#M0N0kRMlC_OD4D_nRR:HCM0oRCs:o=RCM0_k4l_nC5DVP0FC4s_n
2;
b0$CkRF0k_L#$_0b4C_.HUR#sRNsRN$5lMk_DOCD._4UFR8IFM0RRj,I0H8ER-48MFI0jFR2VRFR8#0_oDFH
O;0C$bR0Fk_#Lk_b0$Cc_nRRH#NNss$MR5kOl_C_DDn8cRF0IMF,RjR8IH04E-RI8FMR0FjF2RV0R#8F_Do;HO
b0$CkRF0k_L#$_0bdC_.#RHRsNsN5$RM_klODCD_Rd.8MFI0jFR,HRI8-0E4FR8IFM0RRj2F#VR0D8_FOoH;$
0bFCRkL0_k0#_$_bC4HnR#sRNsRN$5lMk_DOCDn_4RI8FMR0FjI,RHE80-84RF0IMF2RjRRFV#_08DHFoO#;
HNoMDkRF0k_L#._4URR:F_k0L_k#0C$b_U4.;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFV80FkRM5HbRk000FRs#H-0CN0##2
HNoMDkRF0k_L#c_nRF:RkL0_k0#_$_bCnRc;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RVFR8k50RHkMb0FR0RH0s-N#002C#
o#HMRNDF_k0L_k#d:.RR0Fk_#Lk_b0$C._d;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFV80FkRM5HbRk000FRs#H-0CN0##2
HNoMDkRF0k_L#n_4RF:RkL0_k0#_$_bC4Rn;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RVFR8k50RHkMb0FR0RH0s-N#002C#
o#HMRND#k_F0M_CR#:R0D8_FOoH_OPC05FsM_klODCD_U4.RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-C-RMDNLCV#RF0sRs#H-0CN0#H
#oDMNR0Fk__CMn:cRR8#0_oDFH
O;#MHoNFDRkC0_M._dR#:R0D8_FOoH;H
#oDMNR0Fk__CM4:nRR8#0_oDFH
O;#MHoN#DR_0Is_RCM:0R#8F_Do_HOP0COFMs5kOl_C_DD4R.U8MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-sRIHR0CCLMNDRC#VRFsCENORIsFRRFV)RqvODCD#H
#oDMNR0Is__CMn:cRR8#0_oDFH
O;#MHoNIDRsC0_M._dR#:R0D8_FOoH;H
#oDMNR0Is__CM4:nRR8#0_oDFH
O;#MHoN#DR__HMsRCo:0R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-k-R#RC80sFRC#oH0RCs7RQh
o#HMRND#k_F0C_soRR:#_08DHFoOC_POs0F58IH04E-RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--k8#CRR0FsHCo#s0CRz7maH
#oDMNRN#_8C_soRR:#_08DHFoOC_POs0F58N8s8IH04E-RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RCk#8FR0RosCHC#0s7Rq7#)
HNoMDFRDI8_N8:sRR8#0_oDFHPO_CFO0sR5n8MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--Ns88R0LH#MRHbRk00)FRqOvRC#DDRR5cL#H0RJsCkCHs8O2
F0M#NRM0D_#LI0H8ERR:HCM0oRCs:I=RHE80-5U*#H_I8_0ENNss$25d--42c_*#I0H8Es_Ns5N$..2-*I#_HE80_sNsN4$52_-#I0H8Es_Ns5N$j
2;0C$bRb0l_sNsNR$UHN#Rs$sNR_5#I0H8Es_Ns5N$d42-RI8FMR0FjF2RV0R#8F_Do_HOP0COF(s5RI8FMR0Fj
2;#MHoN0DRlUb__,d.Rb0l_4U_nRR:0_lbNNss$
U;-C-RM#8RCODC0NRsllRHblDCCNM00MHFRo#HM#ND
0N0skHL0\CR3lsN_VFV#\C0R#:R0MsHo
;
LHCoMR
R
zRRc:dRRRHV58N8sC_soo2RCsMCNR0C-o-RCsMCNR0CLODF	NRslR
RR-R-RRQVNs88I0H8ERR<OHEFOIC_HE80R#N#HRoM'Rj'0kFRMCk#8HRL0R#
RzRRj:RRRRHV58N8s8IH0=ERRR42oCCMsCN0
RRRRRRRRIDF_8sN8<sR=jR"jjjjjjjjjjjj"RR&q)775;j2
RRRRRRRRIDF_8IN8<sR=jR"jjjjjjjjjjjj"RR&Ns8_Cjo52R;
RCRRMo8RCsMCNR0Cz
j;RRRRzR4R:VRHR85N8HsI8R0E=2R.RMoCC0sNCR
RRRRRRFRDIN_s8R8s<"=Rjjjjjjjjjjjj"RR&q)77584RF0IMF2Rj;R
RRRRRRFRDIN_I8R8s<"=Rjjjjjjjjjjjj"RR&Ns8_C4o5RI8FMR0Fj
2;RRRRCRM8oCCMsCN0R;z4
RRRRRz.RH:RVNR58I8sHE80Rd=R2CRoMNCs0RC
RRRRRDRRFsI_Ns88RR<="jjjjjjjjjjj"RR&q)7758.RF0IMF2Rj;R
RRRRRRFRDIN_I8R8s<"=Rjjjjjjjjj"jjRN&R8C_soR5.8MFI0jFR2R;
RCRRMo8RCsMCNR0Cz
.;RRRRzRdR:VRHR85N8HsI8R0E=2RcRMoCC0sNCR
RRRRRRFRDIN_s8R8s<"=RjjjjjjjjjRj"&7Rq7d)5RI8FMR0Fj
2;RRRRRRRRD_FII8N8s=R<Rj"jjjjjjjjj"RR&Ns8_Cdo5RI8FMR0Fj
2;RRRRCRM8oCCMsCN0R;zd
RRRRRzcRH:RVNR58I8sHE80R6=R2CRoMNCs0RC
RRRRRDRRFsI_Ns88RR<="jjjjjjjjRj"&7Rq7c)5RI8FMR0Fj
2;RRRRRRRRD_FII8N8s=R<Rj"jjjjjj"jjRN&R8C_soR5c8MFI0jFR2R;
RCRRMo8RCsMCNR0Cz
c;RRRRzR6R:VRHR85N8HsI8R0E=2RnRMoCC0sNCR
RRRRRRFRDIN_s8R8s<"=Rjjjjjjjj"RR&q)77586RF0IMF2Rj;R
RRRRRRFRDIN_I8R8s<"=Rjjjjjjjj"RR&Ns8_C6o5RI8FMR0Fj
2;RRRRCRM8oCCMsCN0R;z6
RRRRRznRH:RVNR58I8sHE80R(=R2CRoMNCs0RC
RRRRRDRRFsI_Ns88RR<="jjjjjjj"RR&q)7758nRF0IMF2Rj;R
RRRRRRFRDIN_I8R8s<"=Rjjjjj"jjRN&R8C_soR5n8MFI0jFR2R;
RCRRMo8RCsMCNR0Cz
n;RRRRzR(R:VRHR85N8HsI8R0E=2RURMoCC0sNCR
RRRRRRFRDIN_s8R8s<"=RjjjjjRj"&7Rq7()5RI8FMR0Fj
2;RRRRRRRRD_FII8N8s=R<Rj"jjjjj"RR&Ns8_C(o5RI8FMR0Fj
2;RRRRCRM8oCCMsCN0R;z(
RRRRRzURH:RVNR58I8sHE80Rg=R2CRoMNCs0RC
RRRRRDRRFsI_Ns88RR<="jjjjRj"&7Rq7U)5RI8FMR0Fj
2;RRRRRRRRD_FII8N8s=R<Rj"jj"jjRN&R8C_soR5U8MFI0jFR2R;
RCRRMo8RCsMCNR0Cz
U;RRRRzRgR:VRHR85N8HsI8R0E=jR42CRoMNCs0RC
RRRRRDRRFsI_Ns88RR<="jjjj&"RR7q7)R5g8MFI0jFR2R;
RRRRRDRRFII_Ns88RR<="jjjj&"RR_N8s5CogFR8IFM0R;j2
RRRR8CMRMoCC0sNCgRz;R
RR4Rzj:RRRRHV58N8s8IH0=ERR244RMoCC0sNCR
RRRRRRFRDIN_s8R8s<"=Rj"jjRq&R757)48jRF0IMF2Rj;R
RRRRRRFRDIN_I8R8s<"=Rj"jjRN&R8C_soj54RI8FMR0Fj
2;RRRRCRM8oCCMsCN0Rjz4;R
RR4Rz4:RRRRHV58N8s8IH0=ERR24.RMoCC0sNCR
RRRRRRFRDIN_s8R8s<"=RjRj"&7Rq74)54FR8IFM0R;j2
RRRRRRRRIDF_8IN8<sR=jR"j&"RR_N8s5Co484RF0IMF2Rj;R
RRMRC8CRoMNCs0zCR4
4;RRRRzR4.RH:RVNR58I8sHE80R4=Rdo2RCsMCN
0CRRRRRRRRD_FIs8N8s=R<R''jRq&R757)48.RF0IMF2Rj;R
RRRRRRFRDIN_I8R8s<'=Rj&'RR_N8s5Co48.RF0IMF2Rj;R
RRMRC8CRoMNCs0zCR4
.;RRRRzR4dRH:RVNR58I8sHE80R4>Rdo2RCsMCN
0CRRRRRRRRD_FIs8N8s=R<R7q7)d54RI8FMR0Fj
2;RRRRRRRRD_FII8N8s=R<R_N8s5Co48dRF0IMF2Rj;R
RRMRC8CRoMNCs0zCR4
d;
RRRRR--Q5VR8_HMs2CoRosCHC#0sQR7h#RkHRMoB
piRRRRzR4cRH:RV8R5HsM_CRo2oCCMsCN0
RRRRRRRRFbsO#C#Rp5Bi7,RQRh2LHCoMR
RRRRRRRRRRVRHRp5BiRR='R4'NRM8B'piCMPC002RE
CMRRRRRRRRRRRRRRRRHsM_C<oR="R5jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"RR&72Qh;R
RRRRRRRRRRMRC8VRH;R
RRRRRRMRC8sRbF#OC#R;
RCRRMo8RCsMCNR0Cz;4c
RRRR6z4RRR:H5VRMRF08_HMs2CoRMoCC0sNCR
RRRRRRRRRRMRH_osCRR<=5j"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjRj"&QR7h
2;RRRRCRM8oCCMsCN0R6z4;R

R-RR-VRQR85sF_k0s2CoRosCHC#0s_R)7amzRHk#M)oR_pmBiR
RR4Rzn:RRRRHV5k8F0C_soo2RCsMCN
0CRRRRRRRRbOsFCR##5pmBiF,Rks0_C2o4RoLCHRM
RRRRRRRRRHRRVmR5BRpi=4R''MRN8BRmpCi'P0CM2ER0CRM
RRRRRRRRRRRRR7RRmRza<F=Rks0_C;o4
RRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMRFbsO#C#;R
RRRRRRMRC8CRoMNCs0zCR4
n;RRRRzR4(RH:RVMR5F80RF_k0s2CoRMoCC0sNCR
RRRRRRRRRRmR7z<aR=kRF0C_so
4;RRRRCRM8oCCMsCN0R(z4;R

R-RR-VRQR85N8ss_CRo2sHCo#s0CR7q7)FRVssRIHR0CkM#HopRBiR
RR4RzURIR:VRHR85N8ss_CRo2oCCMsCN0
RRRRRRRRFbsO#C#Rp5Biq,R727)RoLCHRM
RRRRRRRRRHRRVBR5p=iRR''4R8NMRiBp'CCPMR020MEC
RRRRRRRRRRRRRRRR_N8sRCo<q=R757)Ns88I0H8ER-48MFI0jFR2R;
RRRRRRRRRCRRMH8RVR;
RRRRRCRRMb8RsCFO#
#;RRRRCRM8oCCMsCN0RUz4IR;
RzRR4RgI:VRHRF5M08RN8ss_CRo2oCCMsCN0
RRRRRRRRRRRR_N8sRCo<q=R7;7)
RRRR8CMRMoCC0sNC4Rzg
I;
RRRRR-- sG0NFRDoRHOVRFs7DkNRsbF0NRO#RC
RzRRsRCo:sRbF#OC#p5BiL2RCMoH
RRRRHRRVBR5p i'ea hR8NMRiBpR'=R4R'20MEC
RRRRRRR7_Qh0Rlb<7=RQ
h;RRRRR)RRq)77_b0lRR<=q)77;R
RRRRRR7Wq70)_l<bR=8RN_osC;R
RRRRRR_W 0Rlb<W=R R;
RRRRR8CMR;HV
RRRR8CMRFbsO#C#;R

R-RR-VRQRN)C88Rq8#sC#RR=W0sHC8Rq8#sC#L,R$#bN#QR7hFR0R0FkbRk0HWVR #RHRNCML8DC
RRRRkzlGRR:bOsFC5##W0 _lRb,)7q7)l_0bW,Rq)77_b0l,QR7hl_0bF,Rks0_C
o2RRRRRCRLo
HMRRRRRRRRH5VRW7q7)l_0bRR=)7q7)l_0bMRN8 RW_b0lR'=R4R'20MEC
RRRRRRRRFRRks0_CRo4<7=RQ0h_l
b;RRRRRRRRCCD#
RRRRRRRRFRRks0_CRo4<F=Rks0_CIo5HE80-84RF0IMF2Rj;R
RRRRRRMRC8VRH;R
RRMRC8sRbF#OC#R;
RRRRR
RRRRRR-t-RCsMCNR0C0REC)RqvODCD#MRN8CR#D0CORoDFHVORF)sRq4vAn4_1_
14RRRRzR4U:VRHRE5OFCHO_8IH0=ERRR42oCCMsCN0
RRRRRRRRgz4RV:RFHsRRRHM5b8C0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CRRRR-Q-RVNR58I8sHE80R4>RcM2RCRC80OFRs0CNCsRIHR0CCLMNDNCRMF8Rkk0b0MRCNCLDRD#CCRO0DHFoOR
RRRRRRRRRR.RzjRR:H5VRNs88I0H8ERR>4Rc2oCCMsCN0
RRRRRRRRRRRRRRRR0Fk_5CMH<2R=4R''ERIC5MR)7q7)l_0b85N8HsI8-0E4FR8IFM0R24cRH=R2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0CHM52=R<RRW IMECR85N_osC58N8s8IH04E-RI8FMR0F4Rc2=2RHR#CDCjR''R;
RRRRRRRRRCRRMo8RCsMCNR0Cz;.j
RRRRR--Q5VRNs88I0H8E=R<R24.RRMFI0sHCMRCNCLDRRFsFbk0kC0RMDNLCCR#D0CORoDFHMORCCC88R
RRRRRRRRRR.Rz4RR:H5VRNs88I0H8E=R<R24cRMoCC0sNCR
RRRRRRRRRRRRRRkRF0M_C5RH2<'=R4
';RRRRRRRRRRRRRRRRI_s0CHM52=R<R;W 
RRRRRRRRRRRR8CMRMoCC0sNC.Rz4R;
R-RR-CRtMNCs00CRE)CRqOvRC#DDR8NMRH0s-N#00
C#RRRRRRRRRRRRzR..:FRVsRR[H5MRI0H8Ek_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0RC
RRRRRRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)RAq4v_ncdUXR47:NRDLRCDH"#RW
";RRRRRRRRRRRRRRRRLHCoMR
RRRRRRRRRRRRRR)RAq4v_ncdUXR47:qR)vnA4__141R4
RRRRRRRRRRRRRbRRFRs0lRNb5q7Q5Rj2=H>RMC_so25[,7Rq7R)q=D>RFII_Ns885R4d8MFI0jFR27,RQ=AR>jR""q,R7A7)RR=>D_FIs8N8sd54RI8FMR0Fj
2,RRRRRRRRRRRRRRRR Rhq='>R4R',1q1)RR=>',j'RqW RR=>I_s0CHM52B,RpRiq=B>RpRi, RhA='>R4R',1A1)RR=>',j'RAW RR=>',j'RiBpA>R=RiBp,R
RRRRRRRRRRRRRRmR7q>R=RCFbM7,RmjA52>R=R0Fk_#Lk4,5H[;22
R
RRRRRRRRRRRRRRkRF0C_so25[RR<=F_k0L4k#5[H,2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRCRRMo8RCsMCNR0Cz;..
RRRRRRRR8CMRMoCC0sNC4RzgR;
RCRRMo8RCsMCNR0Cz;4URRRR
RRRR
RRRRRR-t-RCsMCNR0C0REC)RqvODCD#MRN8CR#D0CORoDFHVORF)sRq4vAn._1_
1.RRRRzR.d:VRHRE5OFCHO_8IH0=ERRR.2oCCMsCN0
RRRRRRRRcz.RV:RFHsRRRHM5b8C0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CRRRR-Q-RVNR58I8sHE80R4>RdM2RCRC80OFRs0CNCsRIHR0CCLMNDNCRMF8Rkk0b0MRCNCLDRD#CCRO0DHFoOR
RRRRRRRRRR.Rz6RR:H5VRNs88I0H8ERR>4Rd2oCCMsCN0
RRRRRRRRRRRRRRRR0Fk_5CMH<2R=4R''ERIC5MR)7q7)l_0b85N8HsI8-0E4FR8IFM0R24dRH=R2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0CHM52=R<RRW IMECR85N_osC58N8s8IH04E-RI8FMR0F4Rd2=2RHR#CDCjR''R;
RRRRRRRRRCRRMo8RCsMCNR0Cz;.6
RRRRR--Q5VRNs88I0H8E=R<R24dRRMFI0sHCMRCNCLDRRFsFbk0kC0RMDNLCCR#D0CORoDFHMORCCC88R
RRRRRRRRRR.RznRR:H5VRNs88I0H8E=R<R24dRMoCC0sNCR
RRRRRRRRRRRRRRkRF0M_C5RH2<'=R4
';RRRRRRRRRRRRRRRRI_s0CHM52=R<R;W 
RRRRRRRRRRRR8CMRMoCC0sNC.RznR;
R-RR-CRtMNCs00CRE)CRqOvRC#DDR8NMRH0s-N#00
C#RRRRRRRRRRRRzR.(:FRVsRR[H5MRI0H8Ek_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0RC
RRRRRRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)RAqUv_4Xg..:7RRLDNCHDR#WR""R;
RRRRRRRRRRRRRLRRCMoH
RRRRRRRRRRRRRRRRqA)v4_Ug..X7RR:)Aqv41n_.._1
RRRRRRRRRRRRRRRRsbF0NRlb7R5Q=qR>MRH_osC5[.*+84RF0IMF*R.[R2,q)77q>R=RIDF_8IN84s5.FR8IFM0R,j2RA7QRR=>""jj,7Rq7R)A=D>RFsI_Ns885R4.8MFI0jFR2R,
RRRRRRRRRRRRR RRh=qR>4R''1,R1R)q='>RjR',WR q=I>RsC0_M25H,pRBi=qR>pRBi ,Rh=AR>4R''1,R1R)A='>RjR',WR A='>RjR',BApiRR=>B,pi
RRRRRRRRRRRRRRRRq7mRR=>FMbC,mR7A254RR=>F_k0L.k#5.H,*4[+27,RmjA52>R=R0Fk_#Lk.,5HR[.*2
2;RRRRRRRRRRRRRRRRF_k0s5Co.2*[RR<=F_k0L.k#5.H,*R[2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5[.*+R42<F=RkL0_k5#.H*,.[2+4RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRMRC8CRoMNCs0zCR.
(;RRRRRRRRCRM8oCCMsCN0Rcz.;R
RRMRC8CRoMNCs0zCR.Rd;RR

RRRRR-RR-CRtMNCs00CRE)CRqOvRC#DDR8NMRD#CCRO0DHFoOFRVsqR)vnA4__1c1Rc
RzRR.:URRRHV5FOEH_OCI0H8ERR=co2RCsMCN
0CRRRRRRRRzR.g:FRVsRRHH5MR80CbEk_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0RC
R-RR-VRQR85N8HsI8R0E>.R42CRMC08RFsROCCN0RHIs0CCRMDNLCMRN8kRF00bkRNCMLRDC#CCDOD0RFOoH
RRRRRRRRRRRRjzdRH:RVNR58I8sHE80R4>R.o2RCsMCN
0CRRRRRRRRRRRRRRRRF_k0CHM52=R<R''4RCIEM)R5q)77_b0l58N8s8IH04E-RI8FMR0F4R.2=2RHR#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=WI RERCM5_N8s5CoNs88I0H8ER-48MFI04FR.=2RRRH2CCD#R''j;R
RRRRRRRRRRMRC8CRoMNCs0zCRd
j;RRRR-Q-RVNR58I8sHE80RR<=4R.2MIFRsCH0RNCMLRDCFFsRkk0b0MRCNCLDRD#CCRO0DHFoOCRMC88C
RRRRRRRRRRRR4zdRH:RVNR58I8sHE80RR<=4R.2oCCMsCN0
RRRRRRRRRRRRRRRR0Fk_5CMH<2R=4R''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=W
 ;RRRRRRRRRRRRCRM8oCCMsCN0R4zd;R
RR-R-RMtCC0sNCER0CqR)vCRODRD#NRM80-sH#00NCR#
RRRRRRRRRzRRd:.RRsVFRH[RMIR5HE80_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNCR
RRRRRRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqA)vj_cgcnX7RR:DCNLD#RHR""W;R
RRRRRRRRRRRRRRCRLo
HMRRRRRRRRRRRRRRRRAv)q_gcjn7XcR):Rq4vAnc_1_
1cRRRRRRRRRRRRRRRRb0FsRblNRQ57q>R=R_HMs5Coc+*[dFR8IFM0R[c*2q,R7q7)RR=>D_FII8N8s454RI8FMR0FjR2,7RQA=">Rjjjj"q,R7A7)RR=>D_FIs8N8s454RI8FMR0Fj
2,RRRRRRRRRRRRRRRR Rhq='>R4R',1q1)RR=>',j'RqW RR=>I_s0CHM52B,RpRiq=B>RpRi, RhA='>R4R',1A1)RR=>',j'RAW RR=>',j'RiBpA>R=RiBp,R
RRRRRRRRRRRRRRmR7q>R=RCFbM7,RmdA52>R=R0Fk_#Lkc,5HR[c*+,d2RA7m5R.2=F>RkL0_k5#cH*,c[2+.,RR
RRRRRRRRRRRRR7RRm4A52>R=R0Fk_#Lkc,5Hc+*[4R2,75mAj=2R>kRF0k_L#Hc5,*Rc[;22
RRRRRRRRRRRRRRRR0Fk_osC5[c*2=R<R0Fk_#Lkc,5Hc2*[RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so*5c[2+4RR<=F_k0Lck#5cH,*4[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cco5*.[+2=R<R0Fk_#Lkc,5Hc+*[.I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Coc+*[d<2R=kRF0k_L#Hc5,[c*+Rd2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
R
RRRRRRRRRRMRC8CRoMNCs0zCRd
.;RRRRRRRRCRM8oCCMsCN0Rgz.;R
RRMRC8CRoMNCs0zCR.
U;
RRRRRRRRR--tCCMsCN0RC0ERv)qRDOCDN#RM#8RCODC0FRDoRHOVRFs)Aqv41n_gg_1
RRRRdzdRH:RVOR5EOFHCH_I8R0E=2RgRMoCC0sNCR
RRRRRRdRzcRR:VRFsHMRHRC58b_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
RRRRR--Q5VRNs88I0H8ERR>4R42M8CCRR0FONsC0ICRsCH0RNCMLRDCNRM8Fbk0kC0RMDNLCCR#D0CORoDFHRO
RRRRRRRRRzRRd:6RRRHV58N8s8IH0>ERR244RMoCC0sNCR
RRRRRRRRRRRRRRkRF0M_C5RH2<'=R4I'RERCM57)q70)_lNb58I8sHE80-84RF0IMF4R42RR=HC2RDR#C';j'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RWRCIEMNR58C_so85N8HsI8-0E4FR8IFM0R244RH=R2DRC#'CRj
';RRRRRRRRRRRRCRM8oCCMsCN0R6zd;R
RR-R-RRQV58N8s8IH0<ER=4R42FRMRHIs0CCRMDNLCsRFR0FkbRk0CLMND#CRCODC0FRDoRHOM8CCCR8
RRRRRRRRRzRRd:nRRRHV58N8s8IH0<ER=4R42CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_M25HRR<=';4'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RW;R
RRRRRRRRRRMRC8CRoMNCs0zCRd
n;RRRR-t-RCsMCNR0C0REC)RqvODCD#MRN8sR0H0-#N#0C
RRRRRRRRRRRR(zdRV:RF[sRRRHM58IH0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CRRRRRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FAVR)_qv.UjcXRU7:NRDLRCDH"#RW
";RRRRRRRRRRRRRRRRLHCoMR
RRRRRRRRRRRRRR)RAq.v_jXcUU:7RRv)qA_4n11g_gR
RRRRRRRRRRRRRRRRRb0FsRblNRQ57q>R=R_HMs5Cog+*[(FR8IFM0R[g*2q,R7q7)RR=>D_FII8N8sj54RI8FMR0FjR2,7RQA=">Rjjjjjjjj"q,R7A7)RR=>D_FIs8N8sj54RI8FMR0Fj
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRR Rhq='>R4R',1q1)RR=>',j'RqW RR=>I_s0CHM52B,RpRiq=B>RpRi, RhA='>R4R',1A1)RR=>',j'RAW RR=>',j'RiBpA>R=RiBp,RR
RRRRRRRRRRRRRRRRRRRRRRRRR7RRm=qR>bRFCRM,75mA(=2R>kRF0k_L#HU5,[U*+,(2RA7m5Rn2=F>RkL0_k5#UH*,U[2+n,RR
RRRRRRRRRRRRRRRRRRRRRRRRR7RRm6A52>R=R0Fk_#LkU,5HU+*[6R2,75mAc=2R>kRF0k_L#HU5,[U*+,c2RA7m5Rd2=F>RkL0_k5#UH*,U[2+d,RR
RRRRRRRRRRRRRRRRRRRRRRRRR7RRm.A52>R=R0Fk_#LkU,5HU+*[.R2,75mA4=2R>kRF0k_L#HU5,[U*+,42RA7m5Rj2=F>RkL0_k5#UH*,U[
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRR7qQu5Rj2=H>RMC_so*5g[2+U,QR7u=AR>jR""7,RmRuq=F>Rb,CMRu7mA25jRR=>bHNs0L$_k5#UH[,R2
2;RRRRRRRRRRRRRRRRF_k0s5Cog2*[RR<=F_k0LUk#5UH,*R[2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5[g*+R42<F=RkL0_k5#UH*,U[2+4RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so*5g[2+.RR<=F_k0LUk#5UH,*.[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cgo5*d[+2=R<R0Fk_#LkU,5HU+*[dI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cog+*[c<2R=kRF0k_L#HU5,[U*+Rc2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5[g*+R62<F=RkL0_k5#UH*,U[2+6RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so*5g[2+nRR<=F_k0LUk#5UH,*n[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cgo5*([+2=R<R0Fk_#LkU,5HU+*[(I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cog+*[U<2R=NRbs$H0_#LkU,5H[I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRCRM8oCCMsCN0R(zd;R
RRRRRRMRC8CRoMNCs0zCRd
c;RRRRCRM8oCCMsCN0Rdzd;R

RRRRR-RR-CRtMNCs00CRE)CRqOvRC#DDR8NMRD#CCRO0DHFoOFRVsqR)vnA4_U14_U14
RRRRUzdRH:RVOR5EOFHCH_I8R0E=UR42CRoMNCs0RC
RRRRRzRRd:gRRsVFRHHRM8R5CEb0_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNCR
RR-R-RRQV58N8s8IH0>ERR24jRCMC8FR0RCOsNR0CI0sHCMRCNCLDR8NMR0FkbRk0CLMND#CRCODC0FRDo
HORRRRRRRRRRRRzRcj:VRHR85N8HsI8R0E>jR42CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_M25HRR<='R4'IMECRq5)7_7)05lbNs88I0H8ER-48MFI04FRj=2RRRH2CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R ERIC5MRNs8_CNo58I8sHE80-84RF0IMFjR42RR=HC2RDR#C';j'
RRRRRRRRRRRR8CMRMoCC0sNCcRzjR;
R-RR-VRQR85N8HsI8R0E<4=RjM2RFsRIHR0CCLMNDFCRskRF00bkRNCMLRDC#CCDOD0RFOoHRCMC8
C8RRRRRRRRRRRRzRc4:VRHR85N8HsI8R0E<4=Rjo2RCsMCN
0CRRRRRRRRRRRRRRRRF_k0CHM52=R<R''4;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R R;
RRRRRRRRRCRRMo8RCsMCNR0Cz;c4
RRRRR--tCCMsCN0RC0ERv)qRDOCDN#RM08Rs#H-0CN0#R
RRRRRRRRRRcRz.RR:VRFs[MRHRH5I8_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
RRRRRRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVAv)q_.4jcnX47RR:DCNLD#RHR""W;R
RRRRRRRRRRRRRRCRLo
HMRRRRRRRRRRRRRRRRAv)q_.4jcnX47RR:)Aqv41n_41U_4RU
RRRRRRRRRRRRRRRRRsbF0NRlb7R5Q=qR>MRH_osC5*4U[6+4RI8FMR0F4[U*2q,R7q7)RR=>D_FII8N8sR5g8MFI0jFR27,RQ=AR>jR"jjjjjjjjjjjjj"jj,7Rq7R)A=D>RFsI_Ns8858gRF0IMF2Rj,R
RRRRRRRRRRRRRRRRRRRRRRRRRRhR q>R=R''4,1R1)=qR>jR''W,R =qR>sRI0M_C5,H2RiBpq>R=RiBp,hR A>R=R''4,1R1)=AR>jR''W,R =AR>jR''B,RpRiA=B>RpRi,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRq7mRR=>FMbC,mR7A6542>R=R0Fk_#Lk4Hn5,*4n[6+427,Rm4A5c=2R>kRF0k_L#54nHn,4*4[+cR2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRA7m524dRR=>F_k0L4k#n,5H4[n*+24d,mR7A.542>R=R0Fk_#Lk4Hn5,*4n[.+427,Rm4A54=2R>kRF0k_L#54nHn,4*4[+4R2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRA7m524jRR=>F_k0L4k#n,5H4[n*+24j,mR7A25gRR=>F_k0L4k#n,5H4[n*+,g2RA7m5RU2=F>RkL0_kn#454H,n+*[UR2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRA7m5R(2=F>RkL0_kn#454H,n+*[(R2,75mAn=2R>kRF0k_L#54nHn,4*n[+27,Rm6A52>R=R0Fk_#Lk4Hn5,*4n[2+6,RR
RRRRRRRRRRRRRRRRRRRRRRRRR7RRmcA52>R=R0Fk_#Lk4Hn5,*4n[2+c,mR7A25dRR=>F_k0L4k#n,5H4[n*+,d2RA7m5R.2=F>RkL0_kn#454H,n+*[.R2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRA7m5R42=F>RkL0_kn#454H,n+*[4R2,75mAj=2R>kRF0k_L#54nHn,4*,[2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRQR7u=qR>MRH_osC5*4U[(+4RI8FMR0F4[U*+24n,QR7u=AR>jR"j
",RRRRRRRRRRRRRRRRRRRRRRRRRRRR7qmuRR=>FMbC,mR7u4A52>R=RsbNH_0$L4k#n,5HR[.*+,42Ru7mA25jRR=>bHNs0L$_kn#45RH,.2*[2R;
RRRRRRRRRRRRRFRRks0_C4o5U2*[RR<=F_k0L4k#n,5H4[n*2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[4<2R=kRF0k_L#54nHn,4*4[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[.<2R=kRF0k_L#54nHn,4*.[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[d<2R=kRF0k_L#54nHn,4*d[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[c<2R=kRF0k_L#54nHn,4*c[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[6<2R=kRF0k_L#54nHn,4*6[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[n<2R=kRF0k_L#54nHn,4*n[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[(<2R=kRF0k_L#54nHn,4*([+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[U<2R=kRF0k_L#54nHn,4*U[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[g<2R=kRF0k_L#54nHn,4*g[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[4Rj2<F=RkL0_kn#454H,n+*[4Rj2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[4+42=R<R0Fk_#Lk4Hn5,*4n[4+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[4R.2<F=RkL0_kn#454H,n+*[4R.2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[d+42=R<R0Fk_#Lk4Hn5,*4n[d+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[4Rc2<F=RkL0_kn#454H,n+*[4Rc2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[6+42=R<R0Fk_#Lk4Hn5,*4n[6+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[4Rn2<b=RN0sH$k_L#54nH*,.[I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+24(RR<=bHNs0L$_kn#45.H,*4[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRCRRMo8RCsMCNR0Cz;c.
RRRRRRRR8CMRMoCC0sNCdRzgR;
RCRRMo8RCsMCNR0Cz;dU
R
RRRRRR-R-RMtCC0sNCER0CqR)vCRODRD#NRM8#CCDOD0RFOoHRsVFRv)qA_4n1_dn1
dnRRRRzNdURH:RVOR5EOFHCH_I8R0E=nRd2CRoMNCs0RC
RRRRRzRRdRgN:FRVsRRHH5MR80CbEk_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0RC
R-RR-VRQR85N8HsI8R0E>2RgRCMC8FR0RCOsNR0CI0sHCMRCNCLDR8NMR0FkbRk0CLMND#CRCODC0FRDo
HORRRRRRRRRRRRzNcjRH:RVNR58I8sHE80Rg>R2CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_M25HRR<='R4'IMECRq5)7_7)05lbNs88I0H8ER-48MFI0gFR2RR=HC2RDR#C';j'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RWRCIEMNR58C_so85N8HsI8-0E4FR8IFM0RRg2=2RHR#CDCjR''R;
RRRRRRRRRCRRMo8RCsMCNR0CzNcj;R
RR-R-RRQV58N8s8IH0<ER=2RgRRMFI0sHCMRCNCLDRRFsFbk0kC0RMDNLCCR#D0CORoDFHMORCCC88R
RRRRRRRRRRcRz4:NRRRHV58N8s8IH0<ER=2RgRMoCC0sNCR
RRRRRRRRRRRRRRkRF0M_C5RH2<'=R4
';RRRRRRRRRRRRRRRRI_s0CHM52=R<R;W 
RRRRRRRRRRRR8CMRMoCC0sNCcRz4
N;RRRR-t-RCsMCNR0C0REC)RqvODCD#MRN8sR0H0-#N#0C
RRRRRRRRRRRR.zcNRR:VRFs[MRHRH5I8_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
RRRRRRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVAv)q_.64X7d.RD:RNDLCRRH#";W"
RRRRRRRRRRRRRRRRoLCHRM
RRRRRRRRRRRRRARR)_qv6X4.dR.7:qR)vnA4_n1d_n1d
RRRRRRRRRRRRRRRRbRRFRs0lRNb5q7QRR=>HsM_Cdo5n+*[d84RF0IMFnRd*,[2R7q7)=qR>FRDIN_I858sUFR8IFM0R,j2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRQR7A>R=Rj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjj,j"R7q7)=AR>FRDIN_s858sUFR8IFM0R,j2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRq hRR=>',4'R)11q>R=R''j, RWq>R=R0Is_5CMHR2,BqpiRR=>B,piRA hRR=>',4'R)11A>R=R''j, RWA>R=R''j,pRBi=AR>pRBi
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRR7Rmq=F>Rb,CMRA7m52d4RR=>F_k0Ldk#.,5Hd[.*+2d4,mR7Aj5d2>R=R0Fk_#LkdH.5,*d.[j+d2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mA.Rg2=F>RkL0_k.#d5dH,.+*[.,g2RA7m52.URR=>F_k0Ldk#.,5Hd[.*+2.U,mR7A(5.2>R=R0Fk_#LkdH.5,*d.[(+.2R,
RRRRRRRRRRRRRRRRRRRRRRRRR7RRm.A5n=2R>kRF0k_L#5d.H.,d*.[+nR2,75mA.R62=F>RkL0_k.#d5dH,.+*[.,62RA7m52.cRR=>F_k0Ldk#.,5Hd[.*+2.c,R
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7Ad5.2>R=R0Fk_#LkdH.5,*d.[d+.27,Rm.A5.=2R>kRF0k_L#5d.H.,d*.[+.R2,75mA.R42=F>RkL0_k.#d5dH,.+*[.,42
RRRRRRRRRRRRRRRRRRRRRRRRRRRRA7m52.jRR=>F_k0Ldk#.,5Hd[.*+2.j,mR7Ag542>R=R0Fk_#LkdH.5,*d.[g+427,Rm4A5U=2R>kRF0k_L#5d.H.,d*4[+U
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRR75mA4R(2=F>RkL0_k.#d5dH,.+*[4,(2RA7m524nRR=>F_k0Ldk#.,5Hd[.*+24n,mR7A6542>R=R0Fk_#LkdH.5,*d.[6+42R,
RRRRRRRRRRRRRRRRRRRRRRRRR7RRm4A5c=2R>kRF0k_L#5d.H.,d*4[+cR2,75mA4Rd2=F>RkL0_k.#d5dH,.+*[4,d2RA7m524.RR=>F_k0Ldk#.,5Hd[.*+24.,RR
RRRRRRRRRRRRRRRRRRRRRRRRR7RRm4A54=2R>kRF0k_L#5d.H.,d*4[+4R2,75mA4Rj2=F>RkL0_k.#d5dH,.+*[4,j2RA7m5Rg2=F>RkL0_k.#d5dH,.+*[gR2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRA7m5RU2=F>RkL0_k.#d5dH,.+*[UR2,75mA(=2R>kRF0k_L#5d.H.,d*([+27,RmnA52>R=R0Fk_#LkdH.5,*d.[2+n,RR
RRRRRRRRRRRRRRRRRRRRRRRRR7RRm6A52>R=R0Fk_#LkdH.5,*d.[2+6,mR7A25cRR=>F_k0Ldk#.,5Hd[.*+,c2RA7m5Rd2=F>RkL0_k.#d5dH,.+*[dR2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRA7m5R.2=F>RkL0_k.#d5dH,.+*[.R2,75mA4=2R>kRF0k_L#5d.H.,d*4[+27,RmjA52>R=R0Fk_#LkdH.5,*d.[R2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRu7Qq>R=R_HMs5Cod[n*+Rd68MFI0dFRn+*[d,.2Ru7QA>R=Rj"jj,j"Ru7mq>R=RCFbM7,Rm5uAd=2R>NRbs$H0_#LkdH.5,[c*+,d2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7u.A52>R=RsbNH_0$Ldk#.,5Hc+*[.R2,7Amu5R42=b>RN0sH$k_L#5d.H*,c[2+4,mR7ujA52>R=RsbNH_0$Ldk#.,5Hc2*[2R;
RRRRRRRRRRRRRFRRks0_Cdo5n2*[RR<=F_k0Ldk#.,5Hd[.*2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cdo5n+*[4<2R=kRF0k_L#5d.H.,d*4[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cdo5n+*[.<2R=kRF0k_L#5d.H.,d*.[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cdo5n+*[d<2R=kRF0k_L#5d.H.,d*d[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cdo5n+*[c<2R=kRF0k_L#5d.H.,d*c[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cdo5n+*[6<2R=kRF0k_L#5d.H.,d*6[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cdo5n+*[n<2R=kRF0k_L#5d.H.,d*n[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cdo5n+*[(<2R=kRF0k_L#5d.H.,d*([+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cdo5n+*[U<2R=kRF0k_L#5d.H.,d*U[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cdo5n+*[g<2R=kRF0k_L#5d.H.,d*g[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cdo5n+*[4Rj2<F=RkL0_k.#d5dH,.+*[4Rj2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*dn[4+42=R<R0Fk_#LkdH.5,*d.[4+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cdo5n+*[4R.2<F=RkL0_k.#d5dH,.+*[4R.2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*dn[d+42=R<R0Fk_#LkdH.5,*d.[d+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cdo5n+*[4Rc2<F=RkL0_k.#d5dH,.+*[4Rc2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*dn[6+42=R<R0Fk_#LkdH.5,*d.[6+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cdo5n+*[4Rn2<F=RkL0_k.#d5dH,.+*[4Rn2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*dn[(+42=R<R0Fk_#LkdH.5,*d.[(+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cdo5n+*[4RU2<F=RkL0_k.#d5dH,.+*[4RU2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*dn[g+42=R<R0Fk_#LkdH.5,*d.[g+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cdo5n+*[.Rj2<F=RkL0_k.#d5dH,.+*[.Rj2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*dn[4+.2=R<R0Fk_#LkdH.5,*d.[4+.2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cdo5n+*[.R.2<F=RkL0_k.#d5dH,.+*[.R.2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*dn[d+.2=R<R0Fk_#LkdH.5,*d.[d+.2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cdo5n+*[.Rc2<F=RkL0_k.#d5dH,.+*[.Rc2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*dn[6+.2=R<R0Fk_#LkdH.5,*d.[6+.2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cdo5n+*[.Rn2<F=RkL0_k.#d5dH,.+*[.Rn2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*dn[(+.2=R<R0Fk_#LkdH.5,*d.[(+.2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cdo5n+*[.RU2<F=RkL0_k.#d5dH,.+*[.RU2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*dn[g+.2=R<R0Fk_#LkdH.5,*d.[g+.2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cdo5n+*[dRj2<F=RkL0_k.#d5dH,.+*[dRj2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*dn[4+d2=R<R0Fk_#LkdH.5,*d.[4+d2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cdo5n+*[dR.2<b=RN0sH$k_L#5d.H*,c[I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cod[n*+2ddRR<=bHNs0L$_k.#d5cH,*4[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cdo5n+*[dRc2<b=RN0sH$k_L#5d.H*,c[2+.RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_son5d*d[+6<2R=NRbs$H0_#LkdH.5,[c*+Rd2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRR8CMRMoCC0sNCcRz.
N;RRRRRRRRCRM8oCCMsCN0RgzdNR;
RCRRMo8RCsMCNR0CzNdU;R
RCRM8oCCMsCN0Rdzc;R
Rz:ccRRHV50MFR8N8sC_soo2RCsMCNR0C-o-RCsMCNR0C#CCDOs0RNRl
R-RR-VRQR8N8s8IH0<ERRN(R#o#HMjR''FR0RkkM#RC8L#H0
RRRRRzjRH:RVNR58I8sHE80R4=R2CRoMNCs0RC
RRRRRDRRFNI_8R8s<"=RjjjjjRj"&_R#Ns8_Cjo52R;
RCRRMo8RCsMCNR0Cz
j;RRRRzR4R:VRHR85N8HsI8R0E=2R.RMoCC0sNCR
RRRRRRFRDI8_N8<sR=jR"jjjj"RR&#8_N_osC584RF0IMF2Rj;R
RRMRC8CRoMNCs0zCR4R;
RzRR.:RRRRHV58N8s8IH0=ERRRd2oCCMsCN0
RRRRRRRRIDF_8N8s=R<Rj"jjRj"&_R#Ns8_C.o5RI8FMR0Fj
2;RRRRCRM8oCCMsCN0R;z.
RRRRRzdRH:RVNR58I8sHE80Rc=R2CRoMNCs0RC
RRRRRDRRFNI_8R8s<"=Rj"jjR#&R__N8s5CodFR8IFM0R;j2
RRRR8CMRMoCC0sNCdRz;z
ScRS:H5VRNs88I0H8ERR=6o2RCsMCN
0CSFSDI8_N8<sR=jR"j&"RRN#_8C_soR5c8MFI0jFR2S;
CRM8oCCMsCN0R;zc
6SzSH:RVNR58I8sHE80Rn=R2CRoMNCs0SC
SIDF_8N8s=R<R''jR#&R__N8s5Co6FR8IFM0R;j2
RRRR8CMRMoCC0sNC6Rz;R
RRnRzRRR:H5VRNs88I0H8ERR>no2RCsMCN
0CRRRRRRRRD_FINs88RR<=#8_N_osC58nRF0IMF2Rj;R
RRMRC8CRoMNCs0zCRn
;
RRRR-Q-RV8R5HsM_CRo2sHCo#s0CRh7QRHk#MBoRpRi
RzRR(:RRRRHV5M8H_osC2CRoMNCs0RC
RRRRRbRRsCFO#5#RB,piRh7Q2CRLo
HMRRRRRRRRRRRRH5VRBRpi=4R''MRN8pRBiP'CC2M0RC0EMR
RRRRRRRRRRRRRR_R#HsM_C<oR=QR7hR;
RRRRRRRRRCRRMH8RVR;
RRRRRCRRMb8RsCFO#
#;RRRRCRM8oCCMsCN0R;z(
RRRRRzURH:RVMR5F80RHsM_CRo2oCCMsCN0
RRRRRRRRRRRRH#_MC_so=R<Rh7Q;R
RRMRC8CRoMNCs0zCRU
;
RRRR-Q-RV8R5F_k0s2CoRosCHC#0smR7zkaR#oHMRpmBiR
RRgRzRRR:H5VR80Fk_osC2CRoMNCs0RC
RRRRRbRRsCFO#5#RmiBp,kRF0C_soL2RCMoH
RRRRRRRRRRRRRHV5pmBiRR='R4'NRM8miBp'CCPMR020MEC
RRRRRRRRRRRRRRRRz7ma=R<RF#_ks0_C
o;RRRRRRRRRRRRCRM8H
V;RRRRRRRRCRM8bOsFC;##
RRRR8CMRMoCC0sNCgRz;R
RR4Rzj:RRRRHV50MFRk8F0C_soo2RCsMCN
0CRRRRRRRRRRRR7amzRR<=#k_F0C_soR;
RCRRMo8RCsMCNR0Cz;4j
R
RR-R-RRQV58N8sC_sos2RC#oH0RCsq)77RHk#MBoRpRi
RzRR4R4R:VRHR85N8ss_CRo2oCCMsCN0
RRRRRRRRFbsO#C#Rp5Biq,R727)RoLCHRM
RRRRRRRRRHRRVBR5p=iRR''4R8NMRiBp'CCPMR020MEC
RRRRRRRRRRRRRRRRN#_8C_so=R<R7q7)85N8HsI8-0E4FR8IFM0R;j2
RRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMRFbsO#C#;R
RRMRC8CRoMNCs0zCR4
4;RRRRzR4.:VRHRF5M08RN8ss_CRo2oCCMsCN0
RRRRRRRRRRRRN#_8C_so=R<R7q7)R;
RCRRMo8RCsMCNR0Cz;4.
RRRRRRRRR
RR-R-RMtCC0sNCER0CqR)vCRODRD#NRM8#CCDOD0RFOoH
RRRRdz4RV:RFHsRRRHM5lMk_DOCD._4URR-482RF0IMFRRjoCCMsCN0
RRRRR--Q5VRNs88I0H8ERR>6M2RCRC80OFRs0CNCsRIHR0CCLMNDNCRMF8Rkk0b0MRCNCLDRD#CCRO0DHFoOR
RRRRRR4RzcRR:H5VRNs88I0H8ERR>(o2RCsMCN
0CRRRRRRRRRRRRRRRR#k_F0M_C5RH2<'=R4I'RERCM5N#_8C_so85N8HsI8-0E4FR8IFM0RR(2=2RHR#CDCjR''R;
RRRRRRRRRRRRR#RR_0Is_5CMH<2R= RWRCIEM#R5__N8s5CoNs88I0H8ER-48MFI0(FR2RR=HC2RDR#C';j'
RRRRRRRR8CMRMoCC0sNC4RzcR;
R-RR-VRQR85N8HsI8R0E<6=R2FRMRHIs0CCRMDNLCsRFR0FkbRk0CLMND#CRCODC0FRDoRHOM8CCCR8
RRRRRzRR4:6RRRHV58N8s8IH0<ER=2R(RMoCC0sNCR
RRRRRRRRRRRRRR_R#F_k0CHM52=R<R''4;R
RRRRRRRRRRRRRR_R#I_s0CHM52=R<R;W 
RRRRRRRR8CMRMoCC0sNC4Rz6R;
R-RR-CRtMNCs00CRE)CRqOvRC#DDR8NMRH0s-N#00
C#RRRRRRRRzR4n:FRVsRR[H5MRI0H8ERR-482RF0IMFRRjoCCMsCN0
RRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVzv)q4R.U:NRDLRCDH"#R1"1aRH&RMo0CCHs'lCNo58IH0RE2&7R""RR&HCM0o'CsHolNC*5H42.UR"&RW&"RR0HMCsoC'NHlo[C52RR&"R "&MRH0CCosl'HN5oCo_C0C_M880CbEH55+*424,.URb8C02E2R"&RX&"RR0HMCsoC'NHlo[C5+;42
RRRRRRRRRRRRoLCHRM
RRRRRRRRRzRR)4qv.:URRqX)vU4.XR41
RRRRRRRRRRRRRRRRsbF0NRlb7R5RR=>#M_H_osC5,[2RRqj=D>RFNI_858sjR2,q=4R>FRDI8_N84s52q,R.>R=RIDF_8N8s25.,R
RRRRRRRRRRRRRRRRRRRRRRRRRq=dR>FRDI8_N8ds52q,Rc>R=RIDF_8N8s25c,6RqRR=>D_FINs885,62RRqn=D>RFNI_858sn
2,SSSSSRSRW= R>_R#I_s0CHM52W,RBRpi=B>RpRi,m>R=R0Fk_#Lk_U4.5[H,2
2;RRRRRRRRRRRRRRRR#k_F0C_so25[RR<=F_k0L_k#45.UH2,[RCIEM#R5_0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRCRM8oCCMsCN0Rnz4;R
RRCRRMo8RCsMCNR0Cz;4dRRRRRRRRRRRR
RRRR
RRRRRR-t-RCsMCNR0CNnR4RsIF8CR8C)bRqOvRCRDDHNVRbFbsbNsH0RCRRRRRRRRRRRRRRR
RR4Rz(RR:H5VRM_klODCD_Rnc=2R4RMoCC0sNCR
RR-R-RRQV58N8s8IH0>ERRR(2M8CCRR0FONsC0ICRsCH0RNCMLRDCNRM8Fbk0kC0RMDNLCCR#D0CORoDFHRO
RRRRRzRR4RUN:VRHR85N8HsI8R0E>2R(RMoCC0sNCR
RRRRRRRRRRRRRRkRF0M_C_Rnc<'=R4I'RERCM5_5#Ns8_CNo58I8sHE80-84RF0IMF2R(RM=RkOl_C_DD42.UR8NMR_5#Ns8_Cno52RR='2j'2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0CnM_c=R<RRW IMECR#55__N8s5CoNs88I0H8ER-48MFI0(FR2RR=M_klODCD_U4.2MRN8#R5__N8s5Con=2RR''j2C2RDR#C';j'
RRRRRRRR8CMRMoCC0sNC4RzU
N;RRRRRRRRzL4URH:RVNR58I8sHE80R(=RR8NMRlMk_DOCD._4URR=jo2RCsMCN
0CRRRRRRRRRRRRRRRRF_k0CnM_c=R<R''4RCIEM5R5#8_N_osC5Rn2=jR''R22CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C_Rnc<W=R ERIC5MR5N#_8C_so25nR'=Rj2'2R#CDCjR''R;
RRRRRCRRMo8RCsMCNR0CzL4U;R
RR-R-RRQV58N8s8IH0<ER=2R6RRMFI0sHCMRCNCLDRRFsFbk0kC0RMDNLCCR#D0CORoDFHMORCCC88R
RRRRRR4RzgRR:H5VRNs88I0H8E=R<RRn2oCCMsCN0
RRRRRRRRRRRRRRRR0Fk__CMn<cR=4R''R;
RRRRRRRRRRRRRIRRsC0_Mc_nRR<=W
 ;RRRRRRRRCRM8oCCMsCN0Rgz4;R
RR-R-RMtCC0sNCER0CqR)vCRODNDRM08Rs#H-0CN0
RSRRORzE.	_RH:RV#R5_8IH0NE_s$sN_5nc4>2RRRj2oCCMsCN0
RRRRRRRRjz.RV:RF[sRRRHM5I#_HE80_sNsNn$_c254R4-R2FR8IFM0RojRCsMCN
0CRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FzVR)nqvcRR:DCNLD#RHR1"1a&"RR0HMCsoC'NHloIC5HE802RR&"R7"&MRH0CCosl'HN5oCM_klODCD_U4.*U4.2RR&"RW"&MRH0CCosl'HN5oCI0H8ERR-.R*[-2R.R"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05lMk_DOCD._4U.*4URR+nRc,80CbER22&XR""RR&HCM0o'CsHolNCH5I8R0E-*R.[
2;RRRRRRRRRRRRLHCoMR
RRRRRRRRRR)RzqcvnRX:R)nqvc1X.RR
RRRRRRRRRRRRRRFRbsl0RN5bR7=4R>_R#HsM_CIo5HE80-[.*-,42RR7j=#>R__HMs5CoI0H8E*-.[2-.,jRqRR=>D_FINs885,j2RRq4=D>RFNI_858s4R2,q=.R>FRDI8_N8.s52R,
RRRRRRRRRRRRRRRRRRRRRRRRRRqd=D>RFNI_858sdR2,q=cR>FRDI8_N8cs52q,R6>R=RIDF_8N8s256,S
SSSSSR RWRR=>I_s0CnM_cW,RBRpi=B>RpRi,m=4R>kRF0k_L#c_n5lMk_DOCDc_n,8IH0.E-*4[-2m,Rj>R=R0Fk_#Lk_5ncM_klODCD_,ncI0H8E*-.[2-.2R;
RRRRRRRRRRRRR#RR_0Fk_osC58IH0.E-*4[-2=R<R0Fk_#Lk_5ncM_klODCD_,ncI0H8E*-.[2-4RCIEMFR5kC0_Mc_nR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRR_R#F_k0s5CoI0H8E*-.[2-.RR<=F_k0L_k#nMc5kOl_C_DDnIc,HE80-[.*-R.2IMECRk5F0M_C_Rnc=4R''C2RDR#C';Z'
RRRRRRRRMRC8CRoMNCs0zCR.
j;SCSRMo8RCsMCNR0Cz	OE_
.;SzSRO_E	4RR:H5VR#H_I8_0ENNss$c_n5Rj2>2RjRMoCC0sNCR
RRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqz)vRnc:NRDLRCDH"#R1"1aRH&RMo0CCHs'lCNo58IH0RE2&7R""RR&HCM0o'CsHolNCk5MlC_OD4D_.4U*.RU2&WR""RR&HCM0o'CsHolNCH5I8R0E-*R.#H_I8_0ENNss$c_n5R42-2R4R"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05lMk_DOCD._4U.*4URR+nRc,80CbER22&XR""RR&HCM0o'CsHolNCH5I8R0E-*R.#H_I8_0ENNss$c_n5242;R
RRRRRRRRRRCRLo
HMRRRRRRRRRRRRzv)qn:cRRv)qn4cX1RR
RRRRRRRRRRRRRbRRFRs0lRNb5=7R>_R#HsM_CIo5HE80-#.*_8IH0NE_s$sN_5nc442-2q,Rj>R=RIDF_8N8s25j,4RqRR=>D_FINs885,42RRq.=D>RFNI_858s.
2,RRRRRRRRRRRRRRRRRRRRRRRRRdRqRR=>D_FINs885,d2RRqc=D>RFNI_858scR2,q=6R>FRDI8_N86s52S,
SSSSSWRR >R=R0Is__CMnRc,WiBpRR=>B,piR=mR>kRF0k_L#c_n5lMk_DOCDc_n,8IH0.E-*I#_HE80_sNsNn$_c254-242;R
RRRRRRRRRRRRRR_R#F_k0s5CoI0H8E*-.#H_I8_0ENNss$c_n5-424<2R=kRF0k_L#c_n5lMk_DOCDc_n,8IH0.E-*I#_HE80_sNsNn$_c254-R42IMECRk5F0M_C_Rnc=4R''C2RDR#C';Z'
RRRRRRRRMRC8CRoMNCs0zCRO_E	4S;
RRRRR8CMRMoCC0sNC4Rz(R;RRRRRRRRR
R
RR-R-RMtCC0sNCRRN4InRFRs88bCCRv)qRDOCDVRHRbNbssFbHCN0RRRRRRRRRRRRR
RRRRRRzR.4:VRHRk5MlC_ODdD_.RR=4o2RCsMCN
0CRRRR-Q-RVNR58I8sHE80R6>R2CRMC08RFsROCCN0RHIs0CCRMDNLCMRN8kRF00bkRNCMLRDC#CCDOD0RFOoH
RRRRRRRR.z.NRR:H5VRNs88I0H8ERR>(MRN8kRMlC_ODnD_cRR=4o2RCsMCN
0CRRRRRRRRRRRRRRRRF_k0CdM_.=R<R''4RCIEM5R5#8_N_osC58N8s8IH04E-RI8FMR0F(=2RRlMk_DOCD._4UN2RM58R#8_N_osC5Rn2=4R''N2RM58R#8_N_osC5R62=jR''R22CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C_Rd.<W=R ERIC5MR5N#_8C_so85N8HsI8-0E4FR8IFM0RR(2=kRMlC_OD4D_.RU2NRM85N#_8C_so25nR'=R4R'2NRM85N#_8C_so256R'=Rj2'2R#CDCjR''R;
RRRRRCRRMo8RCsMCNR0CzN..;R
RRRRRR.Rz.:LRRRHV58N8s8IH0>ERRN(RMM8RkOl_C_DDn/cR=2R4RMoCC0sNCR
RRRRRRRRRRRRRRkRF0M_C_Rd.<'=R4I'RERCM5_5#Ns8_CNo58I8sHE80-84RF0IMF2R(RM=RkOl_C_DD42.UR8NMR_5#Ns8_Cno52RR='2j'R8NMR_5#Ns8_C6o52RR='2j'2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0CdM_.=R<RRW IMECR#55__N8s5CoNs88I0H8ER-48MFI0(FR2RR=M_klODCD_U4.2MRN8#R5__N8s5Con=2RR''j2MRN8#R5__N8s5Co6=2RR''j2C2RDR#C';j'
RRRRRRRR8CMRMoCC0sNC.Rz.
L;RRRRRRRRzO..RH:RVNR58I8sHE80R(=RR8NMRlMk_DOCDc_nR4=R2CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_M._dRR<='R4'IMECR#55__N8s5Con=2RR''42MRN8#R5__N8s5Co6=2RR''j2C2RDR#C';j'
RRRRRRRRRRRRRRRR0Is__CMd<.R= RWRCIEM5R5#8_N_osC5Rn2=4R''N2RM58R#8_N_osC5R62=jR''R22CCD#R''j;R
RRRRRRMRC8CRoMNCs0zCR.;.O
RRRRRRRR.z.8RR:H5VRNs88I0H8ERR=nMRN8kRMlC_ODnD_c=R/RR42oCCMsCN0
RRRRRRRRRRRRRRRR0Fk__CMd<.R=4R''ERIC5MR5N#_8C_so85N8HsI8-0E4FR8IFM0RR62=kRMlC_ODnD_cR22CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C_Rd.<W=R ERIC5MR5N#_8C_so85N8HsI8-0E4FR8IFM0RR62=kRMlC_ODnD_cR22CCD#R''j;R
RRRRRRMRC8CRoMNCs0zCR.;.8
RRRRR--Q5VRNs88I0H8E=R<RR62MIFRsCH0RNCMLRDCFFsRkk0b0MRCNCLDRD#CCRO0DHFoOCRMC88C
RRRRRRRRdz.RH:RVNR58I8sHE80RR<=6o2RCsMCN
0CRRRRRRRRRRRRRRRRF_k0CdM_.=R<R''4;R
RRRRRRRRRRRRRRsRI0M_C_Rd.<W=R R;
RRRRRCRRMo8RCsMCNR0Cz;.d
RRRRR--tCCMsCN0RC0ERv)qRDOCDMRN8sR0H0-#N
0CSRRRREzO	R_U:VRHR_5#I0H8Es_Ns5N$d>2RRRj2oCCMsCN0
zSSO_E	DRC6:VRHRH5I8R0E>U=R*I#_HE80_sNsNd$52MRN8HRI8R0E>U=R2CRoMNCs0RC
RRRRRRRRRRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)Rzq.vdRD:RNDLCRRH#"a11"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloMC5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*n2RR&"RW"&MRH0CCosl'HN5oCI0H8ERR-D_#LI0H8E&2RR"" RH&RMo0CCHs'lCNo50oC_8CM_b8C0ME5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*nRd+R.8,RCEb02&2RR""XRH&RMo0CCHs'lCNo58IH0-ERRLD#_8IH0+ERR;U2
RRRRRRRRRRRRRRRRRRRRoLCHSM
SRRRRqz)vRd.:)RXq.vdX
U1SRSSRbRRFRs0lRNb5=7R>NRb8_5#HsM_CIo5HE80-84RF0IMFHRI8-0ED_#LI0H8ER2,UD,R#IL_HE80-,42RRqj=D>RFNI_858sj
2,SSSSSRSRq=4R>FRDI8_N84s52q,R.>R=RIDF_8N8s25.,dRqRR=>D_FINs885,d2RRqc=D>RFNI_858scR2,W= R>sRI0M_C_,d.RpWBi>R=RiBp,S
SSSSSRRRm=0>RlUb__5d.j;22
SSSS#N#HRoM:FRVs[RHRRHMI0H8ER-48MFI0IFRHE80-LD#_8IH0oERCsMCN
0CSSSSRkRF0k_L#._d5lMk_DOCD._d,2H[RR<=0_lbU._d55j2HI[-HE80+LD#_8IH0;E2
RRRRRRRRRRRRRRRR#RR_0Fk_osC52H[RR<=F_k0L_k#dM.5kOl_C_DDdH.,[I2RERCM50Fk__CMd=.RR''42DRC#'CRZ
';SSSSCRM8oCCMsCN0R#N#H;oM
RRRRRRRRRRRRUz.RV:RF[sRRRHM#H_I8_0ENNss$25d-84RF0IMFRR4oCCMsCN0
RRRRRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)Rzq.vdRD:RNDLCRRH#"a11"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloMC5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*n2RR&"RW"&MRH0CCosl'HN5oCI0H8ERR-D_#LI0H8ERR-[2*UR"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05lMk_DOCD._4U.*4URR+M_klODCD_*ncn+cRR,d.Rb8C02E2R"&RX&"RR0HMCsoC'NHloIC5HE80RD-R#IL_HE80R5-R[2-4*;U2
RRRRRRRRRRRRLRRCMoH
RRRRRRRRRRRRzRR)dqv.RR:Xv)qdU.X1RR
RRRRRRRRRRRRRbRRFRs0lRNb5=7R>_R#HsM_CIo5HE80-LD#_8IH0UE-*([+RI8FMR0FI0H8E#-DLH_I8-0EU2*[,jRqRR=>D_FINs885,j2RRq4=D>RFNI_858s4R2,q=.R>FRDI8_N8.s52R,
RRRRRRRRRRRRRRRRRRRRRRRRRRqd=D>RFNI_858sdR2,q=cR>FRDI8_N8cs52W,R >R=R0Is__CMdR.,WiBpRR=>B,piR=mR>lR0b__Ud[.52
2;SRSSRNRR#o#HMRR:VRFsHH[RMRR(8MFI0jFRRMoCC0sNCS
SSRSRF_k0L_k#dM.5kOl_C_DDdI.,HE80-LD#_8IH0UE-*H[+[<2R=lR0b__Ud[.52[5H2R;
RRRRRRRRRRRRRRRRRF#_ks0_CIo5HE80-LD#_8IH0UE-*H[+[<2R=kRF0k_L#._d5lMk_DOCD._d,8IH0DE-#IL_HE80-[U*+2H[RCIEMFR5kC0_M._dR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRMRC8CRoMNCs0NCR#o#HMR;
RRRRRRRRRCRRMo8RCsMCNR0Cz;.U
CSSMo8RCsMCNR0Cz	OE_6DC;S
Sz	OE_6o0RH:RVIR5HE80RR>=UMRN8HRI8R0ElRF8U=R>RR62oCCMsCN0
RRRRRRRRRRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVzv)qd:.RRLDNCHDR#1R"1Ra"&MRH0CCosl'HN5oCI0H8E&2RR""7RH&RMo0CCHs'lCNo5lMk_DOCD._4U.*4URR+M_klODCD_*ncnRc2&WR""RR&HCM0o'CsHolNCH5I8R0E-#RDLH_I820ER"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05lMk_DOCD._4U.*4URR+M_klODCD_*ncn+cRR,d.Rb8C02E2R"&RX&"RR0HMCsoC'NHloIC5HE80RD-R#IL_HE80RU+R2R;
RRRRRRRRRRRRRRRRRLRRCMoH
RSSRzRR)dqv.RR:Xv)qdU.X1S
SSRRRRsbF0NRlb7R5RR=>b5N8#M_H_osC58IH04E-RI8FMR0FI0H8E#-DLH_I820E,,RURLD#_8IH04E-2q,Rj>R=RIDF_8N8s25j,S
SSSSSR4RqRR=>D_FINs885,42RRq.=D>RFNI_858s.R2,q=dR>FRDI8_N8ds52q,Rc>R=RIDF_8N8s25c, RWRR=>I_s0CdM_.W,RBRpi=B>Rp
i,SSSSSRSRm>R=Rb0l_dU_._5#I0H8Es_Ns5N$d42-2
2;SSSSNH##o:MRRsVFRRH[HIMRHE80-84RF0IMFHRI8-0ED_#LI0H8ECRoMNCs0SC
SRSSR0Fk_#Lk_5d.M_klODCD_,d.HR[2<0=RlUb__5d.#H_I8_0ENNss$25d-542HI[-HE80+LD#_8IH0;E2
RRRRRRRRRRRRRRRR#RR_0Fk_osC52H[RR<=F_k0L_k#dM.5kOl_C_DDdH.,[I2RERCM50Fk__CMd=.RR''42DRC#'CRZ
';SSSSCRM8oCCMsCN0R#N#H;oM
RRRRRRRRRRRRUz.RV:RF[sRRRHM#H_I8_0ENNss$25d-8.RF0IMFRRjoCCMsCN0
RRRRRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)Rzq.vdRD:RNDLCRRH#"a11"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloMC5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*n2RR&"RW"&MRH0CCosl'HN5oC[2*UR"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05lMk_DOCD._4U.*4URR+M_klODCD_*ncn+cRR,d.Rb8C02E2R"&RX&"RR0HMCsoC'NHlo5C5[2+4*;U2
RRRRRRRRRRRRLRRCMoH
RRRRRRRRRRRRzRR)dqv.RR:Xv)qdU.X1RR
RRRRRRRRRRRRRbRRFRs0lRNb5=7R>_R#HsM_CUo5*([+RI8FMR0FU2*[,jRqRR=>D_FINs885,j2RRq4=D>RFNI_858s4R2,q=.R>FRDI8_N8.s52R,
RRRRRRRRRRRRRRRRRRRRRRRRRRqd=D>RFNI_858sdR2,q=cR>FRDI8_N8cs52W,R >R=R0Is__CMdR.,WiBpRR=>B,piR=mR>lR0b__Ud[.52
2;SSSSNH##o:MRRsVFRRH[H(MRRI8FMR0FjCRoMNCs0SC
SRSSR0Fk_#Lk_5d.M_klODCD_,d.U+*[HR[2<0=RlUb__5d.[H25[
2;RRRRRRRRRRRRRRRRR_R#F_k0s5CoU+*[HR[2<F=RkL0_kd#_.k5MlC_ODdD_.*,U[[+H2ERIC5MRF_k0CdM_.RR='24'R#CDCZR''R;
RRRRRRRRRRRRRCRRMo8RCsMCNR0CNH##o
M;RRRRRRRRRRRRCRM8oCCMsCN0RUz.;S
SCRM8oCCMsCN0REzO	0_o6S;
SEzO	R_M:VRHRH5I8R0E<2RURMoCC0sNCR
RRRRRRRRRRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqz)vRd.:NRDLRCDH"#R1"1aRH&RMo0CCHs'lCNo58IH0RE2&7R""RR&HCM0o'CsHolNCk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*2ncR"&RW&"RR0HMCsoC'NHlojC52RR&"R "&MRH0CCosl'HN5oCo_C0C_M880CbEk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*Rnc+.Rd,CR8b20E2RR&"RX"&MRH0CCosl'HN5oCU
2;RRRRRRRRRRRRRRRRRRRRLHCoMS
SRRRRzv)qd:.RRqX)vXd.US1
SRSRRFRbsl0RN5bR7>R=R8bN5H#_MC_soH5I8-0E4FR8IFM0R8IH0DE-#IL_HE802U,R,#RDLH_I8-0E4R2,q=jR>FRDI8_N8js52S,
SSSSSqRR4>R=RIDF_8N8s254,.RqRR=>D_FINs885,.2RRqd=D>RFNI_858sdR2,q=cR>FRDI8_N8cs52W,R >R=R0Is__CMdR.,WiBpRR=>B,pi
SSSSRSSR=mR>lR0b__Udj.52
2;SSSSNH##o:MRRsVFRRH[HIMRHE80-84RF0IMFRRjoCCMsCN0
SSSSFRRkL0_kd#_.k5MlC_ODdD_.[,H2=R<Rb0l_dU_.25j52H[;R
RRRRRRRRRRRRRRRRR#k_F0C_so[5H2=R<R0Fk_#Lk_5d.M_klODCD_,d.HR[2IMECRk5F0M_C_Rd.=4R''C2RDR#C';Z'
SSSS8CMRMoCC0sNC#RN#MHo;S
SCRM8oCCMsCN0REzO	;_M
CSSMo8RCsMCNR0Cz	OE_
U;SOSzEc	_RH:RV#R5_8IH0NE_s$sN5R.2>2RjRMoCC0sNCR
RRRRRR.RzcR_c:VRHRH5I8R0E>c=R2CRoMNCs0RC
RRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)Rzq.vdRD:RNDLCRRH#"a11"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloMC5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*n2RR&"RW"&MRH0CCosl'HN5oCj&2RR"" RH&RMo0CCHs'lCNo50oC_8CM_b8C0ME5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*nRd+R.8,RCEb02&2RR""XRH&RMo0CCHs'lCNo5;c2
RRRRRRRRRRRRoLCHRM
RRRRRRRRRzRR)dqv.RR:Xv)qdc.X1RR
RRRRRRRRRRRRRbRRFRs0lRNb5R7d=#>R__HMs5CodR2,7=.R>_R#HsM_C.o527,R4>R=RH#_MC_so254,jR7RR=>#M_H_osC5,j2
SSSRRRRRRRRRRRRRjRqRR=>D_FINs885,j2RRq4=D>RFNI_858s4R2,q=.R>FRDI8_N8.s52R,
RRRRRRRRRRRRRRRRRRRRRRRRRRqd=D>RFNI_858sdR2,q=cR>FRDI8_N8cs52W,R >R=R0Is__CMdR.,WiBpRR=>B,piRS
SSSSSRdRmRR=>F_k0L_k#dM.5kOl_C_DDdd.,2m,R.>R=R0Fk_#Lk_5d.M_klODCD_,d..
2,SSSSSRSRm=4R>kRF0k_L#._d5lMk_DOCD._d,,42RRmj=F>RkL0_kd#_.k5MlC_ODdD_.2,j2R;
RRRRRRRRRRRRR#RR_0Fk_osC5Rd2<F=RkL0_kd#_.k5MlC_ODdD_.2,dRCIEMFR5kC0_M._dR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRR_R#F_k0s5Co.<2R=kRF0k_L#._d5lMk_DOCD._d,R.2IMECRk5F0M_C_Rd.=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRF#_ks0_C4o52=R<R0Fk_#Lk_5d.M_klODCD_,d.4I2RERCM50Fk__CMd=.RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRR#k_F0C_so25jRR<=F_k0L_k#dM.5kOl_C_DDdj.,2ERIC5MRF_k0CdM_.RR='24'R#CDCZR''R;
RRRRRCRRMo8RCsMCNR0Cz_.ccR;
RRRRRzRR.dc_RH:RVIR5HE80Rd=R2CRoMNCs0RC
RRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)Rzq.vdRD:RNDLCRRH#"a11"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloMC5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*n2RR&"RW"&MRH0CCosl'HN5oCj&2RR"" RH&RMo0CCHs'lCNo50oC_8CM_b8C0ME5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*nRd+R.8,RCEb02&2RR""XRH&RMo0CCHs'lCNo5;c2
RRRRRRRRRRRRoLCHRM
RRRRRRRRRzRR)dqv.RR:Xv)qdc.X1RR
RRRRRRRRRRRRRbRRFRs0lRNb5R7d='>RjR',7=.R>_R#HsM_C.o527,R4>R=RH#_MC_so254,jR7RR=>#M_H_osC5,j2
SSSRRRRRRRRRRRRRjRqRR=>D_FINs885,j2RRq4=D>RFNI_858s4R2,q=.R>FRDI8_N8.s52R,
RRRRRRRRRRRRRRRRRRRRRRRRRRqd=D>RFNI_858sdR2,q=cR>FRDI8_N8cs52W,R >R=R0Is__CMdR.,WiBpRR=>B,piRS
SSSSSRdRmRR=>FMbC,.RmRR=>F_k0L_k#dM.5kOl_C_DDd..,2S,
SSSSSmRR4>R=R0Fk_#Lk_5d.M_klODCD_,d.4R2,m=jR>kRF0k_L#._d5lMk_DOCD._d,2j2;R
RRRRRRRRRRRRRR_R#F_k0s5Co.<2R=kRF0k_L#._d5lMk_DOCD._d,R.2IMECRk5F0M_C_Rd.=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRF#_ks0_C4o52=R<R0Fk_#Lk_5d.M_klODCD_,d.4I2RERCM50Fk__CMd=.RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRR#k_F0C_so25jRR<=F_k0L_k#dM.5kOl_C_DDdj.,2ERIC5MRF_k0CdM_.RR='24'R#CDCZR''R;
RRRRRCRRMo8RCsMCNR0Cz_.cdS;
S8CMRMoCC0sNCORzEc	_;S
Sz	OE_:.RRRHV5I#_HE80_sNsN4$52RR>jo2RCsMCN
0CRRRRRRRRzR.c:FRVsRR[H5MR#H_I8_0ENNss$254R4-R2FR8IFM0RojRCsMCN
0CRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FzVR)dqv.RR:DCNLD#RHR1"1a&"RR0HMCsoC'NHloIC5HE802RR&"R7"&MRH0CCosl'HN5oCM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*c&2RR""WRH&RMo0CCHs'lCNo58IH0UE-*I#_HE80_sNsNd$52*-.[2-.R"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05lMk_DOCD._4U.*4URR+M_klODCD_*ncn+cRR,d.Rb8C02E2R"&RX&"RR0HMCsoC'NHloIC5HE80-#U*_8IH0NE_s$sN5-d2.2*[;R
RRRRRRRRRRCRLo
HMRRRRRRRRRRRRzv)qd:.RRv)qd..X1RR
RRRRRRRRRRRRRbRRFRs0lRNb5R7j=#>R__HMs5CoI0H8E*-U#H_I8_0ENNss$25d-[.*-,.2RR74=#>R__HMs5CoI0H8E*-U#H_I8_0ENNss$25d-[.*-,42RRqj=D>RFNI_858sjR2,q=4R>FRDI8_N84s52q,R.>R=RIDF_8N8s25.,R
RRRRRRRRRRRRRRRRRRRRRRRRRq=dR>FRDI8_N8ds52q,Rc>R=RIDF_8N8s25c, RWRR=>I_s0CdM_.W,RBRpi=B>RpRi,m=jR>kRF0k_L#._d5lMk_DOCD._d,8IH0UE-*I#_HE80_sNsNd$52*-.[2-.,S
SSSSSR4RmRR=>F_k0L_k#dM.5kOl_C_DDdI.,HE80-#U*_8IH0NE_s$sN5-d2.-*[4;22
RRRRRRRRRRRRRRRRF#_ks0_CIo5HE80-#U*_8IH0NE_s$sN5-d2.-*[4<2R=kRF0k_L#._d5lMk_DOCD._d,8IH0UE-*I#_HE80_sNsNd$52*-.[2-4RCIEMFR5kC0_M._dR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRR_R#F_k0s5CoI0H8E*-U#H_I8_0ENNss$25d-[.*-R.2<F=RkL0_kd#_.k5MlC_ODdD_.H,I8-0EU_*#I0H8Es_Ns5N$d.2-*.[-2ERIC5MRF_k0CdM_.RR='24'R#CDCZR''R;
RRRRRCRRMo8RCsMCNR0Cz;.c
CSSMo8RCsMCNR0Cz	OE_
.;SOSzE4	_RH:RV#R5_8IH0NE_s$sN5Rj2>2RjRMoCC0sNCR
RRRRRR.RzcRR:H5VRI0H8EFRl8RRU=2R4RMoCC0sNCR
RRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqz)vRd.:NRDLRCDH"#R1"1aRH&RMo0CCHs'lCNo58IH0RE2&7R""RR&HCM0o'CsHolNCk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*2ncR"&RW&"RR0HMCsoC'NHlojC52RR&"R "&MRH0CCosl'HN5oCo_C0C_M880CbEk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*Rnc+.Rd,CR8b20E2RR&"RX"&MRH0CCosl'HN5oC4
2;RRRRRRRRRRRRLHCoMR
RRRRRRRRRR)Rzq.vdR):Rq.vdXR41
RRRRRRRRRRRRRRRRsbF0NRlb7R5RR=>#M_H_osC5,j2RRqj=D>RFNI_858sjR2,q=4R>FRDI8_N84s52q,R.>R=RIDF_8N8s25.,R
RRRRRRRRRRRRRRRRRRRRRRRRRq=dR>FRDI8_N8ds52q,Rc>R=RIDF_8N8s25c, RWRR=>I_s0CdM_.W,RBRpi=B>RpRi,m>R=R0Fk_#Lk_5d.M_klODCD_,d.j;22
RRRRRRRRRRRRRRRRF#_ks0_Cjo52=R<R0Fk_#Lk_5d.M_klODCD_,d.jI2RERCM50Fk__CMd=.RR''42DRC#'CRZ
';RRRRRRRRCRM8oCCMsCN0Rcz.;S
SCRM8oCCMsCN0REzO	;_4
RRRR8CMRMoCC0sNC.Rz4R;RRRRRRRRR
R
RR-R-RMtCC0sNCRRN4InRFRs88bCCRv)qRDOCDVRHRbNbssFbHCN0RRRRRRRRRRRRR
RRRRRRzR.6:VRHRk5MlC_OD4D_nRR=4o2RCsMCN
0CRRRR-Q-RVNR58I8sHE80R6>R2CRMC08RFsROCCN0RHIs0CCRMDNLCMRN8kRF00bkRNCMLRDC#CCDOD0RFOoH
RRRRRRRRnz.NRR:H5VRNs88I0H8ERR>(MRN8kRMlC_ODnD_cRR=4MRN8kRMlC_ODdD_.RR=4o2RCsMCN
0CRRRRRRRRRRRRRRRRF_k0C4M_n=R<R''4RCIEM5R5#8_N_osC58N8s8IH04E-RI8FMR0F(=2RRlMk_DOCD._4UN2RM58R#8_N_osC5Rn2=4R''N2RM58R#8_N_osC5R62=4R''N2RM58R#8_N_osC5Rc2=jR''R22CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C_R4n<W=R ERIC5MR5N#_8C_so85N8HsI8-0E4FR8IFM0RR(2=kRMlC_OD4D_.RU2NRM85N#_8C_so25nR'=R4R'2NRM85N#_8C_so256R'=R4R'2NRM85N#_8C_so25cR'=Rj2'2R#CDCjR''R;
RRRRRCRRMo8RCsMCNR0CzN.n;R
RRRRRR.Rzn:LRRRHV58N8s8IH0>ERRN(RMM8RkOl_C_DDn=cRRN4RMM8RkOl_C_DDd=.RRRj2oCCMsCN0
RRRRRRRRRRRRRRRR0Fk__CM4<nR=4R''ERIC5MR5N#_8C_so85N8HsI8-0E4FR8IFM0RR(2=kRMlC_OD4D_.RU2NRM85N#_8C_so25nR'=R4R'2NRM85N#_8C_so256R'=RjR'2NRM85N#_8C_so25cR'=Rj2'2R#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_Mn_4RR<=WI RERCM5_5#Ns8_CNo58I8sHE80-84RF0IMF2R(RM=RkOl_C_DD42.UR8NMR_5#Ns8_Cno52RR='24'R8NMR_5#Ns8_C6o52RR='2j'R8NMR_5#Ns8_Cco52RR='2j'2DRC#'CRj
';RRRRRRRRCRM8oCCMsCN0Rnz.LR;
RRRRRzRR.RnO:VRHR85N8HsI8R0E>RR(NRM8M_klODCD_Rnc=RRjNRM8M_klODCD_Rd.=2R4RMoCC0sNCR
RRRRRRRRRRRRRRkRF0M_C_R4n<'=R4I'RERCM5_5#Ns8_CNo58I8sHE80-84RF0IMF2R(RM=RkOl_C_DD42.UR8NMR_5#Ns8_Cno52RR='2j'R8NMR_5#Ns8_C6o52RR='24'R8NMR_5#Ns8_Cco52RR='2j'2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0C4M_n=R<RRW IMECR#55__N8s5CoNs88I0H8ER-48MFI0(FR2RR=M_klODCD_U4.2MRN8#R5__N8s5Con=2RR''j2MRN8#R5__N8s5Co6=2RR''42MRN8#R5__N8s5Coc=2RR''j2C2RDR#C';j'
RRRRRRRR8CMRMoCC0sNC.Rzn
O;RRRRRRRRz8.nRH:RVNR58I8sHE80R(>RR8NMRlMk_DOCDc_nRj=RR8NMRlMk_DOCD._dRj=R2CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_Mn_4RR<='R4'IMECR#55__N8s5CoNs88I0H8ER-48MFI0(FR2RR=M_klODCD_U4.2MRN8#R5__N8s5Con=2RR''j2MRN8#R5__N8s5Co6=2RR''j2MRN8#R5__N8s5Coc=2RR''j2C2RDR#C';j'
RRRRRRRRRRRRRRRR0Is__CM4<nR= RWRCIEM5R5#8_N_osC58N8s8IH04E-RI8FMR0F(=2RRlMk_DOCD._4UN2RM58R#8_N_osC5Rn2=jR''N2RM58R#8_N_osC5R62=jR''N2RM58R#8_N_osC5Rc2=jR''R22CCD#R''j;R
RRRRRRMRC8CRoMNCs0zCR.;n8
RRRRRRRRnz.CRR:H5VRNs88I0H8ERR=(MRN8kRMlC_ODnD_cRR=4MRN8kRMlC_ODdD_.RR=4o2RCsMCN
0CRRRRRRRRRRRRRRRRF_k0C4M_n=R<R''4RCIEM5R5#8_N_osC5Rn2=4R''N2RM58R#8_N_osC5R62=4R''N2RM58R#8_N_osC5Rc2=jR''R22CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C_R4n<W=R ERIC5MR5N#_8C_so25nR'=R4R'2NRM85N#_8C_so256R'=R4R'2NRM8R_5#Ns8_Cco52RR='2j'2DRC#'CRj
';RRRRRRRRCRM8oCCMsCN0Rnz.CR;
RRRRRzRR.RnV:VRHR85N8HsI8R0E=RR(NRM8M_klODCD_Rnc=RR4NRM8M_klODCD_Rd.=2RjRMoCC0sNCR
RRRRRRRRRRRRRRkRF0M_C_R4n<'=R4I'RERCM5_5#Ns8_Cno52RR='24'R8NMR_5#Ns8_C6o52RR='2j'R8NMR_5#Ns8_Cco52RR='2j'2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0C4M_n=R<RRW IMECR#55__N8s5Con=2RR''42MRN8#R5__N8s5Co6=2RR''j2MRN8#R5__N8s5Coc=2RR''j2C2RDR#C';j'
RRRRRRRR8CMRMoCC0sNC.Rzn
V;RRRRRRRRzo.nRH:RVNR58I8sHE80Rn=RR8NMRlMk_DOCDc_nRj=RR8NMRlMk_DOCD._dR4=R2CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_Mn_4RR<='R4'IMECR#55__N8s5Co6=2RR''42MRN8#R5__N8s5Coc=2RR''j2C2RDR#C';j'
RRRRRRRRRRRRRRRR0Is__CM4<nR= RWRCIEM5R5#8_N_osC5R62=4R''N2RM58R#8_N_osC5Rc2=jR''R22CCD#R''j;R
RRRRRRMRC8CRoMNCs0zCR.;no
RRRRRRRRnz.ERR:H5VRNs88I0H8ERR=6MRN8kRMlC_ODdD_.=R/RR42oCCMsCN0
RRRRRRRRRRRRRRRR0Fk__CM4<nR=4R''ERIC5MR5N#_8C_so85N8HsI8-0E4FR8IFM0RRc2=kRMlC_ODdD_.R22CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C_R4n<W=R ERIC5MR5N#_8C_so85N8HsI8-0E4FR8IFM0RRc2=kRMlC_ODdD_.R22CCD#R''j;R
RRRRRRMRC8CRoMNCs0zCR.;nE
RRRRR--Q5VRNs88I0H8E=R<RR62MIFRsCH0RNCMLRDCFFsRkk0b0MRCNCLDRD#CCRO0DHFoOCRMC88C
RRRRRRRR(z.RH:RVNR58I8sHE80RR<=co2RCsMCN
0CRRRRRRRRRRRRRRRRF_k0C4M_n=R<R''4;R
RRRRRRRRRRRRRRsRI0M_C_R4n<W=R R;
RRRRRCRRMo8RCsMCNR0Cz;.(
RRRRR--tCCMsCN0RC0ERv)qRDOCDMRN8sR0H0-#N
0CSRRRREzO	R_U:VRHR_5#I0H8Es_Ns5N$d>2RRRj2oCCMsCN0
zSSO_E	DRC6:VRHRH5I8R0E>U=R*I#_HE80_sNsNd$52MRN8HRI8R0E>U=R2CRoMNCs0RC
RRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)Rzqnv4RD:RNDLCRRH#"a11"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloMC5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*nRM+RkOl_C_DDdd.*.&2RR""WRH&RMo0CCHs'lCNo58IH0-ERRLD#_8IH0RE2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50EM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*cRR+M_klODCD_*d.d+.RR,4nRb8C02E2R"&RX&"RR0HMCsoC'NHloIC5HE80RD-R#IL_HE80RU+R2R;
RRRRRRRRRLRRCMoH
RSSRzRR)4qvnRR:Xv)q4UnX1S
SSRRRRsbF0NRlb7R5RR=>b5N8#M_H_osC58IH04E-RI8FMR0FI0H8E#-DLH_I820E,,RURLD#_8IH04E-2q,Rj>R=RIDF_8N8s25j,S
SSSSSR4RqRR=>D_FINs885,42RRq.=D>RFNI_858s.R2,q=dR>FRDI8_N8ds52W,R >R=R0Is__CM4Rn,WiBpRR=>B,pi
SSSSRSSR=mR>lR0b__U4jn52
2;SSSSNH##o:MRRsVFRRH[HIMRHE80-84RF0IMFHRI8-0ED_#LI0H8ECRoMNCs0SC
SRSSR0Fk_#Lk_54nM_klODCD_,4nHR[2<0=RlUb__54njH25[H-I8+0ED_#LI0H8E
2;RRRRRRRRRRRRRRRRR_R#F_k0s5CoHR[2<F=RkL0_k4#_nk5MlC_OD4D_n[,H2ERIC5MRF_k0C4M_nRR='24'R#CDCZR''S;
SCSSMo8RCsMCNR0CNH##o
M;RRRRRRRRRRRRzR.U:FRVsRR[H#MR_8IH0NE_s$sN5-d24FR8IFM0Ro4RCsMCN
0CRRRRRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqz)vR4n:NRDLRCDH"#R1"1aRH&RMo0CCHs'lCNo58IH0RE2&7R""RR&HCM0o'CsHolNCk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*Rnc+kRMlC_ODdD_..*d2RR&"RW"&MRH0CCosl'HN5oCI0H8ERR-D_#LI0H8ERR-[2*UR"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05lMk_DOCD._4U.*4URR+M_klODCD_*ncn+cRRlMk_DOCD._d*Rd.+nR4,CR8b20E2RR&"RX"&MRH0CCosl'HN5oCI0H8ERR-D_#LI0H8ERR-54[-22*U;R
RRRRRRRRRRRRRLHCoMR
RRRRRRRRRRRRRzv)q4:nRRqX)vX4nU
1RRRRRRRRRRRRRRRRRb0FsRblNRR57=#>R__HMs5CoI0H8E#-DLH_I8-0EU+*[(FR8IFM0R8IH0DE-#IL_HE80-[U*2q,Rj>R=RIDF_8N8s25j,4RqRR=>D_FINs885,42RRq.=D>RFNI_858s.
2,RRRRRRRRRRRRRRRRRRRRRRRRRdRqRR=>D_FINs885,d2RRW =I>RsC0_Mn_4,BRWp=iR>pRBim,RRR=>0_lbUn_452[2;S
SSRRRR#N#HRoM:FRVs[RHRRHM(FR8IFM0RojRCsMCN
0CSSSSRkRF0k_L#n_45lMk_DOCDn_4,8IH0DE-#IL_HE80-[U*+2H[RR<=0_lbUn_455[2H;[2
RRRRRRRRRRRRRRRR#RR_0Fk_osC58IH0DE-#IL_HE80-[U*+2H[RR<=F_k0L_k#4Mn5kOl_C_DD4In,HE80-LD#_8IH0UE-*H[+[I2RERCM50Fk__CM4=nRR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRCRM8oCCMsCN0R#N#H;oM
RRRRRRRRRRRR8CMRMoCC0sNC.RzUS;
S8CMRMoCC0sNCORzED	_C
6;SOSzEo	_0:6RRRHV58IH0>ER=RRUNRM8I0H8EFRl8RRU>6=R2CRoMNCs0RC
RRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)Rzqnv4RD:RNDLCRRH#"a11"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloMC5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*nRM+RkOl_C_DDdd.*.&2RR""WRH&RMo0CCHs'lCNo58IH0-ERRLD#_8IH0RE2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50EM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*cRR+M_klODCD_*d.d+.RR,4nRb8C02E2R"&RX&"RR0HMCsoC'NHloIC5HE80RD-R#IL_HE80RU+R2R;
RRRRRRRRRLRRCMoH
RSSRzRR)4qvnRR:Xv)q4UnX1S
SSRRRRsbF0NRlb7R5RR=>b5N8#M_H_osC58IH04E-RI8FMR0FI0H8E#-DLH_I820E,,RURLD#_8IH04E-2q,Rj>R=RIDF_8N8s25j,S
SSSSSR4RqRR=>D_FINs885,42RRq.=D>RFNI_858s.R2,q=dR>FRDI8_N8ds52W,R >R=R0Is__CM4Rn,WiBpRR=>B,pi
SSSSRSSR=mR>lR0b__U4#n5_8IH0NE_s$sN5-d24;22
SSSS#N#HRoM:FRVs[RHRRHMI0H8ER-48MFI0IFRHE80-LD#_8IH0oERCsMCN
0CSSSSRkRF0k_L#n_45lMk_DOCDn_4,2H[RR<=0_lbUn_45I#_HE80_sNsNd$522-45-H[I0H8E#+DLH_I820E;R
RRRRRRRRRRRRRRRRR#k_F0C_so[5H2=R<R0Fk_#Lk_54nM_klODCD_,4nHR[2IMECRk5F0M_C_R4n=4R''C2RDR#C';Z'
SSSS8CMRMoCC0sNC#RN#MHo;R
RRRRRRRRRR.RzURR:VRFs[MRHRI#_HE80_sNsNd$52R-.8MFI0jFRRMoCC0sNCR
RRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FzVR)4qvnRR:DCNLD#RHR1"1a&"RR0HMCsoC'NHloIC5HE802RR&"R7"&MRH0CCosl'HN5oCM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*cRR+M_klODCD_*d.dR.2&WR""RR&HCM0o'CsHolNC*5[U&2RR"" RH&RMo0CCHs'lCNo50oC_8CM_b8C0ME5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*nRM+RkOl_C_DDdd.*.RR+4Rn,80CbER22&XR""RR&HCM0o'CsHolNC[55+*42U
2;RRRRRRRRRRRRRCRLo
HMRRRRRRRRRRRRR)Rzqnv4RX:R)4qvn1XURR
RRRRRRRRRRRRRRFRbsl0RN5bR7>R=RH#_MC_so*5U[R+(8MFI0UFR*,[2RRqj=D>RFNI_858sjR2,q=4R>FRDI8_N84s52q,R.>R=RIDF_8N8s25.,R
RRRRRRRRRRRRRRRRRRRRRRRRRq=dR>FRDI8_N8ds52W,R >R=R0Is__CM4Rn,WiBpRR=>B,piR=mR>lR0b__U4[n52
2;SSSSNH##o:MRRsVFRRH[H(MRRI8FMR0FjCRoMNCs0SC
SRSSR0Fk_#Lk_54nM_klODCD_,4nU+*[HR[2<0=RlUb__54n[H25[
2;RRRRRRRRRRRRRRRRR_R#F_k0s5CoU+*[HR[2<F=RkL0_k4#_nk5MlC_OD4D_n*,U[[+H2ERIC5MRF_k0C4M_nRR='24'R#CDCZR''R;
RRRRRRRRRRRRRCRRMo8RCsMCNR0CNH##o
M;RRRRRRRRRRRRCRM8oCCMsCN0RUz.;S
SCRM8oCCMsCN0REzO	0_o6S;
SEzO	R_M:VRHRH5I8R0E<2RURMoCC0sNCR
RRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqz)vR4n:NRDLRCDH"#R1"1aRH&RMo0CCHs'lCNo58IH0RE2&7R""RR&HCM0o'CsHolNCk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*Rnc+kRMlC_ODdD_..*d2RR&"RW"&MRH0CCosl'HN5oCj&2RR"" RH&RMo0CCHs'lCNo50oC_8CM_b8C0ME5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*nRM+RkOl_C_DDdd.*.RR+4Rn,80CbER22&XR""RR&HCM0o'CsHolNC25U;R
RRRRRRRRRRCRLo
HMSRSRR)Rzqnv4RX:R)4qvn1XU
SSSRRRRb0FsRblNRR57=b>RN#85__HMs5CoI0H8ER-48MFI0IFRHE80-LD#_8IH0,E2RRU,D_#LI0H8E2-4,jRqRR=>D_FINs885,j2
SSSSRSSRRq4=D>RFNI_858s4R2,q=.R>FRDI8_N8.s52q,Rd>R=RIDF_8N8s25d, RWRR=>I_s0C4M_nW,RBRpi=B>Rp
i,SSSSSRSRm>R=Rb0l_4U_n25j2S;
SNSS#o#HMRR:VRFsHH[RMHRI8-0E4FR8IFM0RojRCsMCN
0CSSSSRkRF0k_L#n_45lMk_DOCDn_4,2H[RR<=0_lbUn_455j2H;[2
RRRRRRRRRRRRRRRR#RR_0Fk_osC52H[RR<=F_k0L_k#4Mn5kOl_C_DD4Hn,[I2RERCM50Fk__CM4=nRR''42DRC#'CRZ
';SSSSCRM8oCCMsCN0R#N#H;oM
CSSMo8RCsMCNR0Cz	OE_
M;SMSC8CRoMNCs0zCRO_E	US;
SEzO	R_c:VRHR_5#I0H8Es_Ns5N$.>2RRRj2oCCMsCN0
RRRRRRRRgz._:cRRRHV58IH0>ER=2RcRMoCC0sNCR
RRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqz)vR4n:NRDLRCDH"#R1"1aRH&RMo0CCHs'lCNo58IH0RE2&7R""RR&HCM0o'CsHolNCk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*Rnc+kRMlC_ODdD_..*d2RR&"RW"&MRH0CCosl'HN5oCj&2RR"" RH&RMo0CCHs'lCNo50oC_8CM_b8C0ME5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*nRM+RkOl_C_DDdd.*.RR+4Rn,80CbER22&XR""RR&HCM0o'CsHolNC25c;R
RRRRRRRRRRCRLo
HMRRRRRRRRRRRRzv)q4:nRRv)q4cnX1RR
RRRRRRRRRRRRRbRRFRs0lRNb5R7d=#>R__HMs5CodR2,7=.R>_R#HsM_C.o527,R4>R=RH#_MC_so254,jR7RR=>#M_H_osC5,j2
SSSRRRRRRRRRRRRRjRqRR=>D_FINs885,j2RRq4=D>RFNI_858s4R2,q=.R>FRDI8_N8.s52R,
RRRRRRRRRRRRRRRRRRRRRRRRRRqd=D>RFNI_858sdR2,W= R>sRI0M_C_,4nRpWBi>R=RiBp,SR
SSSSSmRRd>R=R0Fk_#Lk_54nM_klODCD_,4ndR2,m=.R>kRF0k_L#n_45lMk_DOCDn_4,,.2
SSSSRSSRRm4=F>RkL0_k4#_nk5MlC_OD4D_n2,4,jRmRR=>F_k0L_k#4Mn5kOl_C_DD4jn,2
2;RRRRRRRRRRRRRRRR#k_F0C_so25dRR<=F_k0L_k#4Mn5kOl_C_DD4dn,2ERIC5MRF_k0C4M_nRR='24'R#CDCZR''R;
RRRRRRRRRRRRR#RR_0Fk_osC5R.2<F=RkL0_k4#_nk5MlC_OD4D_n2,.RCIEMFR5kC0_Mn_4R'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRR_R#F_k0s5Co4<2R=kRF0k_L#n_45lMk_DOCDn_4,R42IMECRk5F0M_C_R4n=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRF#_ks0_Cjo52=R<R0Fk_#Lk_54nM_klODCD_,4njI2RERCM50Fk__CM4=nRR''42DRC#'CRZ
';RRRRRRRRCRM8oCCMsCN0Rgz._
c;RRRRRRRRz_.gdRR:H5VRI0H8ERR=do2RCsMCN
0CRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FzVR)4qvnRR:DCNLD#RHR1"1a&"RR0HMCsoC'NHloIC5HE802RR&"R7"&MRH0CCosl'HN5oCM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*cRR+M_klODCD_*d.dR.2&WR""RR&HCM0o'CsHolNC25jR"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05lMk_DOCD._4U.*4URR+M_klODCD_*ncn+cRRlMk_DOCD._d*Rd.+nR4,CR8b20E2RR&"RX"&MRH0CCosl'HN5oCc
2;RRRRRRRRRRRRLHCoMR
RRRRRRRRRR)Rzqnv4R):Rqnv4XRc1
RRRRRRRRRRRRRRRRsbF0NRlb7R5d>R=R''j,.R7RR=>#M_H_osC5,.2RR74=#>R__HMs5Co4R2,7=jR>_R#HsM_Cjo52S,
SRSRRRRRRRRRRRRRq=jR>FRDI8_N8js52q,R4>R=RIDF_8N8s254,.RqRR=>D_FINs885,.2
RRRRRRRRRRRRRRRRRRRRRRRRqRRd>R=RIDF_8N8s25d, RWRR=>I_s0C4M_nW,RBRpi=B>RpRi,
SSSSRSSRRmd=F>Rb,CMRRm.=F>RkL0_k4#_nk5MlC_OD4D_n2,.,S
SSSSSR4RmRR=>F_k0L_k#4Mn5kOl_C_DD44n,2m,Rj>R=R0Fk_#Lk_54nM_klODCD_,4nj;22
RRRRRRRRRRRRRRRRF#_ks0_C.o52=R<R0Fk_#Lk_54nM_klODCD_,4n.I2RERCM50Fk__CM4=nRR''42DRC#'CRZ
';RRRRRRRRRRRRRRRR#k_F0C_so254RR<=F_k0L_k#4Mn5kOl_C_DD44n,2ERIC5MRF_k0C4M_nRR='24'R#CDCZR''R;
RRRRRRRRRRRRR#RR_0Fk_osC5Rj2<F=RkL0_k4#_nk5MlC_OD4D_n2,jRCIEMFR5kC0_Mn_4R'=R4R'2CCD#R''Z;R
RRRRRRMRC8CRoMNCs0zCR.dg_;S
SCRM8oCCMsCN0REzO	;_c
zSSO_E	.RR:H5VR#H_I8_0ENNss$254Rj>R2CRoMNCs0RC
RRRRRzRRd:jRRsVFRH[RM#R5_8IH0NE_s$sN5R42-2R4RI8FMR0FjCRoMNCs0RC
RRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)Rzqnv4RD:RNDLCRRH#"a11"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloMC5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*nRM+RkOl_C_DDdd.*.&2RR""WRH&RMo0CCHs'lCNo58IH0UE-*I#_HE80_sNsNd$52*-.[2-.R"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05lMk_DOCD._4U.*4URR+M_klODCD_*ncn+cRRlMk_DOCD._d*Rd.+nR4,CR8b20E2RR&"RX"&MRH0CCosl'HN5oCI0H8E*-U#H_I8_0ENNss$25d-[.*2R;
RRRRRRRRRLRRCMoH
RRRRRRRRRRRRqz)vR4n:qR)vX4n.
1RRRRRRRRRRRRRRRRRb0FsRblNRj57RR=>#M_H_osC58IH0UE-*I#_HE80_sNsNd$52*-.[2-.,4R7RR=>#M_H_osC58IH0UE-*I#_HE80_sNsNd$52*-.[2-4,jRqRR=>D_FINs885,j2RRq4=D>RFNI_858s4R2,q=.R>FRDI8_N8.s52R,
RRRRRRRRRRRRRRRRRRRRRRRRRRqd=D>RFNI_858sdR2,W= R>sRI0M_C_,4nRpWBi>R=RiBp,jRmRR=>F_k0L_k#4Mn5kOl_C_DD4In,HE80-#U*_8IH0NE_s$sN5-d2.-*[.
2,SSSSSRSRm=4R>kRF0k_L#n_45lMk_DOCDn_4,8IH0UE-*I#_HE80_sNsNd$52*-.[2-42R;
RRRRRRRRRRRRR#RR_0Fk_osC58IH0UE-*I#_HE80_sNsNd$52*-.[2-4RR<=F_k0L_k#4Mn5kOl_C_DD4In,HE80-#U*_8IH0NE_s$sN5-d2.-*[4I2RERCM50Fk__CM4=nRR''42DRC#'CRZ
';RRRRRRRRRRRRRRRR#k_F0C_soH5I8-0EU_*#I0H8Es_Ns5N$d.2-*.[-2=R<R0Fk_#Lk_54nM_klODCD_,4nI0H8E*-U#H_I8_0ENNss$25d-[.*-R.2IMECRk5F0M_C_R4n=4R''C2RDR#C';Z'
RRRRRRRR8CMRMoCC0sNCdRzjS;
S8CMRMoCC0sNCORzE.	_;S
Sz	OE_:4RRRHV5I#_HE80_sNsNj$52RR>jo2RCsMCN
0CRRRRRRRRzRd4:VRHRH5I8R0ElRF8URR=4o2RCsMCN
0CRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FzVR)4qvnRR:DCNLD#RHR1"1a&"RR0HMCsoC'NHloIC5HE802RR&"R7"&MRH0CCosl'HN5oCM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*cRR+M_klODCD_*d.dR.2&WR""RR&HCM0o'CsHolNC25jR"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05lMk_DOCD._4U.*4URR+M_klODCD_*ncn+cRRlMk_DOCD._d*Rd.+nR4,CR8b20E2RR&"RX"&MRH0CCosl'HN5oC4
2;RRRRRRRRRRRRLHCoMR
RRRRRRRRRR)Rzqnv4R):Rqnv4XR41
RRRRRRRRRRRRRRRRsbF0NRlb7R5RR=>#M_H_osC5,j2RRqj=D>RFNI_858sjR2,q=4R>FRDI8_N84s52q,R.>R=RIDF_8N8s25.,R
RRRRRRRRRRRRRRRRRRRRRRRRRq=dR>FRDI8_N8ds52W,R >R=R0Is__CM4Rn,WiBpRR=>B,piR=mR>kRF0k_L#n_45lMk_DOCDn_4,2j2;R
RRRRRRRRRRRRRR_R#F_k0s5Coj<2R=kRF0k_L#n_45lMk_DOCDn_4,Rj2IMECRk5F0M_C_R4n=4R''C2RDR#C';Z'
RRRRRRRR8CMRMoCC0sNCdRz4S;
S8CMRMoCC0sNCORzE4	_;R
RRCRRMo8RCsMCNR0Cz;.6RRRRRRRRRRR
RMRC8CRoMNCs0zCRc
c;CRM8NEsOHO0C0CksRFLDOs	_N
l;
ONsECH0Os0kCFRM__sIOOEC	VRFRv)q_R)WHO#
FFlbM0CMRqX)vU4.X
41RsbF0
R5RmRRRF:Rk#0R0D8_FOoH;R
RRRqj:MRHR8#0_oDFH
O;RqRR4RR:H#MR0D8_FOoH;R
RRRq.:MRHR8#0_oDFH
O;RqRRdRR:H#MR0D8_FOoH;R
RRRqc:MRHR8#0_oDFH
O;RqRR6RR:H#MR0D8_FOoH;R
RRRqn:MRHR8#0_oDFH
O;R7RRRH:RM0R#8F_Do;HO
RRRWiBpRH:RM0R#8F_Do;HO
RRRW: RRRHM#_08DHFoO2
R;M
C8FROlMbFC;M0
O

FFlbM0CMRqX)vXnc.R1
b0FsRR5
RjRmRF:Rk#0R0D8_FOoH;R
RRRm4:kRF00R#8F_Do;HO
RRRq:jRRRHM#_08DHFoOR;
R4RqRH:RM0R#8F_Do;HO
RRRq:.RRRHM#_08DHFoOR;
RdRqRH:RM0R#8F_Do;HO
RRRq:cRRRHM#_08DHFoOR;
R6RqRH:RM0R#8F_Do;HO
RRR7:jRRRHM#_08DHFoOR;
R4R7RH:RM0R#8F_Do;HO
RRRWiBpRH:RM0R#8F_Do;HO
RRRW: RRRHM#_08DHFoO2
R;M
C8FROlMbFC;M0
F
OlMbFCRM0Xv)qdc.X1b
RFRs05R
RRRmj:kRF00R#8F_Do;HO
RRRm:4RR0FkR8#0_oDFH
O;RmRR.RR:FRk0#_08DHFoOR;
RdRmRF:Rk#0R0D8_FOoH;R
RRRqj:MRHR8#0_oDFH
O;RqRR4RR:H#MR0D8_FOoH;R
RRRq.:MRHR8#0_oDFH
O;RqRRdRR:H#MR0D8_FOoH;R
RRRqc:MRHR8#0_oDFH
O;R7RRjRR:H#MR0D8_FOoH;R
RRR74:MRHR8#0_oDFH
O;R7RR.RR:H#MR0D8_FOoH;R
RRR7d:MRHR8#0_oDFH
O;RWRRBRpi:MRHR8#0_oDFH
O;RWRR RR:H#MR0D8_FOoH
;R2
8CMRlOFbCFMM
0;ObFlFMMC0)RXq.vdX
U1
FRbs50R
RRRmRR:FRk0#_08DHFoOC_POs0F58(RF0IMF2Rj;R
RRRqj:MRHR8#0_oDFH
O;RqRR4RR:H#MR0D8_FOoH;R
RRRq.:MRHR8#0_oDFH
O;RqRRdRR:H#MR0D8_FOoH;R
RRRqc:MRHR8#0_oDFH
O;R7RRRH:RM0R#8F_Do_HOP0COF(s5RI8FMR0Fj
2;RWRRBRpi:MRHR8#0_oDFH
O;RWRR RR:H#MR0D8_FOoH
;R2
8CMRlOFbCFMM
0;
lOFbCFMMX0R)4qvn1XU
FRbs50R
RRRmRR:FRk0#_08DHFoOC_POs0F58(RF0IMF2Rj;R
RRRqj:MRHR8#0_oDFH
O;RqRR4RR:H#MR0D8_FOoH;R
RRRq.:MRHR8#0_oDFH
O;RqRRdRR:H#MR0D8_FOoH;R
RR:7RRRHM#_08DHFoOC_POs0F58(RF0IMF2Rj;R
RRpWBiRR:H#MR0D8_FOoH;R
RRRW :MRHR8#0_oDFHRO
2C;
MO8RFFlbM0CM;k
VMHO0FVMRk_MOH0MH5:LRRFLFDMCN2CRs0MksRs#0HRMoHL#
CMoH
HRRVLR52ER0CRM
RsRRCs0kMh5"FCRsNI8/sCH0RMOFVODH0EROC3O	Rl1Hk0DNHRFMllH#NE0OR#bF#DHLC!R!"
2;RDRC#RC
RsRRCs0kMB5"F8kDR0MFRbHlDCClMA0RD	FORv)q3#RQRC0ERNsC88RN8#sC#CRso0H#C8sCRHk#M0oRE#CRNRlCOODF	#RNRC0ERv)q?;"2
CRRMH8RVC;
MV8Rk_MOH0MH;k
VMHO0FoMRCC0_M88_CEb05x#HCRR:HCM0oRCs;CR8bR0E:MRH0CCoss2RCs0kMMRH0CCos#RH
sPNHDNLCHRlMH_#x:CRR0HMCsoCRR:=jL;
CMoH
lRRH#M_HRxC:8=RCEb0;R
RH5VR#CHxR8<RCEb02ER0CRM
RlRRH#M_HRxC:#=RH;xC
CRRMH8RVR;
R0sCkRsMl_HM#CHx;M
C8CRo0M_C8C_8b;0E
0N0skHL0oCRCsMCNs0F_bsCFRs0:0R#soHM;0
N0LsHkR0CoCCMsFN0sC_sb0FsRRFVMsF_IE_OCRO	:sRNO0EHCkO0sHCR#kRVMHO_M5H0Ns88_osC2-;
-CRLoRHMLODF	NRsllRHblDCCNM00MHFRo#HM#ND
b0$CMRH0s_NsRN$HN#Rs$sNRR5j06FR2VRFR0HMCsoC;F
OMN#0MI0RHE80_sNsN:$RR0HM_sNsN:$R=4R5,,R.RRc,g4,RUd,Rn
2;O#FM00NMRb8C0NE_s$sNRH:RMN0_s$sNRR:=5d4nURc,U.4g,jRcgRn,.Ujc,jR4.Rc,624.;F
OMN#0M80RH.PdRH:RMo0CC:sR=IR5HE80-/42d
n;O#FM00NMRP8H4:nRR0HMCsoCRR:=58IH04E-2U/4;F
OMN#0M80RHRPU:MRH0CCos=R:RH5I8-0E4g2/;F
OMN#0M80RHRPc:MRH0CCos=R:RH5I8-0E4c2/;F
OMN#0M80RHRP.:MRH0CCos=R:RH5I8-0E4.2/;F
OMN#0M80RHRP4:MRH0CCos=R:RH5I8-0E442/;O

F0M#NRM0LDFF4RR:LDFFCRNM:5=R84HPRj>R2O;
F0M#NRM0LDFF.RR:LDFFCRNM:5=R8.HPRj>R2O;
F0M#NRM0LDFFcRR:LDFFCRNM:5=R8cHPRj>R2O;
F0M#NRM0LDFFURR:LDFFCRNM:5=R8UHPRj>R2O;
F0M#NRM0LDFF4:nRRFLFDMCNRR:=5P8H4>nRR;j2
MOF#M0N0FRLF.DdRL:RFCFDN:MR=8R5H.PdRj>R2
;
O#FM00NMRP8H4UndcRR:HCM0oRCs:5=R80CbE2-4/d4nU
c;O#FM00NMRP8HU.4gRH:RMo0CC:sR=8R5CEb0-/42U.4g;F
OMN#0M80RHjPcg:nRR0HMCsoCRR:=5b8C04E-2j/cg
n;O#FM00NMRP8H.UjcRH:RMo0CC:sR=8R5CEb0-/42.Ujc;F
OMN#0M80RHjP4.:cRR0HMCsoCRR:=5b8C04E-2j/4.
c;O#FM00NMRP8H6R4.:MRH0CCos=R:RC58b-0E462/4
.;
MOF#M0N0FRLF4D6.RR:LDFFCRNM:5=R86HP4>.RR;j2
MOF#M0N0FRLFjD4.:cRRFLFDMCNRR:=5P8H4cj.Rj>R2O;
F0M#NRM0LDFF.UjcRL:RFCFDN:MR=8R5HjP.c>URR;j2
MOF#M0N0FRLFjDcg:nRRFLFDMCNRR:=5P8HcnjgRj>R2O;
F0M#NRM0LDFFU.4gRL:RFCFDN:MR=8R5H4PUg>.RR;j2
MOF#M0N0FRLFnD4dRUc:FRLFNDCM=R:RH58Pd4nU>cRR;j2
F
OMN#0M#0RkIl_HE80RH:RMo0CC:sR=mRAmqp hF'b#F5LF2D4RA+Rm mpqbh'FL#5F.FD2RR+Apmm 'qhb5F#LDFFc+2RRmAmph q'#bF5FLFDRU2+mRAmqp hF'b#F5LFnD42O;
F0M#NRM0#_kl80CbERR:HCM0oRCs:6=RR5-RApmm 'qhb5F#LDFF624.RA+Rm mpqbh'FL#5F4FDj2.cRA+Rm mpqbh'FL#5F.FDj2cURA+Rm mpqbh'FL#5FcFDj2gnRA+Rm mpqbh'FL#5FUFD42g.2
;
O#FM00NMROI_EOFHCH_I8R0E:MRH0CCos=R:R8IH0NE_s$sN5l#k_8IH0;E2
MOF#M0N0_RIOHEFO8C_CEb0RH:RMo0CC:sR=CR8b_0ENNss$k5#lH_I820E;F
OMN#0M80R_FOEH_OCI0H8ERR:HCM0oRCs:I=RHE80_sNsN#$5k8l_CEb02O;
F0M#NRM08E_OFCHO_b8C0:ERR0HMCsoCRR:=80CbEs_Ns5N$#_kl80CbE
2;
MOF#M0N0_RII0H8Ek_MlC_ODRD#:MRH0CCos=R:RH5I8-0E4I2/_FOEH_OCI0H8ERR+4O;
F0M#NRM0IC_8b_0EM_klODCD#RR:HCM0oRCs:5=R80CbE2-4/OI_EOFHCC_8bR0E+;R4
F
OMN#0M80R_8IH0ME_kOl_C#DDRH:RMo0CC:sR=IR5HE80-/428E_OFCHO_8IH0+ERR
4;O#FM00NMR88_CEb0_lMk_DOCD:#RR0HMCsoCRR:=5b8C04E-2_/8OHEFO8C_CEb0R4+R;O

F0M#NRM0IH_#x:CRR0HMCsoCRR:=IH_I8_0EM_klODCD#RR*IC_8b_0EM_klODCD#O;
F0M#NRM08H_#x:CRR0HMCsoCRR:=8H_I8_0EM_klODCD#RR*8C_8b_0EM_klODCD#
;
O#FM00NMRFLFDR_8:FRLFNDCM=R:R_58#CHxRI-R_x#HC=R<R;j2
MOF#M0N0FRLFID_RL:RFCFDN:MR=FRM0F5LF8D_2
;
O#FM00NMRFOEH_OCI0H8ERR:HCM0oRCs:5=RApmm 'qhb5F#LDFF_R82*_R8OHEFOIC_HE802RR+5mAmph q'#bF5FLFD2_IRI*R_FOEH_OCI0H8E
2;O#FM00NMRFOEH_OC80CbERR:HCM0oRCs:5=RApmm 'qhb5F#LDFF_R82*_R8OHEFO8C_CEb02RR+5mAmph q'#bF5FLFD2_IRI*R_FOEH_OC80CbE
2;O#FM00NMR8IH0ME_kOl_C#DDRH:RMo0CC:sR=AR5m mpqbh'FL#5F_FD8*2R58IH04E-2_/8OHEFOIC_HE802RR+5mAmph q'#bF5FLFD2_IR5*RI0H8E2-4/OI_EOFHCH_I820ER4+R;F
OMN#0M80RCEb0_lMk_DOCD:#RR0HMCsoCRR:=5mAmph q'#bF5FLFD2_8R8*5CEb0-/428E_OFCHO_b8C0RE2+AR5m mpqbh'FL#5F_FDI*2RRC58b-0E4I2/_FOEH_OC80CbE+2RR
4;-F-OMN#0MM0RkOl_C#DDRH:RMo0CC:sR=5R55b8C0-ERRR42/.Rd2RR+5855CEb0R4-R2FRl8.Rd2RR/42n2;RRR-y-RRRFV)dqv.1X4RDOCDM#RCCC88-R
-MOF#M0N0CRDVF0_PRCs:MRH0CCos=R:R55580CbERR+4R62lRF8dR.2/nR42R;RRRRRRRRRRRRRRRRRRRRRR-RR-RRyF)VRqnv4XR41M8CCCV8RFDsRCRV0FsPCRsIF80#
$RbCF_k0L4k#_b0$C#RHRsNsN5$R80CbEk_MlC_OD-D#4FR8IFM0RRj,I0H8Ek_MlC_OD-D#4FR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNR0Fk_#Lk4RR:F_k0L4k#_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFR8s_FRk05bHMk00RFsR0H0-#N#0C2$
0bFCRkL0_k_#.0C$bRRH#NNss$8R5CEb0_lMk_DOCD4#-RI8FMR0Fj.,R*8IH0ME_kOl_C#DD+84RF0IMF2RjRRFV#_08DHFoO#;
HNoMDkRF0k_L#:.RR0Fk_#Lk.$_0bRC;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RV_Rs80FkRM5HbRk000FRs#H-0CN0#02
$RbCF_k0Lck#_b0$C#RHRsNsN5$R80CbEk_MlC_OD-D#4FR8IFM0RRj,cH*I8_0EM_klODCD#R+d8MFI0jFR2VRFR8#0_oDFH
O;#MHoNFDRkL0_kR#c:kRF0k_L#0c_$;bCRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$FsVR_k8F0HR5M0bkRR0F0-sH#00NC
#20C$bR0Fk_#LkU$_0bHCR#sRNsRN$5b8C0ME_kOl_C#DD-84RF0IMF,RjRIU*HE80_lMk_DOCD(#+RI8FMR0FjF2RV0R#8F_Do;HO
o#HMRNDF_k0LUk#RF:RkL0_k_#U0C$b;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFVsF_8k50RHkMb0FR0RH0s-N#002C#
b0$CNRbs$H0_#LkU$_0bHCR#sRNsRN$5b8C0ME_kOl_C#DD-84RF0IMF,RjR8IH0ME_kOl_C#DD-84RF0IMF2RjRRFV#_08DHFoO#;
HNoMDNRbs$H0_#LkURR:bHNs0L$_k_#U0C$b;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RV_Rs80FkRM5HbRk000FRs#H-0CN0#02
$RbCF_k0L4k#n$_0bHCR#sRNsRN$5b8C0ME_kOl_C#DD-84RF0IMF,RjR*4nI0H8Ek_MlC_OD+D#486RF0IMF2RjRRFV#_08DHFoO#;
HNoMDkRF0k_L#R4n:kRF0k_L#_4n0C$b;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFVsF_8k50RHkMb0FR0RH0s-N#002C#
b0$CNRbs$H0_#Lk40n_$RbCHN#Rs$sNRC58b_0EM_klODCD#R-48MFI0jFR,*R.I0H8Ek_MlC_OD+D#4FR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNRsbNH_0$L4k#nRR:bHNs0L$_kn#4_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$FsVR_k8F0HR5M0bkRR0F0-sH#00NC
#20C$bR0Fk_#Lkd0._$RbCHN#Rs$sNRC58b_0EM_klODCD#R-48MFI0jFR,.Rd*8IH0ME_kOl_C#DD+Rd48MFI0jFR2VRFR8#0_oDFH
O;#MHoNFDRkL0_k.#dRF:RkL0_k.#d_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFR8s_FRk05bHMk00RFsR0H0-#N#0C2$
0bbCRN0sH$k_L#_d.0C$bRRH#NNss$8R5CEb0_lMk_DOCD4#-RI8FMR0Fjc,R*8IH0ME_kOl_C#DD+8dRF0IMF2RjRRFV#_08DHFoO#;
HNoMDNRbs$H0_#Lkd:.RRsbNH_0$Ldk#.$_0bRC;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFVsF_8k50RHkMb0FR0RH0s-N#002C#
o#HMRNDF_k0C:MRR8#0_oDFHPO_CFO0sC58b_0EM_klODCD#R-48MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-MRCNCLD#FRVssR0H0-#N#0C
o#HMRNDI_s0C:MRR8#0_oDFHPO_CFO0sC58b_0EM_klODCD#R-48MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-sRIHR0CCLMNDRC#VRFsCENORIsFRRFV)RqvODCD#H
#oDMNR_HMsRCo:0R#8F_Do_HOP0COFIs5HE80+Rd68MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--k8#CRR0FsHCo#s0CRh7QRH
#oDMNR0Fk_osCR#:R0D8_FOoH_OPC05FsI0H8E6+dRI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--k8#CRR0FsHCo#s0CRz7maH
#oDMNR0Fk_osC4RR:#_08DHFoOC_POs0F58IH04E-RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-k-R#RC80OFRE#FFCCRL0CICMQR7hMRN8kRF00bkRRFVAODF	qR)vH
#oDMNR_N8sRCo:0R#8F_Do_HOP0COFNs58I8sHE80-84RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-k-R#RC80sFRC#oH0RCsq)77RsVFRHIs0#C
HNoMDFRDIN_s8R8s:0R#8F_Do_HOP0COF4s5dFR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-NRs8R8sL#H0RbHMk00RFqR)vCRODRD#5LcRHR0#skCJH8sC2H
#oDMNRIDF_8IN8:sRR8#0_oDFHPO_CFO0sd54RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-R8IN8LsRHR0#HkMb0FR0Rv)qRDOCD5#RcHRL0s#RCHJks2C8
o#HMRNDs8N8sC_soRR:#_08DHFoOC_POs0F58N8s8IH04E-RI8FMR0Fj
2;-C-RML8RD	FORlsNRbHlDCClM00NHRFM#MHoN
D#
R--LHCoMCR#D0CORlsNRbHlDCClM00NHRFM#MHoN
D#0C$bRVDC0CFPsR_0HN#Rs$sNRR5j0dFR2VRFR0HMCsoC;$
0bDCRCFV0P_Cs0R_.HN#Rs$sNRR5j04FR2VRFR0HMCsoC;k
VMHO0FbMRNH85R#:R0D8_FOoH_OPC0;FsR,I4RRI.:MRH0CCoss2RCs0kM0R#8F_Do_HOP0COFHsR#N
PsLHNDPCRN:sRR8#0_oDFHPO_CFO0s45I-84RF0IMF2Rj;C
Lo
HMRFRVsRR[HPMRNss'NCMoRFDFbR
RRVRHRR5[<I=R.02RERCM
RSRP5Ns[:2R=5RHHF'DI2+[;C
SD
#CSPRRN[s52=R:R''j;C
SMH8RVR;
R8CMRFDFbR;
R0sCkRsMP;Ns
8CMR8bN;k
VMHO0FoMRCI0_HE80_IU5HE80:MRH0CCoss2RCs0kMMRH0CCos#RH
sPNHDNLCNRPDRR:HCM0oRCs:j=R;C
Lo
HMRNRPD=R:R8IH0UE/;R
RH5VR58IH0lERFU8R2RR>c02RE
CMRRRRPRND:P=RN+DRR
4;RMRC8VRH;R
RskC0sPMRN
D;CRM8o_C0I0H8E;_U
MVkOF0HMCRo0H_I8_0E.H5I8:0ER0HMCsoC2CRs0MksR0HMCsoCR
H#PHNsNCLDRDPNRH:RMo0CC:sR=;Rj
oLCHRM
RDPNRR:=I0H8E;/.
sRRCs0kMNRPDC;
Mo8RCI0_HE80_
.;VOkM0MHFR0oC_8IH0IE5HE80RH:RMo0CCRs2skC0sDMRCFV0P_Cs0R_.HP#
NNsHLRDCPRND:CRDVP0FC0s__
.;LHCoMR
RP5ND4:2R=CRo0H_I8_0E.H5I820E;R
RH5VRI0H8EFRl8RR.=2RjRC0EMR
RRNRPD25jRR:=jR;
R#CDCR
RRNRPD25jRR:=4R;
R8CMR;HV
sRRCs0kMNRPDC;
Mo8RCI0_HE80;k
VMHO0FoMRCI0_HE8058IH0:ERR0HMCsoC2CRs0MksRVDC0CFPsR_0HP#
NNsHLRDCPRND:CRDVP0FC0s_RR:=5Rj,jj,R,2Rj;C
Lo
HMRNRPD25dRR:=o_C0I0H8E5_UI0H8E
2;RNRO#5CRI0H8EFRl82RUR
H#RERICcMRRd|RRR=>P5ND.:2R=;R4
IRRERCM.>R=RDPN5R42:4=R;R
RIMECR=4R>NRPD25jRR:=4R;
RCIEM0RFE#CsRR=>MDkD;R
RCRM8OCN#;R
RskC0sPMRN
D;CRM8o_C0I0H8EO;
F0M#NRM0#H_I8_0ENNss$RR:D0CVFsPC_:0R=CRo0H_I850EI0H8E
2;O#FM00NMRI#_HE80_sNsNn$_cRR:D0CVFsPC_.0_RR:=o_C0I0H8EH5I820E;k
VMHO0FoMRCM0_k4l_.8U5CEb0:MRH0CCoss2RCs0kMMRH0CCos#RH
sPNHDNLCNRPDRR:HCM0oRCs:j=R;C
Lo
HMRNRPD=R:Rb8C04E/.
U;RVRHR855CEb0R8lFRU4.2RR>424.RC0EMR
RRNRPD=R:RDPNR4+R;R
RCRM8H
V;RCRs0MksRDPN;M
C8CRo0k_Ml._4UV;
k0MOHRFMo_C0D0CVFsPC_5nc80CbERR:HCM0o2CsR0sCkRsMHCM0oRCsHL#
CMoH
sRRCs0kMC58bR0ElRF842.U;M
C8CRo0C_DVP0FCns_cV;
k0MOHRFMo_C0M_kln8c5CEb0RH:RMo0CCRs2skC0sHMRMo0CCHsR#N
PsLHNDPCRN:DRR0HMCsoCRR:=jL;
CMoH
HRRV8R5CEb0RR<=4R4.NRM880CbERR>cRU20MEC
RRRRNRPD=R:R
4;RMRC8VRH;R
RskC0sPMRN
D;CRM8o_C0M_kln
c;VOkM0MHFR0oC_VDC0CFPsC58bR0E:MRH0CCosl;RN:GRR0HMCsoC2CRs0MksR0HMCsoCR
H#PHNsNCLDRDPNRH:RMo0CC:sR=;Rj
oLCHRM
RRHV5b8C0-ERRGlNRR>=j02RE
CMRRRRPRND:8=RCEb0Rl-RN
G;RDRC#RC
RPRRN:DR=CR8b;0E
CRRMH8RVR;
R0sCk5sMP2ND;M
C8CRo0C_DVP0FC
s;VOkM0MHFR0oC_lMk_5d.80CbERR:HCM0o2CsR0sCkRsMHCM0oRCsHP#
NNsHLRDCPRND:MRH0CCos=R:R
j;LHCoMR
RH5VR80CbE=R<RRcUNRM880CbERR>4Rn20MEC
RRRRNRPD=R:R
4;RMRC8VRH;R
RskC0sPMRN
D;CRM8o_C0M_kld
.;VOkM0MHFR0oC_lMk_54n80CbERR:HCM0o2CsR0sCkRsMHCM0oRCsHP#
NNsHLRDCPRND:MRH0CCos=R:R
j;LHCoMR
RH5VR80CbE=R<RR4nNRM880CbERR>j02RE
CMRRRRRDPNRR:=4R;
R8CMR;HV
sRRCs0kMNRPDC;
Mo8RCM0_k4l_n-;
-MOF#M0N0kRMlC_ODRD#:MRH0CCos=R:R55580CbERR-4/2RR2d.R5+R5C58bR0E-2R4R8lFR2d.R4/Rn;22R-RR-RRyF)VRq.vdXR41ODCD#CRMC88CRF
OMN#0MM0RkOl_C_DD4R.U:MRH0CCos=R:R0oC_lMk_U4.5b8C0;E2
MOF#M0N0CRDVP0FCns_cRR:HCM0oRCs:o=RCD0_CFV0P_Csn8c5CEb02O;
F0M#NRM0M_klODCD_Rnc:MRH0CCos=R:R0oC_lMk_5ncD0CVFsPC_2nc;F
OMN#0MD0RCFV0P_Csd:.RR0HMCsoCRR:=o_C0D0CVFsPC5VDC0CFPsc_n,cRn2O;
F0M#NRM0M_klODCD_Rd.:MRH0CCos=R:R0oC_lMk_5d.D0CVFsPC_2d.;F
OMN#0MD0RCFV0P_Cs4:nRR0HMCsoCRR:=o_C0D0CVFsPC5VDC0CFPs._d,.Rd2O;
F0M#NRM0M_klODCD_R4n:MRH0CCos=R:R0oC_lMk_54nD0CVFsPC_24n;0

$RbCF_k0L_k#0C$b_U4.RRH#NNss$MR5kOl_C_DD4R.U8MFI0jFR,HRI8-0E4FR8IFM0RRj2F#VR0D8_FOoH;$
0bFCRkL0_k0#_$_bCnHcR#sRNsRN$5lMk_DOCDc_nRI8FMR0FjI,RHE80-84RF0IMF2RjRRFV#_08DHFoO0;
$RbCF_k0L_k#0C$b_Rd.HN#Rs$sNRk5MlC_ODdD_.FR8IFM0RRj,I0H8ER-48MFI0jFR2VRFR8#0_oDFH
O;0C$bR0Fk_#Lk_b0$Cn_4RRH#NNss$MR5kOl_C_DD48nRF0IMF,RjR8IH04E-RI8FMR0FjF2RV0R#8F_Do;HO
o#HMRNDF_k0L_k#4R.U:kRF0k_L#$_0b4C_.RU;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RVFR8k50RHkMb0FR0RH0s-N#002C#
o#HMRNDF_k0L_k#n:cRR0Fk_#Lk_b0$Cc_n;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFV80FkRM5HbRk000FRs#H-0CN0##2
HNoMDkRF0k_L#._dRF:RkL0_k0#_$_bCdR.;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RVFR8k50RHkMb0FR0RH0s-N#002C#
o#HMRNDF_k0L_k#4:nRR0Fk_#Lk_b0$Cn_4;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFV80FkRM5HbRk000FRs#H-0CN0##2
HNoMD_R#F_k0C:MRR8#0_oDFHPO_CFO0sk5MlC_OD4D_.8URF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RNCML#DCRsVFRH0s-N#00
C##MHoNFDRkC0_Mc_nR#:R0D8_FOoH;H
#oDMNR0Fk__CMd:.RR8#0_oDFH
O;#MHoNFDRkC0_Mn_4R#:R0D8_FOoH;H
#oDMNRI#_sC0_MRR:#_08DHFoOC_POs0F5lMk_DOCD._4UFR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--I0sHCMRCNCLD#FRVsNRCOsERFFIRVqR)vCROD
D##MHoNIDRsC0_Mc_nR#:R0D8_FOoH;H
#oDMNR0Is__CMd:.RR8#0_oDFH
O;#MHoNIDRsC0_Mn_4R#:R0D8_FOoH;H
#oDMNRH#_MC_soRR:#_08DHFoOC_POs0F58IH04E-RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RCk#8FR0RosCHC#0sQR7h#R
HNoMD_R#F_k0sRCo:0R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-#RkC08RFCRso0H#C7sRm
za#MHoN#DR__N8sRCo:0R#8F_Do_HOP0COFNs58I8sHE80-84RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-k-R#RC80sFRC#oH0RCsq)77
o#HMRNDD_FINs88R#:R0D8_FOoH_OPC05FsnFR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-8RN8LsRHR0#HkMb0FR0Rv)qRDOCD5#RcHRL0s#RCHJks2C8
MOF#M0N0#RDLH_I8R0E:MRH0CCos=R:R8IH0UE-*_5#I0H8Es_Ns5N$d42-2*-c#H_I8_0ENNss$25.-#.*_8IH0NE_s$sN5-42#H_I8_0ENNss$25j;$
0b0CRlNb_s$sNU#RHRsNsN5$R#H_I8_0ENNss$25d-84RF0IMF2RjRRFV#_08DHFoOC_POs0F58(RF0IMF2Rj;H
#oDMNRb0l_dU_.0,RlUb__R4n:lR0bs_NsUN$;-
-R8CMRD#CCRO0sRNlHDlbCMlC0HN0F#MRHNoMDN#
0H0sLCk0Rs\3NFl_VCV#0:\RRs#0H;Mo
C
Lo
HMRRR
RdzcRH:RVNR58_8ss2CoRMoCC0sNC-R-RMoCC0sNCDRLFRO	s
NlRRRR-Q-RV8RN8HsI8R0E<EROFCHO_8IH0NER#o#HMjR''FR0RkkM#RC8L#H0
RRRRRzjRH:RVNR58I8sHE80R4=R2CRoMNCs0RC
RRRRRDRRFsI_Ns88RR<="jjjjjjjjjjjjRj"&7Rq7j)52R;
RRRRRDRRFII_Ns88RR<="jjjjjjjjjjjjRj"&8RN_osC5;j2
RRRR8CMRMoCC0sNCjRz;R
RR4RzRRR:H5VRNs88I0H8ERR=.o2RCsMCN
0CRRRRRRRRD_FIs8N8s=R<Rj"jjjjjjjjjjRj"&7Rq74)5RI8FMR0Fj
2;RRRRRRRRD_FII8N8s=R<Rj"jjjjjjjjjjRj"&8RN_osC584RF0IMF2Rj;R
RRMRC8CRoMNCs0zCR4R;
RzRR.:RRRRHV58N8s8IH0=ERRRd2oCCMsCN0
RRRRRRRRIDF_8sN8<sR=jR"jjjjjjjjjRj"&7Rq7.)5RI8FMR0Fj
2;RRRRRRRRD_FII8N8s=R<Rj"jjjjjjjjjj&"RR_N8s5Co.FR8IFM0R;j2
RRRR8CMRMoCC0sNC.Rz;R
RRdRzRRR:H5VRNs88I0H8ERR=co2RCsMCN
0CRRRRRRRRD_FIs8N8s=R<Rj"jjjjjjjjj"RR&q)7758dRF0IMF2Rj;R
RRRRRRFRDIN_I8R8s<"=RjjjjjjjjjRj"&8RN_osC58dRF0IMF2Rj;R
RRMRC8CRoMNCs0zCRdR;
RzRRc:RRRRHV58N8s8IH0=ERRR62oCCMsCN0
RRRRRRRRIDF_8sN8<sR=jR"jjjjjjjj"RR&q)7758cRF0IMF2Rj;R
RRRRRRFRDIN_I8R8s<"=Rjjjjjjjjj&"RR_N8s5CocFR8IFM0R;j2
RRRR8CMRMoCC0sNCcRz;R
RR6RzRRR:H5VRNs88I0H8ERR=no2RCsMCN
0CRRRRRRRRD_FIs8N8s=R<Rj"jjjjjjRj"&7Rq76)5RI8FMR0Fj
2;RRRRRRRRD_FII8N8s=R<Rj"jjjjjjRj"&8RN_osC586RF0IMF2Rj;R
RRMRC8CRoMNCs0zCR6R;
RzRRn:RRRRHV58N8s8IH0=ERRR(2oCCMsCN0
RRRRRRRRIDF_8sN8<sR=jR"jjjjjRj"&7Rq7n)5RI8FMR0Fj
2;RRRRRRRRD_FII8N8s=R<Rj"jjjjjj&"RR_N8s5ConFR8IFM0R;j2
RRRR8CMRMoCC0sNCnRz;R
RR(RzRRR:H5VRNs88I0H8ERR=Uo2RCsMCN
0CRRRRRRRRD_FIs8N8s=R<Rj"jjjjj"RR&q)7758(RF0IMF2Rj;R
RRRRRRFRDIN_I8R8s<"=RjjjjjRj"&8RN_osC58(RF0IMF2Rj;R
RRMRC8CRoMNCs0zCR(R;
RzRRU:RRRRHV58N8s8IH0=ERRRg2oCCMsCN0
RRRRRRRRIDF_8sN8<sR=jR"jjjj"RR&q)7758URF0IMF2Rj;R
RRRRRRFRDIN_I8R8s<"=Rjjjjj&"RR_N8s5CoUFR8IFM0R;j2
RRRR8CMRMoCC0sNCURz;R
RRgRzRRR:H5VRNs88I0H8ERR=4Rj2oCCMsCN0
RRRRRRRRIDF_8sN8<sR=jR"j"jjRq&R757)gFR8IFM0R;j2
RRRRRRRRIDF_8IN8<sR=jR"j"jjRN&R8C_soR5g8MFI0jFR2R;
RCRRMo8RCsMCNR0Cz
g;RRRRzR4jRH:RVNR58I8sHE80R4=R4o2RCsMCN
0CRRRRRRRRD_FIs8N8s=R<Rj"jj&"RR7q7)j54RI8FMR0Fj
2;RRRRRRRRD_FII8N8s=R<Rj"jj&"RR_N8s5Co48jRF0IMF2Rj;R
RRMRC8CRoMNCs0zCR4
j;RRRRzR44RH:RVNR58I8sHE80R4=R.o2RCsMCN
0CRRRRRRRRD_FIs8N8s=R<Rj"j"RR&q)775R448MFI0jFR2R;
RRRRRDRRFII_Ns88RR<=""jjRN&R8C_so454RI8FMR0Fj
2;RRRRCRM8oCCMsCN0R4z4;R
RR4Rz.:RRRRHV58N8s8IH0=ERR24dRMoCC0sNCR
RRRRRRFRDIN_s8R8s<'=Rj&'RR7q7).54RI8FMR0Fj
2;RRRRRRRRD_FII8N8s=R<R''jRN&R8C_so.54RI8FMR0Fj
2;RRRRCRM8oCCMsCN0R.z4;R
RR4Rzd:RRRRHV58N8s8IH0>ERR24dRMoCC0sNCR
RRRRRRFRDIN_s8R8s<q=R757)48dRF0IMF2Rj;R
RRRRRRFRDIN_I8R8s<N=R8C_sod54RI8FMR0Fj
2;RRRRCRM8oCCMsCN0Rdz4;R

R-RR-VRQRH58MC_sos2RC#oH0RCs7RQhkM#HopRBiR
RR4Rzc:RRRRHV5M8H_osC2CRoMNCs0RC
RRRRRbRRsCFO#5#RB,piRh7Q2CRLo
HMRRRRRRRRRRRRH5VRBRpi=4R''MRN8pRBiP'CC2M0RC0EMR
RRRRRRRRRRRRRRMRH_osCRR<=5j"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjRj"&QR7h
2;RRRRRRRRRRRRCRM8H
V;RRRRRRRRCRM8bOsFC;##
RRRR8CMRMoCC0sNC4RzcR;
RzRR4R6R:VRHRF5M0HR8MC_soo2RCsMCN
0CRRRRRRRRRRRRHsM_C<oR="R5jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"RR&72Qh;R
RRMRC8CRoMNCs0zCR4
6;
RRRRR--Q5VRsk8F0C_sos2RC#oH0RCs)m_7zkaR#oHMRm)_B
piRRRRzR4nRH:RV8R5F_k0s2CoRMoCC0sNCR
RRRRRRsRbF#OC#mR5B,piR0Fk_osC4L2RCMoH
RRRRRRRRRRRRRHV5pmBiRR='R4'NRM8miBp'CCPMR020MEC
RRRRRRRRRRRRRRRRz7ma=R<R0Fk_osC4R;
RRRRRRRRRCRRMH8RVR;
RRRRRCRRMb8RsCFO#
#;RRRRRRRRCRM8oCCMsCN0Rnz4;R
RR4Rz(:RRRRHV50MFRk8F0C_soo2RCsMCN
0CRRRRRRRRRRRR7amzRR<=F_k0s4Co;R
RRMRC8CRoMNCs0zCR4
(;
RRRRR--Q5VRNs88_osC2CRso0H#CqsR7R7)VRFsI0sHC#RkHRMoB
piRRRRzI4URRR:H5VRNs88_osC2CRoMNCs0RC
RRRRRbRRsCFO#5#RB,piR7q7)L2RCMoH
RRRRRRRRRRRRRHV5iBpR'=R4N'RMB8RpCi'P0CM2ER0CRM
RRRRRRRRRRRRRNRR8C_so=R<R7q7)85N8HsI8-0E4FR8IFM0R;j2
RRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMRFbsO#C#;R
RRMRC8CRoMNCs0zCR4;UI
RRRRgz4IRR:H5VRMRF0Ns88_osC2CRoMNCs0RC
RRRRRRRRRNRR8C_so=R<R7q7)R;
RCRRMo8RCsMCNR0CzI4g;R

R-RR-GR 0RsNDHFoOFRVskR7NbDRFRs0OCN#
-S-RR7FMRF0M8CCRH0E#FRVsFRMRFoDkDCRFOoHRMOF8HH0F-M
-RRRRCzsoRR:bOsFC5##B2piRoLCH-M
-RRRRHRRVBR5p i'ea hR8NMRiBpR'=R4R'20MEC
R--RRRRRQR7hl_0b=R<Rh7Q;-
-RRRRR)RRq)77_b0lRR<=q)77;-
-RRRRRWRRq)77_b0lRR<=Ns8_C
o;-R-RRRRRR_W 0Rlb<W=R -;
-RRRRCRRMH8RV-;
-RRRR8CMRFbsO#C#;R

RzRRlRkG:sRbF#OC#k5F0C_soR2
RRRRRoLCH-M
-RRRRRRRRRHV57Wq70)_l=bRR7)q70)_lNbRMW8R l_0bRR='24'RC0EM-
-RRRRRRRRRkRF0C_so<4R=QR7hl_0b-;
-RRRRRRRR#CDCR
RRRRRRRRRF_k0s4CoRR<=F_k0s5CoI0H8ER-48MFI0jFR2-;
-RRRRRRRR8CMR;HV
RRRR8CMRFbsO#C#;R
RRRRRRRR
R-RR-CRtMNCs00CRE)CRqOvRC#DDR8NMRD#CCRO0DHFoOFRVsqR)vnA4__141R4
RzRR4:URRRHV5FOEH_OCI0H8ERR=4o2RCsMCN
0CSR--VRHGVRFsODNDRU4dUR(,#CCDOF0RVsR0HN#00MCRFL0RCoHMRosCHC#0s
C8SRRRRzRRORE	:VRHRN5R8I8sHE80R4>Rco2RCsMCN
0CRRRRRRRRRRRRk	OD:sRbF#OC#p5BiR2
RRRRRRRRRRRRLHCoMR
RRRRRRRRRRRRRH5VRB'piCMPC0MRN8pRBiRR='24'RC0EMR
RRRRRRRRRRRRRRNRs8_8ss5CoNs88I0H8ER-48MFI04FRc<2R=7Rq7N)58I8sHE80-84RF0IMFcR42R;
RRRRRRRRRRRRR8CMR;HV
RRRRRRRRRRRR8CMRFbsO#C#;S
SRMRC8CRoMNCs0zCRO;E	
RRRRRRRRgz4RV:RFHsRRRHM5b8C0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CRRRR-Q-RVNR58I8sHE80R4>RcM2RCRC80OFRs0CNCsRIHR0CCLMNDNCRMF8Rkk0b0MRCNCLDRD#CCRO0DHFoOR
RRRRRRRRRR.RzjRR:H5VRNs88I0H8ERR>4Rc2oCCMsCN0
-S-RGVHRsVFRDONDdR4U,U(RD#CCRO0F0VRs0H#NR0CMRF0LMCHoCRso0H#C8sC
RRRRRRRRRRRRRRRR0Fk_5CMH<2R=4R''ERIC5MRs8N8sC_so85N8HsI8-0E4FR8IFM0R24cRH=R2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0CHM52=R<RRW IMECR85N_osC58N8s8IH04E-RI8FMR0F4Rc2=2RHR#CDCjR''R;
RRRRRRRRRCRRMo8RCsMCNR0Cz;.j
RRRRR--Q5VRNs88I0H8E=R<R24cRRMFI0sHCMRCNCLDRRFsFbk0kC0RMDNLCCR#D0CORoDFHMORCCC88R
RRRRRRRRRR.Rz4RR:H5VRNs88I0H8E=R<R24cRMoCC0sNCR
RRRRRRRRRRRRRRkRF0M_C5RH2<'=R4
';RRRRRRRRRRRRRRRRI_s0CHM52=R<R;W 
RRRRRRRRRRRR8CMRMoCC0sNC.Rz4R;
R-RR-CRtMNCs00CRE)CRqOvRC#DDR8NMRH0s-N#00
C#RRRRRRRRRRRRzR..:FRVsRR[H5MRI0H8Ek_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0RC
RRRRRRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)RAq4v_ncdUXR47:NRDLRCDH"#RW
";RRRRRRRRRRRRRRRRLHCoMR
RRRRRRRRRRRRRR)RAq4v_ncdUXR47:qR)vnA4__141R4
RRRRRRRRRRRRRbRRFRs0lRNb5q7Q5Rj2=H>RMC_so25[,7Rq7R)q=D>RFII_Ns885R4d8MFI0jFR27,RQ=AR>jR""q,R7A7)RR=>D_FIs8N8sd54RI8FMR0Fj
2,RRRRRRRRRRRRRRRR Rhq='>R4R',1q1)RR=>',j'RqW RR=>I_s0CHM52B,RpRiq=B>RpRi, RhA='>R4R',1A1)RR=>',j'RAW RR=>',j'RiBpA>R=RiBp,R
RRRRRRRRRRRRRRmR7q>R=RCFbM7,RmjA52>R=R0Fk_#Lk4,5H[;22
R
RRRRRRRRRRRRRRkRF0C_so25[RR<=F_k0L4k#5[H,2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRCRRMo8RCsMCNR0Cz;..
RRRRRRRR8CMRMoCC0sNC4RzgR;
RCRRMo8RCsMCNR0Cz;4URRRR
RRRR
RRRRRR-t-RCsMCNR0C0REC)RqvODCD#MRN8CR#D0CORoDFHVORF)sRq4vAn._1_
1.RRRRzR.d:VRHRE5OFCHO_8IH0=ERRR.2oCCMsCN0
-S-RGVHRsVFRDONDdR4U,U(RD#CCRO0F0VRs0H#NR0CMRF0LMCHoCRso0H#C8sC
RSRRzRRO:E	RRHV58N8s8IH0>ERR24dRMoCC0sNCR
RRRRRRRRRRORkDR	:bOsFC5##B2pi
RRRRRRRRRRRRCRLo
HMRRRRRRRRRRRRRVRHRp5BiP'CCRM0NRM8BRpi=4R''02RE
CMRRRRRRRRRRRRRRRRs8N8sC_so85N8HsI8-0E4FR8IFM0R24dRR<=q)7758N8s8IH04E-RI8FMR0F4;d2
RRRRRRRRRRRRCRRMH8RVR;
RRRRRRRRRCRRMb8RsCFO#
#;SCSRMo8RCsMCNR0Cz	OE;R
RRRRRR.RzcRR:VRFsHMRHRC58b_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
RRRRR--Q5VRNs88I0H8ERR>4Rd2M8CCRR0FONsC0ICRsCH0RNCMLRDCNRM8Fbk0kC0RMDNLCCR#D0CORoDFHRO
RRRRRRRRRzRR.:6RRRHV58N8s8IH0>ERR24dRMoCC0sNC-
S-HRVGFRVsNROD4DRd(UU,CR#D0CORRFV0#sH0CN0R0MFRHLCMsoRC#oH0CCs8R
RRRRRRRRRRRRRRkRF0M_C5RH2<'=R4I'RERCM58sN8ss_CNo58I8sHE80-84RF0IMFdR42RR=HC2RDR#C';j'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RWRCIEMNR58C_so85N8HsI8-0E4FR8IFM0R24dRH=R2DRC#'CRj
';RRRRRRRRRRRRCRM8oCCMsCN0R6z.;R
RR-R-RRQV58N8s8IH0<ER=dR42FRMRHIs0CCRMDNLCsRFR0FkbRk0CLMND#CRCODC0FRDoRHOM8CCCR8
RRRRRRRRRzRR.:nRRRHV58N8s8IH0<ER=dR42CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_M25HRR<=';4'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RW;R
RRRRRRRRRRMRC8CRoMNCs0zCR.
n;RRRR-t-RCsMCNR0C0REC)RqvODCD#MRN8sR0H0-#N#0C
RRRRRRRRRRRR(z.RV:RF[sRRRHM58IH0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CRRRRRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FAVR)_qvU.4gXR.7:NRDLRCDH"#RW
";RRRRRRRRRRRRRRRRLHCoMR
RRRRRRRRRRRRRR)RAqUv_4Xg..:7RRv)qA_4n11._.R
RRRRRRRRRRRRRRFRbsl0RN5bR7RQq=H>RMC_so*5.[R+48MFI0.FR*,[2R7q7)=qR>FRDIN_I858s48.RF0IMF2Rj,QR7A>R=Rj"j"q,R7A7)RR=>D_FIs8N8s.54RI8FMR0Fj
2,RRRRRRRRRRRRRRRR Rhq='>R4R',1q1)RR=>',j'RqW RR=>I_s0CHM52B,RpRiq=B>RpRi, RhA='>R4R',1A1)RR=>',j'RAW RR=>',j'RiBpA>R=RiBp,R
RRRRRRRRRRRRRRmR7q>R=RCFbM7,Rm4A52>R=R0Fk_#Lk.,5H.+*[4R2,75mAj=2R>kRF0k_L#H.5,*R.[;22
RRRRRRRRRRRRRRRR0Fk_osC5[.*2=R<R0Fk_#Lk.,5H.2*[RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so*5.[2+4RR<=F_k0L.k#5.H,*4[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRCRRMo8RCsMCNR0Cz;.(
RRRRRRRR8CMRMoCC0sNC.RzcR;
RCRRMo8RCsMCNR0Cz;.dR
R
RRRRRRRR-t-RCsMCNR0C0REC)RqvODCD#MRN8CR#D0CORoDFHVORF)sRq4vAnc_1_
1cRRRRzR.U:VRHRE5OFCHO_8IH0=ERRRc2oCCMsCN0
-S-RGVHRsVFRDONDdR4U,U(RD#CCRO0F0VRs0H#NR0CMRF0LMCHoCRso0H#C8sC
RSRRRRRz	OE:VRHR85N8HsI8R0E>.R42CRoMNCs0RC
RRRRRRRRRkRRO:D	RFbsO#C#5iBp2R
RRRRRRRRRRLRRCMoH
RRRRRRRRRRRRHRRVBR5pCi'P0CMR8NMRiBpR'=R4R'20MEC
RRRRRRRRRRRRRRRR8sN8ss_CNo58I8sHE80-84RF0IMF.R42=R<R7q7)85N8HsI8-0E4FR8IFM0R24.;R
RRRRRRRRRRRRRCRM8H
V;RRRRRRRRRRRRCRM8bOsFC;##
RSSR8CMRMoCC0sNCORzE
	;RRRRRRRRzR.g:FRVsRRHH5MR80CbEk_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0RC
R-RR-VRQR85N8HsI8R0E>.R42CRMC08RFsROCCN0RHIs0CCRMDNLCMRN8kRF00bkRNCMLRDC#CCDOD0RFOoH
RRRRRRRRRRRRjzdRH:RVNR58I8sHE80R4>R.o2RCsMCN
0CSR--VRHGVRFsODNDRU4dUR(,#CCDOF0RVsR0HN#00MCRFL0RCoHMRosCHC#0s
C8RRRRRRRRRRRRRRRRF_k0CHM52=R<R''4RCIEMsR5Ns88_osC58N8s8IH04E-RI8FMR0F4R.2=2RHR#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=WI RERCM5_N8s5CoNs88I0H8ER-48MFI04FR.=2RRRH2CCD#R''j;R
RRRRRRRRRRMRC8CRoMNCs0zCRd
j;RRRR-Q-RVNR58I8sHE80RR<=4R.2MIFRsCH0RNCMLRDCFFsRkk0b0MRCNCLDRD#CCRO0DHFoOCRMC88C
RRRRRRRRRRRR4zdRH:RVNR58I8sHE80RR<=4R.2oCCMsCN0
RRRRRRRRRRRRRRRR0Fk_5CMH<2R=4R''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=W
 ;RRRRRRRRRRRRCRM8oCCMsCN0R4zd;R
RR-R-RMtCC0sNCER0CqR)vCRODRD#NRM80-sH#00NCR#
RRRRRRRRRzRRd:.RRsVFRH[RMIR5HE80_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNCR
RRRRRRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqA)vj_cgcnX7RR:DCNLD#RHR""W;R
RRRRRRRRRRRRRRCRLo
HMRRRRRRRRRRRRRRRRAv)q_gcjn7XcR):Rq4vAnc_1_
1cRRRRRRRRRRRRRRRRb0FsRblNRQ57q>R=R_HMs5Coc+*[dFR8IFM0R[c*2q,R7q7)RR=>D_FII8N8s454RI8FMR0FjR2,7RQA=">Rjjjj"q,R7A7)RR=>D_FIs8N8s454RI8FMR0Fj
2,RRRRRRRRRRRRRRRR Rhq='>R4R',1q1)RR=>',j'RqW RR=>I_s0CHM52B,RpRiq=B>RpRi, RhA='>R4R',1A1)RR=>',j'RAW RR=>',j'RiBpA>R=RiBp,R
RRRRRRRRRRRRRRmR7q>R=RCFbM7,RmdA52>R=R0Fk_#Lkc,5HR[c*+,d2RA7m5R.2=F>RkL0_k5#cH*,c[2+.,RR
RRRRRRRRRRRRR7RRm4A52>R=R0Fk_#Lkc,5Hc+*[4R2,75mAj=2R>kRF0k_L#Hc5,*Rc[;22
RRRRRRRRRRRRRRRR0Fk_osC5[c*2=R<R0Fk_#Lkc,5Hc2*[RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so*5c[2+4RR<=F_k0Lck#5cH,*4[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cco5*.[+2=R<R0Fk_#Lkc,5Hc+*[.I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Coc+*[d<2R=kRF0k_L#Hc5,[c*+Rd2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
R
RRRRRRRRRRMRC8CRoMNCs0zCRd
.;RRRRRRRRCRM8oCCMsCN0Rgz.;R
RRMRC8CRoMNCs0zCR.
U;
RRRRRRRRR--tCCMsCN0RC0ERv)qRDOCDN#RM#8RCODC0FRDoRHOVRFs)Aqv41n_gg_1
RRRRdzdRH:RVOR5EOFHCH_I8R0E=2RgRMoCC0sNC-
S-HRVGFRVsNROD4DRd(UU,CR#D0CORRFV0#sH0CN0R0MFRHLCMsoRC#oH0CCs8R
SRRRRREzO	H:RVNR58I8sHE80R4>R4o2RCsMCN
0CRRRRRRRRRRRRk	OD:sRbF#OC#p5BiR2
RRRRRRRRRRRRLHCoMR
RRRRRRRRRRRRRH5VRB'piCMPC0MRN8pRBiRR='24'RC0EMR
RRRRRRRRRRRRRRNRs8_8ss5CoNs88I0H8ER-48MFI04FR4<2R=7Rq7N)58I8sHE80-84RF0IMF4R42R;
RRRRRRRRRRRRR8CMR;HV
RRRRRRRRRRRR8CMRFbsO#C#;S
SRMRC8CRoMNCs0zCRO;E	
RRRRRRRRczdRV:RFHsRRRHM5b8C0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CRRRR-Q-RVNR58I8sHE80R4>R4M2RCRC80OFRs0CNCsRIHR0CCLMNDNCRMF8Rkk0b0MRCNCLDRD#CCRO0DHFoOR
RRRRRRRRRRdRz6RR:H5VRNs88I0H8ERR>4R42oCCMsCN0
-S-RGVHRsVFRDONDdR4U,U(RD#CCRO0F0VRs0H#NR0CMRF0LMCHoCRso0H#C8sC
RRRRRRRRRRRRRRRR0Fk_5CMH<2R=4R''ERIC5MRs8N8sC_so85N8HsI8-0E4FR8IFM0R244RH=R2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0CHM52=R<RRW IMECR85N_osC58N8s8IH04E-RI8FMR0F4R42=2RHR#CDCjR''R;
RRRRRRRRRCRRMo8RCsMCNR0Cz;d6
RRRRR--Q5VRNs88I0H8E=R<R244RRMFI0sHCMRCNCLDRRFsFbk0kC0RMDNLCCR#D0CORoDFHMORCCC88R
RRRRRRRRRRdRznRR:H5VRNs88I0H8E=R<R244RMoCC0sNCR
RRRRRRRRRRRRRRkRF0M_C5RH2<'=R4
';RRRRRRRRRRRRRRRRI_s0CHM52=R<R;W 
RRRRRRRRRRRR8CMRMoCC0sNCdRznR;
R-RR-CRtMNCs00CRE)CRqOvRC#DDR8NMRH0s-N#00
C#RRRRRRRRRRRRzRd(:FRVsRR[H5MRI0H8Ek_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0RC
RRRRRRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)RAq.v_jXcUU:7RRLDNCHDR#WR""R;
RRRRRRRRRRRRRLRRCMoH
RRRRRRRRRRRRRRRRqA)vj_.cUUX7RR:)Aqv41n_gg_1
RRRRRRRRRRRRRRRRbRRFRs0lRNb5q7QRR=>HsM_Cgo5*([+RI8FMR0Fg2*[,7Rq7R)q=D>RFII_Ns885R4j8MFI0jFR27,RQ=AR>jR"jjjjj"jj,7Rq7R)A=D>RFsI_Ns885R4j8MFI0jFR2R,
RRRRRRRRRRRRR RRh=qR>4R''1,R1R)q='>RjR',WR q=I>RsC0_M25H,pRBi=qR>pRBi ,Rh=AR>4R''1,R1R)A='>RjR',WR A='>RjR',BApiRR=>B,piRR
RRRRRRRRRRRRRRmR7q>R=RCFbM7,Rm(A52>R=R0Fk_#LkU,5HU+*[(R2,75mAn=2R>kRF0k_L#HU5,[U*+,n2RR
RRRRRRRRRRRRRRmR7A256RR=>F_k0LUk#5UH,*6[+27,RmcA52>R=R0Fk_#LkU,5HU+*[cR2,75mAd=2R>kRF0k_L#HU5,[U*+,d2RR
RRRRRRRRRRRRRRmR7A25.RR=>F_k0LUk#5UH,*.[+27,Rm4A52>R=R0Fk_#LkU,5HU+*[4R2,75mAj=2R>kRF0k_L#HU5,[U*2R,
RRRRRRRRRRRRRRRRRRRRRRRRR7RRQ5uqj=2R>MRH_osC5[g*+,U2Ru7QA>R=R""j,mR7u=qR>bRFCRM,7Amu5Rj2=b>RN0sH$k_L#HU5,2R[2R;
RRRRRRRRRRRRRFRRks0_Cgo5*R[2<F=RkL0_k5#UH*,U[I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cog+*[4<2R=kRF0k_L#HU5,[U*+R42IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5[g*+R.2<F=RkL0_k5#UH*,U[2+.RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so*5g[2+dRR<=F_k0LUk#5UH,*d[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cgo5*c[+2=R<R0Fk_#LkU,5HU+*[cI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cog+*[6<2R=kRF0k_L#HU5,[U*+R62IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5[g*+Rn2<F=RkL0_k5#UH*,U[2+nRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so*5g[2+(RR<=F_k0LUk#5UH,*([+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cgo5*U[+2=R<RsbNH_0$LUk#5[H,2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRCRRMo8RCsMCNR0Cz;d(
RRRRRRRR8CMRMoCC0sNCdRzcR;
RCRRMo8RCsMCNR0Cz;dd
R
RRRRRR-R-RMtCC0sNCER0CqR)vCRODRD#NRM8#CCDOD0RFOoHRsVFRv)qA_4n1_4U1
4URRRRzRdU:VRHRE5OFCHO_8IH0=ERR24URMoCC0sNC-
S-HRVGFRVsNROD4DRd(UU,CR#D0CORRFV0#sH0CN0R0MFRHLCMsoRC#oH0CCs8R
SRRRRREzO	H:RVNR58I8sHE80R4>Rjo2RCsMCN
0CRRRRRRRRRRRRk	OD:sRbF#OC#p5BiR2
RRRRRRRRRRRRLHCoMR
RRRRRRRRRRRRRH5VRB'piCMPC0MRN8pRBiRR='24'RC0EMR
RRRRRRRRRRRRRRNRs8_8ss5CoNs88I0H8ER-48MFI04FRj<2R=7Rq7N)58I8sHE80-84RF0IMFjR42R;
RRRRRRRRRRRRR8CMR;HV
RRRRRRRRRRRR8CMRFbsO#C#;S
SRMRC8CRoMNCs0zCRO;E	
RRRRRRRRgzdRV:RFHsRRRHM5b8C0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CRRRR-Q-RVNR58I8sHE80R4>RjM2RCRC80OFRs0CNCsRIHR0CCLMNDNCRMF8Rkk0b0MRCNCLDRD#CCRO0DHFoOR
RRRRRRRRRRcRzjRR:H5VRNs88I0H8ERR>4Rj2oCCMsCN0
-S-RGVHRsVFRDONDdR4U,U(RD#CCRO0F0VRs0H#NR0CMRF0LMCHoCRso0H#C8sC
RRRRRRRRRRRRRRRR0Fk_5CMH<2R=4R''ERIC5MRs8N8sC_so85N8HsI8-0E4FR8IFM0R24jRH=R2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0CHM52=R<RRW IMECR85N_osC58N8s8IH04E-RI8FMR0F4Rj2=2RHR#CDCjR''R;
RRRRRRRRRCRRMo8RCsMCNR0Cz;cj
RRRRR--Q5VRNs88I0H8E=R<R24jRRMFI0sHCMRCNCLDRRFsFbk0kC0RMDNLCCR#D0CORoDFHMORCCC88R
RRRRRRRRRRcRz4RR:H5VRNs88I0H8E=R<R24jRMoCC0sNCR
RRRRRRRRRRRRRRkRF0M_C5RH2<'=R4
';RRRRRRRRRRRRRRRRI_s0CHM52=R<R;W 
RRRRRRRRRRRR8CMRMoCC0sNCcRz4R;
R-RR-CRtMNCs00CRE)CRqOvRC#DDR8NMRH0s-N#00
C#RRRRRRRRRRRRzRc.:FRVsRR[H5MRI0H8Ek_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0RC
RRRRRRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)RAq4v_jX.c4Rn7:NRDLRCDH"#RW
";RRRRRRRRRRRRRRRRLHCoMR
RRRRRRRRRRRRRR)RAq4v_jX.c4Rn7:qR)vnA4_U14_U14
RRRRRRRRRRRRRRRRbRRFRs0lRNb5q7QRR=>HsM_C4o5U+*[486RF0IMFUR4*,[2R7q7)=qR>FRDIN_I858sgFR8IFM0R,j2RA7QRR=>"jjjjjjjjjjjjjjjjR",q)77A>R=RIDF_8sN8gs5RI8FMR0Fj
2,RRRRRRRRRRRRRRRR Rhq='>R4R',1q1)RR=>',j'RqW RR=>I_s0CHM52B,RpRiq=B>RpRi, RhA='>R4R',1A1)RR=>',j'RAW RR=>',j'RiBpA>R=RiBp,RR
RRRRRRRRRRRRR7RRm=qR>bRFCRM,75mA4R62=F>RkL0_kn#454H,n+*[4,62RA7m524cRR=>F_k0L4k#n,5H4[n*+24c,RR
RRRRRRRRRRRRR7RRm4A5d=2R>kRF0k_L#54nHn,4*4[+dR2,75mA4R.2=F>RkL0_kn#454H,n+*[4,.2RA7m5244RR=>F_k0L4k#n,5H4[n*+244,RR
RRRRRRRRRRRRR7RRm4A5j=2R>kRF0k_L#54nHn,4*4[+jR2,75mAg=2R>kRF0k_L#54nHn,4*g[+27,RmUA52>R=R0Fk_#Lk4Hn5,*4n[2+U,RR
RRRRRRRRRRRRR7RRm(A52>R=R0Fk_#Lk4Hn5,*4n[2+(,mR7A25nRR=>F_k0L4k#n,5H4[n*+,n2RA7m5R62=F>RkL0_kn#454H,n+*[6R2,
RRRRRRRRRRRRRRRRA7m5Rc2=F>RkL0_kn#454H,n+*[cR2,75mAd=2R>kRF0k_L#54nHn,4*d[+27,Rm.A52>R=R0Fk_#Lk4Hn5,*4n[2+.,RR
RRRRRRRRRRRRR7RRm4A52>R=R0Fk_#Lk4Hn5,*4n[2+4,mR7A25jRR=>F_k0L4k#n,5H4[n*2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRR7qQuRR=>HsM_C4o5U+*[48(RF0IMFUR4*4[+nR2,7AQuRR=>""jj,R
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7u=qR>bRFCRM,7Amu5R42=b>RN0sH$k_L#54nH.,R*4[+27,Rm5uAj=2R>NRbs$H0_#Lk4Hn5,*R.[;22
RRRRRRRRRRRRRRRR0Fk_osC5*4U[<2R=kRF0k_L#54nHn,4*R[2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[2+4RR<=F_k0L4k#n,5H4[n*+R42IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[2+.RR<=F_k0L4k#n,5H4[n*+R.2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[2+dRR<=F_k0L4k#n,5H4[n*+Rd2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[2+cRR<=F_k0L4k#n,5H4[n*+Rc2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[2+6RR<=F_k0L4k#n,5H4[n*+R62IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[2+nRR<=F_k0L4k#n,5H4[n*+Rn2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[2+(RR<=F_k0L4k#n,5H4[n*+R(2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[2+URR<=F_k0L4k#n,5H4[n*+RU2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[2+gRR<=F_k0L4k#n,5H4[n*+Rg2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[j+42=R<R0Fk_#Lk4Hn5,*4n[j+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[4R42<F=RkL0_kn#454H,n+*[4R42IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[.+42=R<R0Fk_#Lk4Hn5,*4n[.+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[4Rd2<F=RkL0_kn#454H,n+*[4Rd2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[c+42=R<R0Fk_#Lk4Hn5,*4n[c+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[4R62<F=RkL0_kn#454H,n+*[4R62IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[n+42=R<RsbNH_0$L4k#n,5H.2*[RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*4[+(<2R=NRbs$H0_#Lk4Hn5,[.*+R42IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRR8CMRMoCC0sNCcRz.R;
RRRRRCRRMo8RCsMCNR0Cz;dg
RRRR8CMRMoCC0sNCdRzU
;
SRRRRR--tCCMsCN0RC0ERv)qRDOCDN#RM#8RCODC0FRDoRHOVRFs)Aqv41n_d1n_dSn
zNdURH:RVOR5EOFHCH_I8R0E=nRd2CRoMNCs0SC
-V-RHVGRFOsRNRDD4UdU(#,RCODC0VRFRH0s#00NCFRM0CRLHRMosHCo#s0CCS8
RRRRRORzER	:H5VRNs88I0H8ERR>go2RCsMCN
0CSRSRRORkDR	:bOsFC5##B2pi
SSSRoLCHSM
SRSRH5VRB'piCMPC0MRN8pRBiRR='24'RC0EMS
SSRRRR8sN8ss_CNo58I8sHE80-84RF0IMF2RgRR<=q)7758N8s8IH04E-RI8FMR0Fg
2;SRSSR8CMR;HV
SSSCRM8bOsFC;##
RSSR8CMRMoCC0sNCORzE
	;SRRRRgzdNRR:VRFsHMRHRC58b_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
-S-RRQV58N8s8IH0>ERRRg2M8CCRR0FONsC0ICRsCH0RNCMLRDCNRM8Fbk0kC0RMDNLCCR#D0CORoDFHSO
ScSzj:NRRRHV58N8s8IH0>ERRRg2oCCMsCN0
-S-RGVHRsVFRDONDdR4U,U(RD#CCRO0F0VRs0H#NR0CMRF0LMCHoCRso0H#C8sC
SSSRRRRF_k0CHM52=R<R''4RCIEMsR5Ns88_osC58N8s8IH04E-RI8FMR0Fg=2RRRH2CCD#R''j;S
SSsSI0M_C5RH2<W=R ERIC5MRNs8_CNo58I8sHE80-84RF0IMF2RgRH=R2DRC#'CRj
';SCSSMo8RCsMCNR0CzNcj;-
S-VRQR85N8HsI8R0E<g=R2FRMRHIs0CCRMDNLCsRFR0FkbRk0CLMND#CRCODC0FRDoRHOM8CCCS8
ScSz4:NRRRHV58N8s8IH0<ER=2RgRMoCC0sNCS
SSkSF0M_C5RH2<'=R4
';SSSSI_s0CHM52=R<R;W 
SSSCRM8oCCMsCN0R4zcNS;
-t-RCsMCNR0C0REC)RqvODCD#MRN8sR0H0-#N#0C
SSSzNc.RV:RF[sRRRHM58IH0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CRRRRRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FAVR)_qv6X4.dR.7:NRDLRCDH"#RW
";RRRRRRRRRRRRRRRRLHCoMS
SS)SAq6v_4d.X.:7RRv)qA_4n1_dn1
dnRRRRRRRRRRRRRRRRRFRbsl0RN5bR7RQq=H>RMC_son5d*d[+4FR8IFM0R*dn[R2,q)77q>R=RIDF_8IN8Us5RI8FMR0FjR2,
SSSSA7QRR=>"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjR",q)77A>R=RIDF_8sN8Us5RI8FMR0Fj
2,SSSS Rhq='>R4R',1q1)RR=>',j'RqW RR=>I_s0CHM52B,RpRiq=B>RpRi, RhA='>R4R',1A1)RR=>',j'RAW RR=>',j'RiBpA>R=RiBp,S
SSmS7q>R=RCFbM7,RmdA54=2R>kRF0k_L#5d.H.,d*d[+4R2,75mAdRj2=F>RkL0_k.#d5dH,.+*[d,j2
SSSSA7m52.gRR=>F_k0Ldk#.,5Hd[.*+2.g,mR7AU5.2>R=R0Fk_#LkdH.5,*d.[U+.27,Rm.A5(=2R>kRF0k_L#5d.H.,d*.[+(
2,SSSS75mA.Rn2=F>RkL0_k.#d5dH,.+*[.,n2RA7m52.6RR=>F_k0Ldk#.,5Hd[.*+2.6,mR7Ac5.2>R=R0Fk_#LkdH.5,*d.[c+.2S,
S7SSm.A5d=2R>kRF0k_L#5d.H.,d*.[+dR2,75mA.R.2=F>RkL0_k.#d5dH,.+*[.,.2RA7m52.4RR=>F_k0Ldk#.,5Hd[.*+2.4,S
SSmS7Aj5.2>R=R0Fk_#LkdH.5,*d.[j+.27,Rm4A5g=2R>kRF0k_L#5d.H.,d*4[+gR2,75mA4RU2=F>RkL0_k.#d5dH,.+*[4,U2
SSSSA7m524(RR=>F_k0Ldk#.,5Hd[.*+24(,mR7An542>R=R0Fk_#LkdH.5,*d.[n+427,Rm4A56=2R>kRF0k_L#5d.H.,d*4[+6
2,SSSS75mA4Rc2=F>RkL0_k.#d5dH,.+*[4,c2RA7m524dRR=>F_k0Ldk#.,5Hd[.*+24d,mR7A.542>R=R0Fk_#LkdH.5,*d.[.+42
,RSSSS75mA4R42=F>RkL0_k.#d5dH,.+*[4,42RA7m524jRR=>F_k0Ldk#.,5Hd[.*+24j,mR7A25gRR=>F_k0Ldk#.,5Hd[.*+,g2RS
SSmS7A25URR=>F_k0Ldk#.,5Hd[.*+,U2RA7m5R(2=F>RkL0_k.#d5dH,.+*[(R2,75mAn=2R>kRF0k_L#5d.H.,d*n[+2
,RSSSS75mA6=2R>kRF0k_L#5d.H.,d*6[+27,RmcA52>R=R0Fk_#LkdH.5,*d.[2+c,mR7A25dRR=>F_k0Ldk#.,5Hd[.*+,d2RS
SSmS7A25.RR=>F_k0Ldk#.,5Hd[.*+,.2RA7m5R42=F>RkL0_k.#d5dH,.+*[4R2,75mAj=2R>kRF0k_L#5d.H.,d*,[2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRQR7u=qR>MRH_osC5*dn[6+dRI8FMR0Fd[n*+2d.,QR7u=AR>jR"j"jj,mR7u=qR>bRFCRM,7Amu5Rd2=b>RN0sH$k_L#5d.H*,c[2+d,R
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7u.A52>R=RsbNH_0$Ldk#.,5Hc+*[.R2,7Amu5R42=b>RN0sH$k_L#5d.H*,c[2+4,mR7ujA52>R=RsbNH_0$Ldk#.,5Hc2*[2R;
RRRRRRRRRRRRRFRRks0_Cdo5n2*[RR<=F_k0Ldk#.,5Hd[.*2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cdo5n+*[4<2R=kRF0k_L#5d.H.,d*4[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cdo5n+*[.<2R=kRF0k_L#5d.H.,d*.[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cdo5n+*[d<2R=kRF0k_L#5d.H.,d*d[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cdo5n+*[c<2R=kRF0k_L#5d.H.,d*c[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cdo5n+*[6<2R=kRF0k_L#5d.H.,d*6[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cdo5n+*[n<2R=kRF0k_L#5d.H.,d*n[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cdo5n+*[(<2R=kRF0k_L#5d.H.,d*([+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cdo5n+*[U<2R=kRF0k_L#5d.H.,d*U[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cdo5n+*[g<2R=kRF0k_L#5d.H.,d*g[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cdo5n+*[4Rj2<F=RkL0_k.#d5dH,.+*[4Rj2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*dn[4+42=R<R0Fk_#LkdH.5,*d.[4+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cdo5n+*[4R.2<F=RkL0_k.#d5dH,.+*[4R.2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*dn[d+42=R<R0Fk_#LkdH.5,*d.[d+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cdo5n+*[4Rc2<F=RkL0_k.#d5dH,.+*[4Rc2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*dn[6+42=R<R0Fk_#LkdH.5,*d.[6+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cdo5n+*[4Rn2<F=RkL0_k.#d5dH,.+*[4Rn2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*dn[(+42=R<R0Fk_#LkdH.5,*d.[(+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cdo5n+*[4RU2<F=RkL0_k.#d5dH,.+*[4RU2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*dn[g+42=R<R0Fk_#LkdH.5,*d.[g+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cdo5n+*[.Rj2<F=RkL0_k.#d5dH,.+*[.Rj2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*dn[4+.2=R<R0Fk_#LkdH.5,*d.[4+.2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cdo5n+*[.R.2<F=RkL0_k.#d5dH,.+*[.R.2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*dn[d+.2=R<R0Fk_#LkdH.5,*d.[d+.2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cdo5n+*[.Rc2<F=RkL0_k.#d5dH,.+*[.Rc2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*dn[6+.2=R<R0Fk_#LkdH.5,*d.[6+.2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cdo5n+*[.Rn2<F=RkL0_k.#d5dH,.+*[.Rn2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*dn[(+.2=R<R0Fk_#LkdH.5,*d.[(+.2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cdo5n+*[.RU2<F=RkL0_k.#d5dH,.+*[.RU2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*dn[g+.2=R<R0Fk_#LkdH.5,*d.[g+.2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cdo5n+*[dRj2<F=RkL0_k.#d5dH,.+*[dRj2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*dn[4+d2=R<R0Fk_#LkdH.5,*d.[4+d2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cdo5n+*[dR.2<b=RN0sH$k_L#5d.H*,c[I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cod[n*+2ddRR<=bHNs0L$_k.#d5cH,*4[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cdo5n+*[dRc2<b=RN0sH$k_L#5d.H*,c[2+.RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_son5d*d[+6<2R=NRbs$H0_#LkdH.5,[c*+Rd2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRR8CMRMoCC0sNCcRz.
N;RRRRRRRRCRM8oCCMsCN0RgzdNR;
RCRRMo8RCsMCNR0CzNdU;R
RCRM8oCCMsCN0Rdzc;R
Rz:ccRRHV50MFR8N8sC_soo2RCsMCNR0C-o-RCsMCNR0C#CCDOs0RNRl
R-RR-VRQR8N8s8IH0<ERRN(R#o#HMjR''FR0RkkM#RC8L#H0
RRRRRzjRH:RVNR58I8sHE80R4=R2CRoMNCs0RC
RRRRRDRRFNI_8R8s<"=RjjjjjRj"&_R#Ns8_Cjo52R;
RCRRMo8RCsMCNR0Cz
j;RRRRzR4R:VRHR85N8HsI8R0E=2R.RMoCC0sNCR
RRRRRRFRDI8_N8<sR=jR"jjjj"RR&#8_N_osC584RF0IMF2Rj;R
RRMRC8CRoMNCs0zCR4R;
RzRR.:RRRRHV58N8s8IH0=ERRRd2oCCMsCN0
RRRRRRRRIDF_8N8s=R<Rj"jjRj"&_R#Ns8_C.o5RI8FMR0Fj
2;RRRRCRM8oCCMsCN0R;z.
RRRRRzdRH:RVNR58I8sHE80Rc=R2CRoMNCs0RC
RRRRRDRRFNI_8R8s<"=Rj"jjR#&R__N8s5CodFR8IFM0R;j2
RRRR8CMRMoCC0sNCdRz;z
ScRS:H5VRNs88I0H8ERR=6o2RCsMCN
0CSFSDI8_N8<sR=jR"j&"RRN#_8C_soR5c8MFI0jFR2S;
CRM8oCCMsCN0R;zc
6SzSH:RVNR58I8sHE80Rn=R2CRoMNCs0SC
SIDF_8N8s=R<R''jR#&R__N8s5Co6FR8IFM0R;j2
RRRR8CMRMoCC0sNC6Rz;R
RRnRzRRR:H5VRNs88I0H8ERR>no2RCsMCN
0CRRRRRRRRD_FINs88RR<=#8_N_osC58nRF0IMF2Rj;R
RRMRC8CRoMNCs0zCRn
;
RRRR-Q-RV8R5HsM_CRo2sHCo#s0CRh7QRHk#MBoRpRi
RzRR(:RRRRHV5M8H_osC2CRoMNCs0RC
RRRRRbRRsCFO#5#RB,piRh7Q2CRLo
HMRRRRRRRRRRRRH5VRBRpi=4R''MRN8pRBiP'CC2M0RC0EMR
RRRRRRRRRRRRRR_R#HsM_C<oR=QR7hR;
RRRRRRRRRCRRMH8RVR;
RRRRRCRRMb8RsCFO#
#;RRRRCRM8oCCMsCN0R;z(
RRRRRzURH:RVMR5F80RHsM_CRo2oCCMsCN0
RRRRRRRRRRRRH#_MC_so=R<Rh7Q;R
RRMRC8CRoMNCs0zCRU
;
RRRR-Q-RV8R5F_k0s2CoRosCHC#0smR7zkaR#oHMRpmBiR
RRgRzRRR:H5VR80Fk_osC2CRoMNCs0RC
RRRRRbRRsCFO#5#RmiBp,kRF0C_soL2RCMoH
RRRRRRRRRRRRRHV5pmBiRR='R4'NRM8miBp'CCPMR020MEC
RRRRRRRRRRRRRRRRz7ma=R<RF#_ks0_C
o;RRRRRRRRRRRRCRM8H
V;RRRRRRRRCRM8bOsFC;##
RRRR8CMRMoCC0sNCgRz;R
RR4Rzj:RRRRHV50MFRk8F0C_soo2RCsMCN
0CRRRRRRRRRRRR7amzRR<=#k_F0C_soR;
RCRRMo8RCsMCNR0Cz;4j
R
RR-R-RRQV58N8sC_sos2RC#oH0RCsq)77RHk#MBoRpRi
RzRR4R4R:VRHR85N8ss_CRo2oCCMsCN0
RRRRRRRRFbsO#C#Rp5Biq,R727)RoLCHRM
RRRRRRRRRHRRVBR5p=iRR''4R8NMRiBp'CCPMR020MEC
RRRRRRRRRRRRRRRRN#_8C_so=R<R7q7)85N8HsI8-0E4FR8IFM0R;j2
RRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMRFbsO#C#;R
RRMRC8CRoMNCs0zCR4
4;RRRRzR4.:VRHRF5M08RN8ss_CRo2oCCMsCN0
RRRRRRRRRRRRN#_8C_so=R<R7q7)R;
RCRRMo8RCsMCNR0Cz;4.
RRRRRRRRR
RR-R-RMtCC0sNCER0CqR)vCRODRD#NRM8#CCDOD0RFOoH
RRRRdz4RV:RFHsRRRHM5lMk_DOCD._4URR-482RF0IMFRRjoCCMsCN0
RRRRR--Q5VRNs88I0H8ERR>6M2RCRC80OFRs0CNCsRIHR0CCLMNDNCRMF8Rkk0b0MRCNCLDRD#CCRO0DHFoOR
RRRRRR4RzcRR:H5VRNs88I0H8ERR>(o2RCsMCN
0CRRRRRRRRRRRRRRRR#k_F0M_C5RH2<'=R4I'RERCM5N#_8C_so85N8HsI8-0E4FR8IFM0RR(2=2RHR#CDCjR''R;
RRRRRRRRRRRRR#RR_0Is_5CMH<2R= RWRCIEM#R5__N8s5CoNs88I0H8ER-48MFI0(FR2RR=HC2RDR#C';j'
RRRRRRRR8CMRMoCC0sNC4RzcR;
R-RR-VRQR85N8HsI8R0E<6=R2FRMRHIs0CCRMDNLCsRFR0FkbRk0CLMND#CRCODC0FRDoRHOM8CCCR8
RRRRRzRR4:6RRRHV58N8s8IH0<ER=2R(RMoCC0sNCR
RRRRRRRRRRRRRR_R#F_k0CHM52=R<R''4;R
RRRRRRRRRRRRRR_R#I_s0CHM52=R<R;W 
RRRRRRRR8CMRMoCC0sNC4Rz6R;
R-RR-CRtMNCs00CRE)CRqOvRC#DDR8NMRH0s-N#00
C#RRRRRRRRzR4n:FRVsRR[H5MRI0H8ERR-482RF0IMFRRjoCCMsCN0
RRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVzv)q4R.U:NRDLRCDH"#R1"1aRH&RMo0CCHs'lCNo58IH0RE2&7R""RR&HCM0o'CsHolNC*5H42.UR"&RW&"RR0HMCsoC'NHlo[C52RR&"R "&MRH0CCosl'HN5oCo_C0C_M880CbEH55+*424,.URb8C02E2R"&RX&"RR0HMCsoC'NHlo[C5+;42
RRRRRRRRRRRRoLCHRM
RRRRRRRRRzRR)4qv.:URRqX)vU4.XR41
RRRRRRRRRRRRRRRRsbF0NRlb7R5RR=>#M_H_osC5,[2RRqj=D>RFNI_858sjR2,q=4R>FRDI8_N84s52q,R.>R=RIDF_8N8s25.,R
RRRRRRRRRRRRRRRRRRRRRRRRRq=dR>FRDI8_N8ds52q,Rc>R=RIDF_8N8s25c,6RqRR=>D_FINs885,62RRqn=D>RFNI_858sn
2,SSSSSRSRW= R>_R#I_s0CHM52W,RBRpi=B>RpRi,m>R=R0Fk_#Lk_U4.5[H,2
2;RRRRRRRRRRRRRRRR#k_F0C_so25[RR<=F_k0L_k#45.UH2,[RCIEM#R5_0Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRCRM8oCCMsCN0Rnz4;R
RRCRRMo8RCsMCNR0Cz;4dRRRRRRRRRRRR
RRRR
RRRRRR-t-RCsMCNR0CNnR4RsIF8CR8C)bRqOvRCRDDHNVRbFbsbNsH0RCRRRRRRRRRRRRRRR
RR4Rz(RR:H5VRM_klODCD_Rnc=2R4RMoCC0sNCR
RR-R-RRQV58N8s8IH0>ERRR(2M8CCRR0FONsC0ICRsCH0RNCMLRDCNRM8Fbk0kC0RMDNLCCR#D0CORoDFHRO
RRRRRzRR4RUN:VRHR85N8HsI8R0E>2R(RMoCC0sNCR
RRRRRRRRRRRRRRkRF0M_C_Rnc<'=R4I'RERCM5_5#Ns8_CNo58I8sHE80-84RF0IMF2R(RM=RkOl_C_DD42.UR8NMR_5#Ns8_Cno52RR='2j'2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0CnM_c=R<RRW IMECR#55__N8s5CoNs88I0H8ER-48MFI0(FR2RR=M_klODCD_U4.2MRN8#R5__N8s5Con=2RR''j2C2RDR#C';j'
RRRRRRRR8CMRMoCC0sNC4RzU
N;RRRRRRRRzL4URH:RVNR58I8sHE80R(=RR8NMRlMk_DOCD._4URR=jo2RCsMCN
0CRRRRRRRRRRRRRRRRF_k0CnM_c=R<R''4RCIEM5R5#8_N_osC5Rn2=jR''R22CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C_Rnc<W=R ERIC5MR5N#_8C_so25nR'=Rj2'2R#CDCjR''R;
RRRRRCRRMo8RCsMCNR0CzL4U;R
RR-R-RRQV58N8s8IH0<ER=2R6RRMFI0sHCMRCNCLDRRFsFbk0kC0RMDNLCCR#D0CORoDFHMORCCC88R
RRRRRR4RzgRR:H5VRNs88I0H8E=R<RRn2oCCMsCN0
RRRRRRRRRRRRRRRR0Fk__CMn<cR=4R''R;
RRRRRRRRRRRRRIRRsC0_Mc_nRR<=W
 ;RRRRRRRRCRM8oCCMsCN0Rgz4;R
RR-R-RMtCC0sNCER0CqR)vCRODNDRM08Rs#H-0CN0
RSRRORzE.	_RH:RV#R5_8IH0NE_s$sN_5nc4>2RRRj2oCCMsCN0
RRRRRRRRjz.RV:RF[sRRRHM5I#_HE80_sNsNn$_c254R4-R2FR8IFM0RojRCsMCN
0CRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FzVR)nqvcRR:DCNLD#RHR1"1a&"RR0HMCsoC'NHloIC5HE802RR&"R7"&MRH0CCosl'HN5oCM_klODCD_U4.*U4.2RR&"RW"&MRH0CCosl'HN5oCI0H8ERR-.R*[-2R.R"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05lMk_DOCD._4U.*4URR+nRc,80CbER22&XR""RR&HCM0o'CsHolNCH5I8R0E-*R.[
2;RRRRRRRRRRRRLHCoMR
RRRRRRRRRR)RzqcvnRX:R)nqvc1X.RR
RRRRRRRRRRRRRRFRbsl0RN5bR7=4R>_R#HsM_CIo5HE80-[.*-,42RR7j=#>R__HMs5CoI0H8E*-.[2-.,jRqRR=>D_FINs885,j2RRq4=D>RFNI_858s4R2,q=.R>FRDI8_N8.s52R,
RRRRRRRRRRRRRRRRRRRRRRRRRRqd=D>RFNI_858sdR2,q=cR>FRDI8_N8cs52q,R6>R=RIDF_8N8s256,S
SSSSSR RWRR=>I_s0CnM_cW,RBRpi=B>RpRi,m=4R>kRF0k_L#c_n5lMk_DOCDc_n,8IH0.E-*4[-2m,Rj>R=R0Fk_#Lk_5ncM_klODCD_,ncI0H8E*-.[2-.2R;
RRRRRRRRRRRRR#RR_0Fk_osC58IH0.E-*4[-2=R<R0Fk_#Lk_5ncM_klODCD_,ncI0H8E*-.[2-4RCIEMFR5kC0_Mc_nR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRR_R#F_k0s5CoI0H8E*-.[2-.RR<=F_k0L_k#nMc5kOl_C_DDnIc,HE80-[.*-R.2IMECRk5F0M_C_Rnc=4R''C2RDR#C';Z'
RRRRRRRRMRC8CRoMNCs0zCR.
j;SCSRMo8RCsMCNR0Cz	OE_
.;SzSRO_E	4RR:H5VR#H_I8_0ENNss$c_n5Rj2>2RjRMoCC0sNCR
RRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqz)vRnc:NRDLRCDH"#R1"1aRH&RMo0CCHs'lCNo58IH0RE2&7R""RR&HCM0o'CsHolNCk5MlC_OD4D_.4U*.RU2&WR""RR&HCM0o'CsHolNCH5I8R0E-*R.#H_I8_0ENNss$c_n5R42-2R4R"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05lMk_DOCD._4U.*4URR+nRc,80CbER22&XR""RR&HCM0o'CsHolNCH5I8R0E-*R.#H_I8_0ENNss$c_n5242;R
RRRRRRRRRRCRLo
HMRRRRRRRRRRRRzv)qn:cRRv)qn4cX1RR
RRRRRRRRRRRRRbRRFRs0lRNb5=7R>_R#HsM_CIo5HE80-#.*_8IH0NE_s$sN_5nc442-2q,Rj>R=RIDF_8N8s25j,4RqRR=>D_FINs885,42RRq.=D>RFNI_858s.
2,RRRRRRRRRRRRRRRRRRRRRRRRRdRqRR=>D_FINs885,d2RRqc=D>RFNI_858scR2,q=6R>FRDI8_N86s52S,
SSSSSWRR >R=R0Is__CMnRc,WiBpRR=>B,piR=mR>kRF0k_L#c_n5lMk_DOCDc_n,8IH0.E-*I#_HE80_sNsNn$_c254-242;R
RRRRRRRRRRRRRR_R#F_k0s5CoI0H8E*-.#H_I8_0ENNss$c_n5-424<2R=kRF0k_L#c_n5lMk_DOCDc_n,8IH0.E-*I#_HE80_sNsNn$_c254-R42IMECRk5F0M_C_Rnc=4R''C2RDR#C';Z'
RRRRRRRRMRC8CRoMNCs0zCRO_E	4S;
RRRRR8CMRMoCC0sNC4Rz(R;RRRRRRRRR
R
RR-R-RMtCC0sNCRRN4InRFRs88bCCRv)qRDOCDVRHRbNbssFbHCN0RRRRRRRRRRRRR
RRRRRRzR.4:VRHRk5MlC_ODdD_.RR=4o2RCsMCN
0CRRRR-Q-RVNR58I8sHE80R6>R2CRMC08RFsROCCN0RHIs0CCRMDNLCMRN8kRF00bkRNCMLRDC#CCDOD0RFOoH
RRRRRRRR.z.NRR:H5VRNs88I0H8ERR>(MRN8kRMlC_ODnD_cRR=4o2RCsMCN
0CRRRRRRRRRRRRRRRRF_k0CdM_.=R<R''4RCIEM5R5#8_N_osC58N8s8IH04E-RI8FMR0F(=2RRlMk_DOCD._4UN2RM58R#8_N_osC5Rn2=4R''N2RM58R#8_N_osC5R62=jR''R22CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C_Rd.<W=R ERIC5MR5N#_8C_so85N8HsI8-0E4FR8IFM0RR(2=kRMlC_OD4D_.RU2NRM85N#_8C_so25nR'=R4R'2NRM85N#_8C_so256R'=Rj2'2R#CDCjR''R;
RRRRRCRRMo8RCsMCNR0CzN..;R
RRRRRR.Rz.:LRRRHV58N8s8IH0>ERRN(RMM8RkOl_C_DDn/cR=2R4RMoCC0sNCR
RRRRRRRRRRRRRRkRF0M_C_Rd.<'=R4I'RERCM5_5#Ns8_CNo58I8sHE80-84RF0IMF2R(RM=RkOl_C_DD42.UR8NMR_5#Ns8_Cno52RR='2j'R8NMR_5#Ns8_C6o52RR='2j'2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0CdM_.=R<RRW IMECR#55__N8s5CoNs88I0H8ER-48MFI0(FR2RR=M_klODCD_U4.2MRN8#R5__N8s5Con=2RR''j2MRN8#R5__N8s5Co6=2RR''j2C2RDR#C';j'
RRRRRRRR8CMRMoCC0sNC.Rz.
L;RRRRRRRRzO..RH:RVNR58I8sHE80R(=RR8NMRlMk_DOCDc_nR4=R2CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_M._dRR<='R4'IMECR#55__N8s5Con=2RR''42MRN8#R5__N8s5Co6=2RR''j2C2RDR#C';j'
RRRRRRRRRRRRRRRR0Is__CMd<.R= RWRCIEM5R5#8_N_osC5Rn2=4R''N2RM58R#8_N_osC5R62=jR''R22CCD#R''j;R
RRRRRRMRC8CRoMNCs0zCR.;.O
RRRRRRRR.z.8RR:H5VRNs88I0H8ERR=nMRN8kRMlC_ODnD_c=R/RR42oCCMsCN0
RRRRRRRRRRRRRRRR0Fk__CMd<.R=4R''ERIC5MR5N#_8C_so85N8HsI8-0E4FR8IFM0RR62=kRMlC_ODnD_cR22CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C_Rd.<W=R ERIC5MR5N#_8C_so85N8HsI8-0E4FR8IFM0RR62=kRMlC_ODnD_cR22CCD#R''j;R
RRRRRRMRC8CRoMNCs0zCR.;.8
RRRRR--Q5VRNs88I0H8E=R<RR62MIFRsCH0RNCMLRDCFFsRkk0b0MRCNCLDRD#CCRO0DHFoOCRMC88C
RRRRRRRRdz.RH:RVNR58I8sHE80RR<=6o2RCsMCN
0CRRRRRRRRRRRRRRRRF_k0CdM_.=R<R''4;R
RRRRRRRRRRRRRRsRI0M_C_Rd.<W=R R;
RRRRRCRRMo8RCsMCNR0Cz;.d
RRRRR--tCCMsCN0RC0ERv)qRDOCDMRN8sR0H0-#N
0CSRRRREzO	R_U:VRHR_5#I0H8Es_Ns5N$d>2RRRj2oCCMsCN0
zSSO_E	DRC6:VRHRH5I8R0E>U=R*I#_HE80_sNsNd$52MRN8HRI8R0E>U=R2CRoMNCs0RC
RRRRRRRRRRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)Rzq.vdRD:RNDLCRRH#"a11"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloMC5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*n2RR&"RW"&MRH0CCosl'HN5oCI0H8ERR-D_#LI0H8E&2RR"" RH&RMo0CCHs'lCNo50oC_8CM_b8C0ME5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*nRd+R.8,RCEb02&2RR""XRH&RMo0CCHs'lCNo58IH0-ERRLD#_8IH0+ERR;U2
RRRRRRRRRRRRRRRRRRRRoLCHSM
SRRRRqz)vRd.:)RXq.vdX
U1SRSSRbRRFRs0lRNb5=7R>NRb8_5#HsM_CIo5HE80-84RF0IMFHRI8-0ED_#LI0H8ER2,UD,R#IL_HE80-,42RRqj=D>RFNI_858sj
2,SSSSSRSRq=4R>FRDI8_N84s52q,R.>R=RIDF_8N8s25.,dRqRR=>D_FINs885,d2RRqc=D>RFNI_858scR2,W= R>sRI0M_C_,d.RpWBi>R=RiBp,S
SSSSSRRRm=0>RlUb__5d.j;22
SSSS#N#HRoM:FRVs[RHRRHMI0H8ER-48MFI0IFRHE80-LD#_8IH0oERCsMCN
0CSSSSRkRF0k_L#._d5lMk_DOCD._d,2H[RR<=0_lbU._d55j2HI[-HE80+LD#_8IH0;E2
RRRRRRRRRRRRRRRR#RR_0Fk_osC52H[RR<=F_k0L_k#dM.5kOl_C_DDdH.,[I2RERCM50Fk__CMd=.RR''42DRC#'CRZ
';SSSSCRM8oCCMsCN0R#N#H;oM
RRRRRRRRRRRRUz.RV:RF[sRRRHM#H_I8_0ENNss$25d-84RF0IMFRR4oCCMsCN0
RRRRRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)Rzq.vdRD:RNDLCRRH#"a11"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloMC5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*n2RR&"RW"&MRH0CCosl'HN5oCI0H8ERR-D_#LI0H8ERR-[2*UR"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05lMk_DOCD._4U.*4URR+M_klODCD_*ncn+cRR,d.Rb8C02E2R"&RX&"RR0HMCsoC'NHloIC5HE80RD-R#IL_HE80R5-R[2-4*;U2
RRRRRRRRRRRRLRRCMoH
RRRRRRRRRRRRzRR)dqv.RR:Xv)qdU.X1RR
RRRRRRRRRRRRRbRRFRs0lRNb5=7R>_R#HsM_CIo5HE80-LD#_8IH0UE-*([+RI8FMR0FI0H8E#-DLH_I8-0EU2*[,jRqRR=>D_FINs885,j2RRq4=D>RFNI_858s4R2,q=.R>FRDI8_N8.s52R,
RRRRRRRRRRRRRRRRRRRRRRRRRRqd=D>RFNI_858sdR2,q=cR>FRDI8_N8cs52W,R >R=R0Is__CMdR.,WiBpRR=>B,piR=mR>lR0b__Ud[.52
2;SRSSRNRR#o#HMRR:VRFsHH[RMRR(8MFI0jFRRMoCC0sNCS
SSRSRF_k0L_k#dM.5kOl_C_DDdI.,HE80-LD#_8IH0UE-*H[+[<2R=lR0b__Ud[.52[5H2R;
RRRRRRRRRRRRRRRRRF#_ks0_CIo5HE80-LD#_8IH0UE-*H[+[<2R=kRF0k_L#._d5lMk_DOCD._d,8IH0DE-#IL_HE80-[U*+2H[RCIEMFR5kC0_M._dR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRMRC8CRoMNCs0NCR#o#HMR;
RRRRRRRRRCRRMo8RCsMCNR0Cz;.U
CSSMo8RCsMCNR0Cz	OE_6DC;S
Sz	OE_6o0RH:RVIR5HE80RR>=UMRN8HRI8R0ElRF8U=R>RR62oCCMsCN0
RRRRRRRRRRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVzv)qd:.RRLDNCHDR#1R"1Ra"&MRH0CCosl'HN5oCI0H8E&2RR""7RH&RMo0CCHs'lCNo5lMk_DOCD._4U.*4URR+M_klODCD_*ncnRc2&WR""RR&HCM0o'CsHolNCH5I8R0E-#RDLH_I820ER"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05lMk_DOCD._4U.*4URR+M_klODCD_*ncn+cRR,d.Rb8C02E2R"&RX&"RR0HMCsoC'NHloIC5HE80RD-R#IL_HE80RU+R2R;
RRRRRRRRRRRRRRRRRLRRCMoH
RSSRzRR)dqv.RR:Xv)qdU.X1S
SSRRRRsbF0NRlb7R5RR=>b5N8#M_H_osC58IH04E-RI8FMR0FI0H8E#-DLH_I820E,,RURLD#_8IH04E-2q,Rj>R=RIDF_8N8s25j,S
SSSSSR4RqRR=>D_FINs885,42RRq.=D>RFNI_858s.R2,q=dR>FRDI8_N8ds52q,Rc>R=RIDF_8N8s25c, RWRR=>I_s0CdM_.W,RBRpi=B>Rp
i,SSSSSRSRm>R=Rb0l_dU_._5#I0H8Es_Ns5N$d42-2
2;SSSSNH##o:MRRsVFRRH[HIMRHE80-84RF0IMFHRI8-0ED_#LI0H8ECRoMNCs0SC
SRSSR0Fk_#Lk_5d.M_klODCD_,d.HR[2<0=RlUb__5d.#H_I8_0ENNss$25d-542HI[-HE80+LD#_8IH0;E2
RRRRRRRRRRRRRRRR#RR_0Fk_osC52H[RR<=F_k0L_k#dM.5kOl_C_DDdH.,[I2RERCM50Fk__CMd=.RR''42DRC#'CRZ
';SSSSCRM8oCCMsCN0R#N#H;oM
RRRRRRRRRRRRUz.RV:RF[sRRRHM#H_I8_0ENNss$25d-8.RF0IMFRRjoCCMsCN0
RRRRRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)Rzq.vdRD:RNDLCRRH#"a11"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloMC5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*n2RR&"RW"&MRH0CCosl'HN5oC[2*UR"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05lMk_DOCD._4U.*4URR+M_klODCD_*ncn+cRR,d.Rb8C02E2R"&RX&"RR0HMCsoC'NHlo5C5[2+4*;U2
RRRRRRRRRRRRLRRCMoH
RRRRRRRRRRRRzRR)dqv.RR:Xv)qdU.X1RR
RRRRRRRRRRRRRbRRFRs0lRNb5=7R>_R#HsM_CUo5*([+RI8FMR0FU2*[,jRqRR=>D_FINs885,j2RRq4=D>RFNI_858s4R2,q=.R>FRDI8_N8.s52R,
RRRRRRRRRRRRRRRRRRRRRRRRRRqd=D>RFNI_858sdR2,q=cR>FRDI8_N8cs52W,R >R=R0Is__CMdR.,WiBpRR=>B,piR=mR>lR0b__Ud[.52
2;SSSSNH##o:MRRsVFRRH[H(MRRI8FMR0FjCRoMNCs0SC
SRSSR0Fk_#Lk_5d.M_klODCD_,d.U+*[HR[2<0=RlUb__5d.[H25[
2;RRRRRRRRRRRRRRRRR_R#F_k0s5CoU+*[HR[2<F=RkL0_kd#_.k5MlC_ODdD_.*,U[[+H2ERIC5MRF_k0CdM_.RR='24'R#CDCZR''R;
RRRRRRRRRRRRRCRRMo8RCsMCNR0CNH##o
M;RRRRRRRRRRRRCRM8oCCMsCN0RUz.;S
SCRM8oCCMsCN0REzO	0_o6S;
SEzO	R_M:VRHRH5I8R0E<2RURMoCC0sNCR
RRRRRRRRRRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqz)vRd.:NRDLRCDH"#R1"1aRH&RMo0CCHs'lCNo58IH0RE2&7R""RR&HCM0o'CsHolNCk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*2ncR"&RW&"RR0HMCsoC'NHlojC52RR&"R "&MRH0CCosl'HN5oCo_C0C_M880CbEk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*Rnc+.Rd,CR8b20E2RR&"RX"&MRH0CCosl'HN5oCU
2;RRRRRRRRRRRRRRRRRRRRLHCoMS
SRRRRzv)qd:.RRqX)vXd.US1
SRSRRFRbsl0RN5bR7>R=R8bN5H#_MC_soH5I8-0E4FR8IFM0R8IH0DE-#IL_HE802U,R,#RDLH_I8-0E4R2,q=jR>FRDI8_N8js52S,
SSSSSqRR4>R=RIDF_8N8s254,.RqRR=>D_FINs885,.2RRqd=D>RFNI_858sdR2,q=cR>FRDI8_N8cs52W,R >R=R0Is__CMdR.,WiBpRR=>B,pi
SSSSRSSR=mR>lR0b__Udj.52
2;SSSSNH##o:MRRsVFRRH[HIMRHE80-84RF0IMFRRjoCCMsCN0
SSSSFRRkL0_kd#_.k5MlC_ODdD_.[,H2=R<Rb0l_dU_.25j52H[;R
RRRRRRRRRRRRRRRRR#k_F0C_so[5H2=R<R0Fk_#Lk_5d.M_klODCD_,d.HR[2IMECRk5F0M_C_Rd.=4R''C2RDR#C';Z'
SSSS8CMRMoCC0sNC#RN#MHo;S
SCRM8oCCMsCN0REzO	;_M
CSSMo8RCsMCNR0Cz	OE_
U;SOSzEc	_RH:RV#R5_8IH0NE_s$sN5R.2>2RjRMoCC0sNCR
RRRRRR.RzcR_c:VRHRH5I8R0E>c=R2CRoMNCs0RC
RRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)Rzq.vdRD:RNDLCRRH#"a11"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloMC5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*n2RR&"RW"&MRH0CCosl'HN5oCj&2RR"" RH&RMo0CCHs'lCNo50oC_8CM_b8C0ME5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*nRd+R.8,RCEb02&2RR""XRH&RMo0CCHs'lCNo5;c2
RRRRRRRRRRRRoLCHRM
RRRRRRRRRzRR)dqv.RR:Xv)qdc.X1RR
RRRRRRRRRRRRRbRRFRs0lRNb5R7d=#>R__HMs5CodR2,7=.R>_R#HsM_C.o527,R4>R=RH#_MC_so254,jR7RR=>#M_H_osC5,j2
SSSRRRRRRRRRRRRRjRqRR=>D_FINs885,j2RRq4=D>RFNI_858s4R2,q=.R>FRDI8_N8.s52R,
RRRRRRRRRRRRRRRRRRRRRRRRRRqd=D>RFNI_858sdR2,q=cR>FRDI8_N8cs52W,R >R=R0Is__CMdR.,WiBpRR=>B,piRS
SSSSSRdRmRR=>F_k0L_k#dM.5kOl_C_DDdd.,2m,R.>R=R0Fk_#Lk_5d.M_klODCD_,d..
2,SSSSSRSRm=4R>kRF0k_L#._d5lMk_DOCD._d,,42RRmj=F>RkL0_kd#_.k5MlC_ODdD_.2,j2R;
RRRRRRRRRRRRR#RR_0Fk_osC5Rd2<F=RkL0_kd#_.k5MlC_ODdD_.2,dRCIEMFR5kC0_M._dR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRR_R#F_k0s5Co.<2R=kRF0k_L#._d5lMk_DOCD._d,R.2IMECRk5F0M_C_Rd.=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRF#_ks0_C4o52=R<R0Fk_#Lk_5d.M_klODCD_,d.4I2RERCM50Fk__CMd=.RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRR#k_F0C_so25jRR<=F_k0L_k#dM.5kOl_C_DDdj.,2ERIC5MRF_k0CdM_.RR='24'R#CDCZR''R;
RRRRRCRRMo8RCsMCNR0Cz_.ccR;
RRRRRzRR.dc_RH:RVIR5HE80Rd=R2CRoMNCs0RC
RRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)Rzq.vdRD:RNDLCRRH#"a11"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloMC5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*n2RR&"RW"&MRH0CCosl'HN5oCj&2RR"" RH&RMo0CCHs'lCNo50oC_8CM_b8C0ME5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*nRd+R.8,RCEb02&2RR""XRH&RMo0CCHs'lCNo5;c2
RRRRRRRRRRRRoLCHRM
RRRRRRRRRzRR)dqv.RR:Xv)qdc.X1RR
RRRRRRRRRRRRRbRRFRs0lRNb5R7d='>RjR',7=.R>_R#HsM_C.o527,R4>R=RH#_MC_so254,jR7RR=>#M_H_osC5,j2
SSSRRRRRRRRRRRRRjRqRR=>D_FINs885,j2RRq4=D>RFNI_858s4R2,q=.R>FRDI8_N8.s52R,
RRRRRRRRRRRRRRRRRRRRRRRRRRqd=D>RFNI_858sdR2,q=cR>FRDI8_N8cs52W,R >R=R0Is__CMdR.,WiBpRR=>B,piRS
SSSSSRdRmRR=>FMbC,.RmRR=>F_k0L_k#dM.5kOl_C_DDd..,2S,
SSSSSmRR4>R=R0Fk_#Lk_5d.M_klODCD_,d.4R2,m=jR>kRF0k_L#._d5lMk_DOCD._d,2j2;R
RRRRRRRRRRRRRR_R#F_k0s5Co.<2R=kRF0k_L#._d5lMk_DOCD._d,R.2IMECRk5F0M_C_Rd.=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRF#_ks0_C4o52=R<R0Fk_#Lk_5d.M_klODCD_,d.4I2RERCM50Fk__CMd=.RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRR#k_F0C_so25jRR<=F_k0L_k#dM.5kOl_C_DDdj.,2ERIC5MRF_k0CdM_.RR='24'R#CDCZR''R;
RRRRRCRRMo8RCsMCNR0Cz_.cdS;
S8CMRMoCC0sNCORzEc	_;S
Sz	OE_:.RRRHV5I#_HE80_sNsN4$52RR>jo2RCsMCN
0CRRRRRRRRzR.c:FRVsRR[H5MR#H_I8_0ENNss$254R4-R2FR8IFM0RojRCsMCN
0CRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FzVR)dqv.RR:DCNLD#RHR1"1a&"RR0HMCsoC'NHloIC5HE802RR&"R7"&MRH0CCosl'HN5oCM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*c&2RR""WRH&RMo0CCHs'lCNo58IH0UE-*I#_HE80_sNsNd$52*-.[2-.R"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05lMk_DOCD._4U.*4URR+M_klODCD_*ncn+cRR,d.Rb8C02E2R"&RX&"RR0HMCsoC'NHloIC5HE80-#U*_8IH0NE_s$sN5-d2.2*[;R
RRRRRRRRRRCRLo
HMRRRRRRRRRRRRzv)qd:.RRv)qd..X1RR
RRRRRRRRRRRRRbRRFRs0lRNb5R7j=#>R__HMs5CoI0H8E*-U#H_I8_0ENNss$25d-[.*-,.2RR74=#>R__HMs5CoI0H8E*-U#H_I8_0ENNss$25d-[.*-,42RRqj=D>RFNI_858sjR2,q=4R>FRDI8_N84s52q,R.>R=RIDF_8N8s25.,R
RRRRRRRRRRRRRRRRRRRRRRRRRq=dR>FRDI8_N8ds52q,Rc>R=RIDF_8N8s25c, RWRR=>I_s0CdM_.W,RBRpi=B>RpRi,m=jR>kRF0k_L#._d5lMk_DOCD._d,8IH0UE-*I#_HE80_sNsNd$52*-.[2-.,S
SSSSSR4RmRR=>F_k0L_k#dM.5kOl_C_DDdI.,HE80-#U*_8IH0NE_s$sN5-d2.-*[4;22
RRRRRRRRRRRRRRRRF#_ks0_CIo5HE80-#U*_8IH0NE_s$sN5-d2.-*[4<2R=kRF0k_L#._d5lMk_DOCD._d,8IH0UE-*I#_HE80_sNsNd$52*-.[2-4RCIEMFR5kC0_M._dR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRR_R#F_k0s5CoI0H8E*-U#H_I8_0ENNss$25d-[.*-R.2<F=RkL0_kd#_.k5MlC_ODdD_.H,I8-0EU_*#I0H8Es_Ns5N$d.2-*.[-2ERIC5MRF_k0CdM_.RR='24'R#CDCZR''R;
RRRRRCRRMo8RCsMCNR0Cz;.c
CSSMo8RCsMCNR0Cz	OE_
.;SOSzE4	_RH:RV#R5_8IH0NE_s$sN5Rj2>2RjRMoCC0sNCR
RRRRRR.RzcRR:H5VRI0H8EFRl8RRU=2R4RMoCC0sNCR
RRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqz)vRd.:NRDLRCDH"#R1"1aRH&RMo0CCHs'lCNo58IH0RE2&7R""RR&HCM0o'CsHolNCk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*2ncR"&RW&"RR0HMCsoC'NHlojC52RR&"R "&MRH0CCosl'HN5oCo_C0C_M880CbEk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*Rnc+.Rd,CR8b20E2RR&"RX"&MRH0CCosl'HN5oC4
2;RRRRRRRRRRRRLHCoMR
RRRRRRRRRR)Rzq.vdR):Rq.vdXR41
RRRRRRRRRRRRRRRRsbF0NRlb7R5RR=>#M_H_osC5,j2RRqj=D>RFNI_858sjR2,q=4R>FRDI8_N84s52q,R.>R=RIDF_8N8s25.,R
RRRRRRRRRRRRRRRRRRRRRRRRRq=dR>FRDI8_N8ds52q,Rc>R=RIDF_8N8s25c, RWRR=>I_s0CdM_.W,RBRpi=B>RpRi,m>R=R0Fk_#Lk_5d.M_klODCD_,d.j;22
RRRRRRRRRRRRRRRRF#_ks0_Cjo52=R<R0Fk_#Lk_5d.M_klODCD_,d.jI2RERCM50Fk__CMd=.RR''42DRC#'CRZ
';RRRRRRRRCRM8oCCMsCN0Rcz.;S
SCRM8oCCMsCN0REzO	;_4
RRRR8CMRMoCC0sNC.Rz4R;RRRRRRRRR
R
RR-R-RMtCC0sNCRRN4InRFRs88bCCRv)qRDOCDVRHRbNbssFbHCN0RRRRRRRRRRRRR
RRRRRRzR.6:VRHRk5MlC_OD4D_nRR=4o2RCsMCN
0CRRRR-Q-RVNR58I8sHE80R6>R2CRMC08RFsROCCN0RHIs0CCRMDNLCMRN8kRF00bkRNCMLRDC#CCDOD0RFOoH
RRRRRRRRnz.NRR:H5VRNs88I0H8ERR>(MRN8kRMlC_ODnD_cRR=4MRN8kRMlC_ODdD_.RR=4o2RCsMCN
0CRRRRRRRRRRRRRRRRF_k0C4M_n=R<R''4RCIEM5R5#8_N_osC58N8s8IH04E-RI8FMR0F(=2RRlMk_DOCD._4UN2RM58R#8_N_osC5Rn2=4R''N2RM58R#8_N_osC5R62=4R''N2RM58R#8_N_osC5Rc2=jR''R22CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C_R4n<W=R ERIC5MR5N#_8C_so85N8HsI8-0E4FR8IFM0RR(2=kRMlC_OD4D_.RU2NRM85N#_8C_so25nR'=R4R'2NRM85N#_8C_so256R'=R4R'2NRM85N#_8C_so25cR'=Rj2'2R#CDCjR''R;
RRRRRCRRMo8RCsMCNR0CzN.n;R
RRRRRR.Rzn:LRRRHV58N8s8IH0>ERRN(RMM8RkOl_C_DDn=cRRN4RMM8RkOl_C_DDd=.RRRj2oCCMsCN0
RRRRRRRRRRRRRRRR0Fk__CM4<nR=4R''ERIC5MR5N#_8C_so85N8HsI8-0E4FR8IFM0RR(2=kRMlC_OD4D_.RU2NRM85N#_8C_so25nR'=R4R'2NRM85N#_8C_so256R'=RjR'2NRM85N#_8C_so25cR'=Rj2'2R#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_Mn_4RR<=WI RERCM5_5#Ns8_CNo58I8sHE80-84RF0IMF2R(RM=RkOl_C_DD42.UR8NMR_5#Ns8_Cno52RR='24'R8NMR_5#Ns8_C6o52RR='2j'R8NMR_5#Ns8_Cco52RR='2j'2DRC#'CRj
';RRRRRRRRCRM8oCCMsCN0Rnz.LR;
RRRRRzRR.RnO:VRHR85N8HsI8R0E>RR(NRM8M_klODCD_Rnc=RRjNRM8M_klODCD_Rd.=2R4RMoCC0sNCR
RRRRRRRRRRRRRRkRF0M_C_R4n<'=R4I'RERCM5_5#Ns8_CNo58I8sHE80-84RF0IMF2R(RM=RkOl_C_DD42.UR8NMR_5#Ns8_Cno52RR='2j'R8NMR_5#Ns8_C6o52RR='24'R8NMR_5#Ns8_Cco52RR='2j'2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0C4M_n=R<RRW IMECR#55__N8s5CoNs88I0H8ER-48MFI0(FR2RR=M_klODCD_U4.2MRN8#R5__N8s5Con=2RR''j2MRN8#R5__N8s5Co6=2RR''42MRN8#R5__N8s5Coc=2RR''j2C2RDR#C';j'
RRRRRRRR8CMRMoCC0sNC.Rzn
O;RRRRRRRRz8.nRH:RVNR58I8sHE80R(>RR8NMRlMk_DOCDc_nRj=RR8NMRlMk_DOCD._dRj=R2CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_Mn_4RR<='R4'IMECR#55__N8s5CoNs88I0H8ER-48MFI0(FR2RR=M_klODCD_U4.2MRN8#R5__N8s5Con=2RR''j2MRN8#R5__N8s5Co6=2RR''j2MRN8#R5__N8s5Coc=2RR''j2C2RDR#C';j'
RRRRRRRRRRRRRRRR0Is__CM4<nR= RWRCIEM5R5#8_N_osC58N8s8IH04E-RI8FMR0F(=2RRlMk_DOCD._4UN2RM58R#8_N_osC5Rn2=jR''N2RM58R#8_N_osC5R62=jR''N2RM58R#8_N_osC5Rc2=jR''R22CCD#R''j;R
RRRRRRMRC8CRoMNCs0zCR.;n8
RRRRRRRRnz.CRR:H5VRNs88I0H8ERR=(MRN8kRMlC_ODnD_cRR=4MRN8kRMlC_ODdD_.RR=4o2RCsMCN
0CRRRRRRRRRRRRRRRRF_k0C4M_n=R<R''4RCIEM5R5#8_N_osC5Rn2=4R''N2RM58R#8_N_osC5R62=4R''N2RM58R#8_N_osC5Rc2=jR''R22CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C_R4n<W=R ERIC5MR5N#_8C_so25nR'=R4R'2NRM85N#_8C_so256R'=R4R'2NRM8R_5#Ns8_Cco52RR='2j'2DRC#'CRj
';RRRRRRRRCRM8oCCMsCN0Rnz.CR;
RRRRRzRR.RnV:VRHR85N8HsI8R0E=RR(NRM8M_klODCD_Rnc=RR4NRM8M_klODCD_Rd.=2RjRMoCC0sNCR
RRRRRRRRRRRRRRkRF0M_C_R4n<'=R4I'RERCM5_5#Ns8_Cno52RR='24'R8NMR_5#Ns8_C6o52RR='2j'R8NMR_5#Ns8_Cco52RR='2j'2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0C4M_n=R<RRW IMECR#55__N8s5Con=2RR''42MRN8#R5__N8s5Co6=2RR''j2MRN8#R5__N8s5Coc=2RR''j2C2RDR#C';j'
RRRRRRRR8CMRMoCC0sNC.Rzn
V;RRRRRRRRzo.nRH:RVNR58I8sHE80Rn=RR8NMRlMk_DOCDc_nRj=RR8NMRlMk_DOCD._dR4=R2CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_Mn_4RR<='R4'IMECR#55__N8s5Co6=2RR''42MRN8#R5__N8s5Coc=2RR''j2C2RDR#C';j'
RRRRRRRRRRRRRRRR0Is__CM4<nR= RWRCIEM5R5#8_N_osC5R62=4R''N2RM58R#8_N_osC5Rc2=jR''R22CCD#R''j;R
RRRRRRMRC8CRoMNCs0zCR.;no
RRRRRRRRnz.ERR:H5VRNs88I0H8ERR=6MRN8kRMlC_ODdD_.=R/RR42oCCMsCN0
RRRRRRRRRRRRRRRR0Fk__CM4<nR=4R''ERIC5MR5N#_8C_so85N8HsI8-0E4FR8IFM0RRc2=kRMlC_ODdD_.R22CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C_R4n<W=R ERIC5MR5N#_8C_so85N8HsI8-0E4FR8IFM0RRc2=kRMlC_ODdD_.R22CCD#R''j;R
RRRRRRMRC8CRoMNCs0zCR.;nE
RRRRR--Q5VRNs88I0H8E=R<RR62MIFRsCH0RNCMLRDCFFsRkk0b0MRCNCLDRD#CCRO0DHFoOCRMC88C
RRRRRRRR(z.RH:RVNR58I8sHE80RR<=co2RCsMCN
0CRRRRRRRRRRRRRRRRF_k0C4M_n=R<R''4;R
RRRRRRRRRRRRRRsRI0M_C_R4n<W=R R;
RRRRRCRRMo8RCsMCNR0Cz;.(
RRRRR--tCCMsCN0RC0ERv)qRDOCDMRN8sR0H0-#N
0CSRRRREzO	R_U:VRHR_5#I0H8Es_Ns5N$d>2RRRj2oCCMsCN0
zSSO_E	DRC6:VRHRH5I8R0E>U=R*I#_HE80_sNsNd$52MRN8HRI8R0E>U=R2CRoMNCs0RC
RRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)Rzqnv4RD:RNDLCRRH#"a11"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloMC5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*nRM+RkOl_C_DDdd.*.&2RR""WRH&RMo0CCHs'lCNo58IH0-ERRLD#_8IH0RE2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50EM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*cRR+M_klODCD_*d.d+.RR,4nRb8C02E2R"&RX&"RR0HMCsoC'NHloIC5HE80RD-R#IL_HE80RU+R2R;
RRRRRRRRRLRRCMoH
RSSRzRR)4qvnRR:Xv)q4UnX1S
SSRRRRsbF0NRlb7R5RR=>b5N8#M_H_osC58IH04E-RI8FMR0FI0H8E#-DLH_I820E,,RURLD#_8IH04E-2q,Rj>R=RIDF_8N8s25j,S
SSSSSR4RqRR=>D_FINs885,42RRq.=D>RFNI_858s.R2,q=dR>FRDI8_N8ds52W,R >R=R0Is__CM4Rn,WiBpRR=>B,pi
SSSSRSSR=mR>lR0b__U4jn52
2;SSSSNH##o:MRRsVFRRH[HIMRHE80-84RF0IMFHRI8-0ED_#LI0H8ECRoMNCs0SC
SRSSR0Fk_#Lk_54nM_klODCD_,4nHR[2<0=RlUb__54njH25[H-I8+0ED_#LI0H8E
2;RRRRRRRRRRRRRRRRR_R#F_k0s5CoHR[2<F=RkL0_k4#_nk5MlC_OD4D_n[,H2ERIC5MRF_k0C4M_nRR='24'R#CDCZR''S;
SCSSMo8RCsMCNR0CNH##o
M;RRRRRRRRRRRRzR.U:FRVsRR[H#MR_8IH0NE_s$sN5-d24FR8IFM0Ro4RCsMCN
0CRRRRRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqz)vR4n:NRDLRCDH"#R1"1aRH&RMo0CCHs'lCNo58IH0RE2&7R""RR&HCM0o'CsHolNCk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*Rnc+kRMlC_ODdD_..*d2RR&"RW"&MRH0CCosl'HN5oCI0H8ERR-D_#LI0H8ERR-[2*UR"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05lMk_DOCD._4U.*4URR+M_klODCD_*ncn+cRRlMk_DOCD._d*Rd.+nR4,CR8b20E2RR&"RX"&MRH0CCosl'HN5oCI0H8ERR-D_#LI0H8ERR-54[-22*U;R
RRRRRRRRRRRRRLHCoMR
RRRRRRRRRRRRRzv)q4:nRRqX)vX4nU
1RRRRRRRRRRRRRRRRRb0FsRblNRR57=#>R__HMs5CoI0H8E#-DLH_I8-0EU+*[(FR8IFM0R8IH0DE-#IL_HE80-[U*2q,Rj>R=RIDF_8N8s25j,4RqRR=>D_FINs885,42RRq.=D>RFNI_858s.
2,RRRRRRRRRRRRRRRRRRRRRRRRRdRqRR=>D_FINs885,d2RRW =I>RsC0_Mn_4,BRWp=iR>pRBim,RRR=>0_lbUn_452[2;S
SSRRRR#N#HRoM:FRVs[RHRRHM(FR8IFM0RojRCsMCN
0CSSSSRkRF0k_L#n_45lMk_DOCDn_4,8IH0DE-#IL_HE80-[U*+2H[RR<=0_lbUn_455[2H;[2
RRRRRRRRRRRRRRRR#RR_0Fk_osC58IH0DE-#IL_HE80-[U*+2H[RR<=F_k0L_k#4Mn5kOl_C_DD4In,HE80-LD#_8IH0UE-*H[+[I2RERCM50Fk__CM4=nRR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRCRM8oCCMsCN0R#N#H;oM
RRRRRRRRRRRR8CMRMoCC0sNC.RzUS;
S8CMRMoCC0sNCORzED	_C
6;SOSzEo	_0:6RRRHV58IH0>ER=RRUNRM8I0H8EFRl8RRU>6=R2CRoMNCs0RC
RRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)Rzqnv4RD:RNDLCRRH#"a11"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloMC5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*nRM+RkOl_C_DDdd.*.&2RR""WRH&RMo0CCHs'lCNo58IH0-ERRLD#_8IH0RE2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50EM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*cRR+M_klODCD_*d.d+.RR,4nRb8C02E2R"&RX&"RR0HMCsoC'NHloIC5HE80RD-R#IL_HE80RU+R2R;
RRRRRRRRRLRRCMoH
RSSRzRR)4qvnRR:Xv)q4UnX1S
SSRRRRsbF0NRlb7R5RR=>b5N8#M_H_osC58IH04E-RI8FMR0FI0H8E#-DLH_I820E,,RURLD#_8IH04E-2q,Rj>R=RIDF_8N8s25j,S
SSSSSR4RqRR=>D_FINs885,42RRq.=D>RFNI_858s.R2,q=dR>FRDI8_N8ds52W,R >R=R0Is__CM4Rn,WiBpRR=>B,pi
SSSSRSSR=mR>lR0b__U4#n5_8IH0NE_s$sN5-d24;22
SSSS#N#HRoM:FRVs[RHRRHMI0H8ER-48MFI0IFRHE80-LD#_8IH0oERCsMCN
0CSSSSRkRF0k_L#n_45lMk_DOCDn_4,2H[RR<=0_lbUn_45I#_HE80_sNsNd$522-45-H[I0H8E#+DLH_I820E;R
RRRRRRRRRRRRRRRRR#k_F0C_so[5H2=R<R0Fk_#Lk_54nM_klODCD_,4nHR[2IMECRk5F0M_C_R4n=4R''C2RDR#C';Z'
SSSS8CMRMoCC0sNC#RN#MHo;R
RRRRRRRRRR.RzURR:VRFs[MRHRI#_HE80_sNsNd$52R-.8MFI0jFRRMoCC0sNCR
RRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FzVR)4qvnRR:DCNLD#RHR1"1a&"RR0HMCsoC'NHloIC5HE802RR&"R7"&MRH0CCosl'HN5oCM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*cRR+M_klODCD_*d.dR.2&WR""RR&HCM0o'CsHolNC*5[U&2RR"" RH&RMo0CCHs'lCNo50oC_8CM_b8C0ME5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*nRM+RkOl_C_DDdd.*.RR+4Rn,80CbER22&XR""RR&HCM0o'CsHolNC[55+*42U
2;RRRRRRRRRRRRRCRLo
HMRRRRRRRRRRRRR)Rzqnv4RX:R)4qvn1XURR
RRRRRRRRRRRRRRFRbsl0RN5bR7>R=RH#_MC_so*5U[R+(8MFI0UFR*,[2RRqj=D>RFNI_858sjR2,q=4R>FRDI8_N84s52q,R.>R=RIDF_8N8s25.,R
RRRRRRRRRRRRRRRRRRRRRRRRRq=dR>FRDI8_N8ds52W,R >R=R0Is__CM4Rn,WiBpRR=>B,piR=mR>lR0b__U4[n52
2;SSSSNH##o:MRRsVFRRH[H(MRRI8FMR0FjCRoMNCs0SC
SRSSR0Fk_#Lk_54nM_klODCD_,4nU+*[HR[2<0=RlUb__54n[H25[
2;RRRRRRRRRRRRRRRRR_R#F_k0s5CoU+*[HR[2<F=RkL0_k4#_nk5MlC_OD4D_n*,U[[+H2ERIC5MRF_k0C4M_nRR='24'R#CDCZR''R;
RRRRRRRRRRRRRCRRMo8RCsMCNR0CNH##o
M;RRRRRRRRRRRRCRM8oCCMsCN0RUz.;S
SCRM8oCCMsCN0REzO	0_o6S;
SEzO	R_M:VRHRH5I8R0E<2RURMoCC0sNCR
RRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqz)vR4n:NRDLRCDH"#R1"1aRH&RMo0CCHs'lCNo58IH0RE2&7R""RR&HCM0o'CsHolNCk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*Rnc+kRMlC_ODdD_..*d2RR&"RW"&MRH0CCosl'HN5oCj&2RR"" RH&RMo0CCHs'lCNo50oC_8CM_b8C0ME5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*nRM+RkOl_C_DDdd.*.RR+4Rn,80CbER22&XR""RR&HCM0o'CsHolNC25U;R
RRRRRRRRRRCRLo
HMSRSRR)Rzqnv4RX:R)4qvn1XU
SSSRRRRb0FsRblNRR57=b>RN#85__HMs5CoI0H8ER-48MFI0IFRHE80-LD#_8IH0,E2RRU,D_#LI0H8E2-4,jRqRR=>D_FINs885,j2
SSSSRSSRRq4=D>RFNI_858s4R2,q=.R>FRDI8_N8.s52q,Rd>R=RIDF_8N8s25d, RWRR=>I_s0C4M_nW,RBRpi=B>Rp
i,SSSSSRSRm>R=Rb0l_4U_n25j2S;
SNSS#o#HMRR:VRFsHH[RMHRI8-0E4FR8IFM0RojRCsMCN
0CSSSSRkRF0k_L#n_45lMk_DOCDn_4,2H[RR<=0_lbUn_455j2H;[2
RRRRRRRRRRRRRRRR#RR_0Fk_osC52H[RR<=F_k0L_k#4Mn5kOl_C_DD4Hn,[I2RERCM50Fk__CM4=nRR''42DRC#'CRZ
';SSSSCRM8oCCMsCN0R#N#H;oM
CSSMo8RCsMCNR0Cz	OE_
M;SMSC8CRoMNCs0zCRO_E	US;
SEzO	R_c:VRHR_5#I0H8Es_Ns5N$.>2RRRj2oCCMsCN0
RRRRRRRRgz._:cRRRHV58IH0>ER=2RcRMoCC0sNCR
RRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqz)vR4n:NRDLRCDH"#R1"1aRH&RMo0CCHs'lCNo58IH0RE2&7R""RR&HCM0o'CsHolNCk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*Rnc+kRMlC_ODdD_..*d2RR&"RW"&MRH0CCosl'HN5oCj&2RR"" RH&RMo0CCHs'lCNo50oC_8CM_b8C0ME5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*nRM+RkOl_C_DDdd.*.RR+4Rn,80CbER22&XR""RR&HCM0o'CsHolNC25c;R
RRRRRRRRRRCRLo
HMRRRRRRRRRRRRzv)q4:nRRv)q4cnX1RR
RRRRRRRRRRRRRbRRFRs0lRNb5R7d=#>R__HMs5CodR2,7=.R>_R#HsM_C.o527,R4>R=RH#_MC_so254,jR7RR=>#M_H_osC5,j2
SSSRRRRRRRRRRRRRjRqRR=>D_FINs885,j2RRq4=D>RFNI_858s4R2,q=.R>FRDI8_N8.s52R,
RRRRRRRRRRRRRRRRRRRRRRRRRRqd=D>RFNI_858sdR2,W= R>sRI0M_C_,4nRpWBi>R=RiBp,SR
SSSSSmRRd>R=R0Fk_#Lk_54nM_klODCD_,4ndR2,m=.R>kRF0k_L#n_45lMk_DOCDn_4,,.2
SSSSRSSRRm4=F>RkL0_k4#_nk5MlC_OD4D_n2,4,jRmRR=>F_k0L_k#4Mn5kOl_C_DD4jn,2
2;RRRRRRRRRRRRRRRR#k_F0C_so25dRR<=F_k0L_k#4Mn5kOl_C_DD4dn,2ERIC5MRF_k0C4M_nRR='24'R#CDCZR''R;
RRRRRRRRRRRRR#RR_0Fk_osC5R.2<F=RkL0_k4#_nk5MlC_OD4D_n2,.RCIEMFR5kC0_Mn_4R'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRR_R#F_k0s5Co4<2R=kRF0k_L#n_45lMk_DOCDn_4,R42IMECRk5F0M_C_R4n=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRF#_ks0_Cjo52=R<R0Fk_#Lk_54nM_klODCD_,4njI2RERCM50Fk__CM4=nRR''42DRC#'CRZ
';RRRRRRRRCRM8oCCMsCN0Rgz._
c;RRRRRRRRz_.gdRR:H5VRI0H8ERR=do2RCsMCN
0CRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FzVR)4qvnRR:DCNLD#RHR1"1a&"RR0HMCsoC'NHloIC5HE802RR&"R7"&MRH0CCosl'HN5oCM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*cRR+M_klODCD_*d.dR.2&WR""RR&HCM0o'CsHolNC25jR"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05lMk_DOCD._4U.*4URR+M_klODCD_*ncn+cRRlMk_DOCD._d*Rd.+nR4,CR8b20E2RR&"RX"&MRH0CCosl'HN5oCc
2;RRRRRRRRRRRRLHCoMR
RRRRRRRRRR)Rzqnv4R):Rqnv4XRc1
RRRRRRRRRRRRRRRRsbF0NRlb7R5d>R=R''j,.R7RR=>#M_H_osC5,.2RR74=#>R__HMs5Co4R2,7=jR>_R#HsM_Cjo52S,
SRSRRRRRRRRRRRRRq=jR>FRDI8_N8js52q,R4>R=RIDF_8N8s254,.RqRR=>D_FINs885,.2
RRRRRRRRRRRRRRRRRRRRRRRRqRRd>R=RIDF_8N8s25d, RWRR=>I_s0C4M_nW,RBRpi=B>RpRi,
SSSSRSSRRmd=F>Rb,CMRRm.=F>RkL0_k4#_nk5MlC_OD4D_n2,.,S
SSSSSR4RmRR=>F_k0L_k#4Mn5kOl_C_DD44n,2m,Rj>R=R0Fk_#Lk_54nM_klODCD_,4nj;22
RRRRRRRRRRRRRRRRF#_ks0_C.o52=R<R0Fk_#Lk_54nM_klODCD_,4n.I2RERCM50Fk__CM4=nRR''42DRC#'CRZ
';RRRRRRRRRRRRRRRR#k_F0C_so254RR<=F_k0L_k#4Mn5kOl_C_DD44n,2ERIC5MRF_k0C4M_nRR='24'R#CDCZR''R;
RRRRRRRRRRRRR#RR_0Fk_osC5Rj2<F=RkL0_k4#_nk5MlC_OD4D_n2,jRCIEMFR5kC0_Mn_4R'=R4R'2CCD#R''Z;R
RRRRRRMRC8CRoMNCs0zCR.dg_;S
SCRM8oCCMsCN0REzO	;_c
zSSO_E	.RR:H5VR#H_I8_0ENNss$254Rj>R2CRoMNCs0RC
RRRRRzRRd:jRRsVFRH[RM#R5_8IH0NE_s$sN5R42-2R4RI8FMR0FjCRoMNCs0RC
RRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)Rzqnv4RD:RNDLCRRH#"a11"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloMC5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*nRM+RkOl_C_DDdd.*.&2RR""WRH&RMo0CCHs'lCNo58IH0UE-*I#_HE80_sNsNd$52*-.[2-.R"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05lMk_DOCD._4U.*4URR+M_klODCD_*ncn+cRRlMk_DOCD._d*Rd.+nR4,CR8b20E2RR&"RX"&MRH0CCosl'HN5oCI0H8E*-U#H_I8_0ENNss$25d-[.*2R;
RRRRRRRRRLRRCMoH
RRRRRRRRRRRRqz)vR4n:qR)vX4n.
1RRRRRRRRRRRRRRRRRb0FsRblNRj57RR=>#M_H_osC58IH0UE-*I#_HE80_sNsNd$52*-.[2-.,4R7RR=>#M_H_osC58IH0UE-*I#_HE80_sNsNd$52*-.[2-4,jRqRR=>D_FINs885,j2RRq4=D>RFNI_858s4R2,q=.R>FRDI8_N8.s52R,
RRRRRRRRRRRRRRRRRRRRRRRRRRqd=D>RFNI_858sdR2,W= R>sRI0M_C_,4nRpWBi>R=RiBp,jRmRR=>F_k0L_k#4Mn5kOl_C_DD4In,HE80-#U*_8IH0NE_s$sN5-d2.-*[.
2,SSSSSRSRm=4R>kRF0k_L#n_45lMk_DOCDn_4,8IH0UE-*I#_HE80_sNsNd$52*-.[2-42R;
RRRRRRRRRRRRR#RR_0Fk_osC58IH0UE-*I#_HE80_sNsNd$52*-.[2-4RR<=F_k0L_k#4Mn5kOl_C_DD4In,HE80-#U*_8IH0NE_s$sN5-d2.-*[4I2RERCM50Fk__CM4=nRR''42DRC#'CRZ
';RRRRRRRRRRRRRRRR#k_F0C_soH5I8-0EU_*#I0H8Es_Ns5N$d.2-*.[-2=R<R0Fk_#Lk_54nM_klODCD_,4nI0H8E*-U#H_I8_0ENNss$25d-[.*-R.2IMECRk5F0M_C_R4n=4R''C2RDR#C';Z'
RRRRRRRR8CMRMoCC0sNCdRzjS;
S8CMRMoCC0sNCORzE.	_;S
Sz	OE_:4RRRHV5I#_HE80_sNsNj$52RR>jo2RCsMCN
0CRRRRRRRRzRd4:VRHRH5I8R0ElRF8URR=4o2RCsMCN
0CRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FzVR)4qvnRR:DCNLD#RHR1"1a&"RR0HMCsoC'NHloIC5HE802RR&"R7"&MRH0CCosl'HN5oCM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*cRR+M_klODCD_*d.dR.2&WR""RR&HCM0o'CsHolNC25jR"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05lMk_DOCD._4U.*4URR+M_klODCD_*ncn+cRRlMk_DOCD._d*Rd.+nR4,CR8b20E2RR&"RX"&MRH0CCosl'HN5oC4
2;RRRRRRRRRRRRLHCoMR
RRRRRRRRRR)Rzqnv4R):Rqnv4XR41
RRRRRRRRRRRRRRRRsbF0NRlb7R5RR=>#M_H_osC5,j2RRqj=D>RFNI_858sjR2,q=4R>FRDI8_N84s52q,R.>R=RIDF_8N8s25.,R
RRRRRRRRRRRRRRRRRRRRRRRRRq=dR>FRDI8_N8ds52W,R >R=R0Is__CM4Rn,WiBpRR=>B,piR=mR>kRF0k_L#n_45lMk_DOCDn_4,2j2;R
RRRRRRRRRRRRRR_R#F_k0s5Coj<2R=kRF0k_L#n_45lMk_DOCDn_4,Rj2IMECRk5F0M_C_R4n=4R''C2RDR#C';Z'
RRRRRRRR8CMRMoCC0sNCdRz4S;
S8CMRMoCC0sNCORzE4	_;R
RRCRRMo8RCsMCNR0Cz;.6RRRRRRRRRRR
RMRC8CRoMNCs0zCRc
c;CRM8NEsOHO0C0CksR_MFsOI_E	CO;-

--
-
----NRp#H0RlCbDl0CMNF0HM#RHRV8CN0kD

--NEsOHO0C0CksRD#CC_O0sRNlF)VRq)v_W#RH
lOFbCFMMX0R)4qv.4UX1b
RFRs05R
RR:mRR0FkR8#0_oDFH
O;RqRRjRR:H#MR0D8_FOoH;R
RRRq4:MRHR8#0_oDFH
O;RqRR.RR:H#MR0D8_FOoH;R
RRRqd:MRHR8#0_oDFH
O;RqRRcRR:H#MR0D8_FOoH;R
RRRq6:MRHR8#0_oDFH
O;RqRRnRR:H#MR0D8_FOoH;R
RR:7RRRHM#_08DHFoOR;
RBRWp:iRRRHM#_08DHFoOR;
R RWRH:RM0R#8F_Do
HOR
2;CRM8ObFlFMMC0
;

lOFbCFMMX0R)nqvc1X.
FRbs50R
RRRm:jRR0FkR8#0_oDFH
O;RmRR4RR:FRk0#_08DHFoOR;
RjRqRH:RM0R#8F_Do;HO
RRRq:4RRRHM#_08DHFoOR;
R.RqRH:RM0R#8F_Do;HO
RRRq:dRRRHM#_08DHFoOR;
RcRqRH:RM0R#8F_Do;HO
RRRq:6RRRHM#_08DHFoOR;
RjR7RH:RM0R#8F_Do;HO
RRR7:4RRRHM#_08DHFoOR;
RBRWp:iRRRHM#_08DHFoOR;
R RWRH:RM0R#8F_Do
HOR
2;CRM8ObFlFMMC0
;
ObFlFMMC0)RXq.vdX
c1RsbF0
R5RmRRjRR:FRk0#_08DHFoOR;
R4RmRF:Rk#0R0D8_FOoH;R
RRRm.:kRF00R#8F_Do;HO
RRRm:dRR0FkR8#0_oDFH
O;RqRRjRR:H#MR0D8_FOoH;R
RRRq4:MRHR8#0_oDFH
O;RqRR.RR:H#MR0D8_FOoH;R
RRRqd:MRHR8#0_oDFH
O;RqRRcRR:H#MR0D8_FOoH;R
RRR7j:MRHR8#0_oDFH
O;R7RR4RR:H#MR0D8_FOoH;R
RRR7.:MRHR8#0_oDFH
O;R7RRdRR:H#MR0D8_FOoH;R
RRpWBiRR:H#MR0D8_FOoH;R
RRRW :MRHR8#0_oDFHRO
2C;
MO8RFFlbM0CM;F
OlMbFCRM0Xv)qdU.X1R

b0FsRR5
RRRm:kRF00R#8F_Do_HOP0COF(s5RI8FMR0Fj
2;RqRRjRR:H#MR0D8_FOoH;R
RRRq4:MRHR8#0_oDFH
O;RqRR.RR:H#MR0D8_FOoH;R
RRRqd:MRHR8#0_oDFH
O;RqRRcRR:H#MR0D8_FOoH;R
RR:7RRRHM#_08DHFoOC_POs0F58(RF0IMF2Rj;R
RRpWBiRR:H#MR0D8_FOoH;R
RRRW :MRHR8#0_oDFHRO
2C;
MO8RFFlbM0CM;O

FFlbM0CMRqX)vX4nUR1
b0FsRR5
RRRm:kRF00R#8F_Do_HOP0COF(s5RI8FMR0Fj
2;RqRRjRR:H#MR0D8_FOoH;R
RRRq4:MRHR8#0_oDFH
O;RqRR.RR:H#MR0D8_FOoH;R
RRRqd:MRHR8#0_oDFH
O;R7RRRH:RM0R#8F_Do_HOP0COF(s5RI8FMR0Fj
2;RWRRBRpi:MRHR8#0_oDFH
O;RWRR RR:H#MR0D8_FOoH
;R2
8CMRlOFbCFMM
0;
b0$CCRDVP0FC0s_RRH#NNss$jR5RR0FdF2RVMRH0CCos0;
$RbCD0CVFsPC_.0_RRH#NNss$jR5RR0F4F2RVMRH0CCosV;
k0MOHRFMb5N8HRR:#_08DHFoOC_POs0F;4RI,.RIRH:RMo0CCRs2skC0s#MR0D8_FOoH_OPC0RFsHP#
NNsHLRDCPRNs:0R#8F_Do_HOP0COFIs54R-48MFI0jFR2L;
CMoH
VRRF[sRRRHMP'NssoNMCFRDFRb
RHRRV[R5RR<=IR.20MECRR
SRsPN5R[2:H=R5DH'F[I+2S;
CCD#
RSRP5Ns[:2R=jR''S;
CRM8H
V;RMRC8FRDF
b;RCRs0MksRsPN;M
C8NRb8V;
k0MOHRFMo_C0I0H8E5_UI0H8EH:RMo0CCRs2skC0sHMRMo0CCHsR#N
PsLHNDPCRN:DRR0HMCsoCRR:=jL;
CMoH
PRRN:DR=HRI8/0EUR;
RRHV5H5I8R0ElRF8U>2RRRc20MEC
RRRRDPNRR:=PRND+;R4
CRRMH8RVR;
R0sCkRsMP;ND
8CMR0oC_8IH0UE_;k
VMHO0FoMRCI0_HE80_I.5HE80:MRH0CCoss2RCs0kMMRH0CCos#RH
sPNHDNLCNRPDRR:HCM0oRCs:j=R;C
Lo
HMRNRPD=R:R8IH0.E/;R
RskC0sPMRN
D;CRM8o_C0I0H8E;_.
MVkOF0HMCRo0H_I850EI0H8ERR:HCM0o2CsR0sCkRsMD0CVFsPC_.0_R
H#PHNsNCLDRDPNRD:RCFV0P_Cs0;_.
oLCHRM
RDPN5R42:o=RCI0_HE80_I.5HE802R;
RRHV58IH0lERF.8RRj=R2ER0CRM
RPRRNjD52=R:R
j;RDRC#RC
RPRRNjD52=R:R
4;RMRC8VRH;R
RskC0sPMRN
D;CRM8o_C0I0H8EV;
k0MOHRFMo_C0I0H8EH5I8R0E:MRH0CCoss2RCs0kMCRDVP0FC0s_R
H#PHNsNCLDRDPNRD:RCFV0P_Cs0=R:R,5jRRj,jj,R2L;
CMoH
PRRNdD52=R:R0oC_8IH0UE_58IH0;E2
ORRNR#C58IH0lERFU8R2#RH
IRRERCMcRR|d>R=RDPN5R.2:4=R;R
RIMECR=.R>NRPD254RR:=4R;
RCIEMRR4=P>RNjD52=R:R
4;RERICFMR0sEC#>R=RDMkDR;
R8CMR#ONCR;
R0sCkRsMP;ND
8CMR0oC_8IH0
E;O#FM00NMR8IH0NE_s$sNRD:RCFV0P_Cs0=R:R0oC_8IH0IE5HE802O;
F0M#NRM0I0H8Es_Ns_N$n:cRRVDC0CFPs__0.=R:R0oC_8IH0IE5HE802V;
k0MOHRFMo_C0M_kl45.U80CbEH:RMo0CCRs2skC0sHMRMo0CCHsR#N
PsLHNDPCRN:DRR0HMCsoCRR:=jL;
CMoH
PRRN:DR=CR8b/0E4;.U
HRRV5R580CbEFRl8.R4U>2RR.442ER0CRM
RPRRN:DR=NRPDRR+4R;
R8CMR;HV
sRRCs0kMNRPDC;
Mo8RCM0_k4l_.
U;VOkM0MHFR0oC_VDC0CFPsc_n5b8C0:ERR0HMCsoC2CRs0MksR0HMCsoCR
H#LHCoMR
RskC0s8M5CEb0R8lFRU4.2C;
Mo8RCD0_CFV0P_Csn
c;VOkM0MHFR0oC_lMk_5nc80CbERR:HCM0o2CsR0sCkRsMHCM0oRCsHP#
NNsHLRDCPRND:MRH0CCos=R:R
j;LHCoMR
RH5VR80CbE=R<R.44R8NMRb8C0>ERR2cURC0EMR
RRPRRN:DR=;R4
CRRMH8RVR;
R0sCkRsMP;ND
8CMR0oC_lMk_;nc
MVkOF0HMCRo0C_DVP0FC8s5CEb0RH:RMo0CCRs;lRNG:MRH0CCoss2RCs0kMMRH0CCos#RH
sPNHDNLCNRPDRR:HCM0oRCs:j=R;C
Lo
HMRVRHRC58bR0E-NRlG=R>RRj20MEC
RRRRDPNRR:=80CbERR-l;NG
CRRD
#CRRRRPRND:8=RCEb0;R
RCRM8H
V;RCRs0Mks5DPN2C;
Mo8RCD0_CFV0P;Cs
MVkOF0HMCRo0k_Ml._d5b8C0:ERR0HMCsoC2CRs0MksR0HMCsoCR
H#PHNsNCLDRDPNRH:RMo0CC:sR=;Rj
oLCHRM
RRHV5b8C0<ER=URcR8NMRb8C0>ERR24nRC0EMR
RRPRRN:DR=;R4
CRRMH8RVR;
R0sCkRsMP;ND
8CMR0oC_lMk_;d.
MVkOF0HMCRo0k_Mln_45b8C0:ERR0HMCsoC2CRs0MksR0HMCsoCR
H#PHNsNCLDRDPNRH:RMo0CC:sR=;Rj
oLCHRM
RRHV5b8C0<ER=nR4R8NMRb8C0>ERRRj20MEC
RRRRNRPD=R:R
4;RMRC8VRH;R
RskC0sPMRN
D;CRM8o_C0M_kl4
n;VOkM0MHFR0oC_8CM_b8C0#E5HRxC:MRH0CCosRR;80CbERR:HCM0o2CsR0sCkRsMHCM0oRCsHP#
NNsHLRDCl_HM#CHxRH:RMo0CC:sR=;Rj
oLCHRM
RMlH_x#HC=R:Rb8C0
E;RVRHRH5#x<CRRb8C0RE20MEC
RRRRMlH_x#HC=R:Rx#HCR;
R8CMR;HV
sRRCs0kMHRlMH_#x
C;CRM8o_C0C_M880CbE-;
-MOF#M0N0kRMlC_ODRD#:MRH0CCos=R:R55580CbERR-4/2RR2d.R5+R5C58bR0E-2R4R8lFR2d.R4/Rn;22R-RR-RRyF)VRq.vdXR41ODCD#CRMC88CRF
OMN#0MM0RkOl_C_DD4R.U:MRH0CCos=R:R0oC_lMk_U4.5b8C0;E2
MOF#M0N0CRDVP0FCns_cRR:HCM0oRCs:o=RCD0_CFV0P_Csn8c5CEb02O;
F0M#NRM0M_klODCD_Rnc:MRH0CCos=R:R0oC_lMk_5ncD0CVFsPC_2nc;F
OMN#0MD0RCFV0P_Csd:.RR0HMCsoCRR:=o_C0D0CVFsPC5VDC0CFPsc_n,cRn2O;
F0M#NRM0M_klODCD_Rd.:MRH0CCos=R:R0oC_lMk_5d.D0CVFsPC_2d.;F
OMN#0MD0RCFV0P_Cs4:nRR0HMCsoCRR:=o_C0D0CVFsPC5VDC0CFPs._d,.Rd2O;
F0M#NRM0M_klODCD_R4n:MRH0CCos=R:R0oC_lMk_54nD0CVFsPC_24n;0

$RbCF_k0L_k#0C$b_U4.RRH#NNss$MR5kOl_C_DD4R.U8MFI0jFR,HRI8-0E4FR8IFM0RRj2F#VR0D8_FOoH;$
0bFCRkL0_k0#_$_bCnHcR#sRNsRN$5lMk_DOCDc_nRI8FMR0FjI,RHE80-84RF0IMF2RjRRFV#_08DHFoO0;
$RbCF_k0L_k#0C$b_Rd.HN#Rs$sNRk5MlC_ODdD_.FR8IFM0RRj,I0H8ER-48MFI0jFR2VRFR8#0_oDFH
O;0C$bR0Fk_#Lk_b0$Cn_4RRH#NNss$MR5kOl_C_DD48nRF0IMF,RjR8IH04E-RI8FMR0FjF2RV0R#8F_Do;HO
o#HMRNDF_k0L_k#4R.U:kRF0k_L#$_0b4C_.RU;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RVFR8k50RHkMb0FR0RH0s-N#002C#
o#HMRNDF_k0L_k#n:cRR0Fk_#Lk_b0$Cc_n;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFV80FkRM5HbRk000FRs#H-0CN0##2
HNoMDkRF0k_L#._dRF:RkL0_k0#_$_bCdR.;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RVFR8k50RHkMb0FR0RH0s-N#002C#
o#HMRNDF_k0L_k#4:nRR0Fk_#Lk_b0$Cn_4;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFV80FkRM5HbRk000FRs#H-0CN0##2
HNoMDkRF0M_CR#:R0D8_FOoH_OPC05FsM_klODCD_U4.RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-C-RMDNLCV#RF0sRs#H-0CN0#H
#oDMNR0Fk__CMn:cRR8#0_oDFH
O;#MHoNFDRkC0_M._dR#:R0D8_FOoH;H
#oDMNR0Fk__CM4:nRR8#0_oDFH
O;#MHoNIDRsC0_MRR:#_08DHFoOC_POs0F5lMk_DOCD._4UFR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--I0sHCMRCNCLD#FRVsNRCOsERFFIRVqR)vCROD
D##MHoNIDRsC0_Mc_nR#:R0D8_FOoH;H
#oDMNR0Is__CMd:.RR8#0_oDFH
O;#MHoNIDRsC0_Mn_4R#:R0D8_FOoH;H
#oDMNR_HMsRCo:0R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-k-R#RC80sFRC#oH0RCs7RQh
o#HMRNDF_k0sRCo:0R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-#RkC08RFCRso0H#C7sRm
za#MHoNNDR8C_soRR:#_08DHFoOC_POs0F58N8s8IH04E-RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RCk#8FR0RosCHC#0s7Rq7#)
HNoMDFRDI8_N8:sRR8#0_oDFHPO_CFO0sR5n8MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--Ns88R0LH#MRHbRk00)FRqOvRC#DDRR5cL#H0RJsCkCHs8O2
F0M#NRM0D_#LI0H8ERR:HCM0oRCs:I=RHE80-5U*I0H8Es_Ns5N$d42-2*-cI0H8Es_Ns5N$..2-*8IH0NE_s$sN5-42I0H8Es_Ns5N$j
2;0C$bRb0l_sNsNR$UHN#Rs$sNRH5I8_0ENNss$25d-84RF0IMF2RjRRFV#_08DHFoOC_POs0F58(RF0IMF2Rj;H
#oDMNRb0l_dU_.0,RlUb__R4n:lR0bs_NsUN$;0
N0LsHkR0C\N3slV_FV0#C\RR:#H0sM
o;LHCoMR

R-RR-VRQR8N8s8IH0<ERRN(R#o#HMjR''FR0RkkM#RC8L#H0
RRRRRzjRH:RVNR58I8sHE80R4=R2CRoMNCs0RC
RRRRRDRRFNI_8R8s<"=RjjjjjRj"&8RN_osC5;j2
RRRR8CMRMoCC0sNCjRz;R
RR4RzRRR:H5VRNs88I0H8ERR=.o2RCsMCN
0CRRRRRRRRD_FINs88RR<="jjjjRj"&8RN_osC584RF0IMF2Rj;R
RRMRC8CRoMNCs0zCR4R;
RzRR.:RRRRHV58N8s8IH0=ERRRd2oCCMsCN0
RRRRRRRRIDF_8N8s=R<Rj"jjRj"&8RN_osC58.RF0IMF2Rj;R
RRMRC8CRoMNCs0zCR.R;
RzRRd:RRRRHV58N8s8IH0=ERRRc2oCCMsCN0
RRRRRRRRIDF_8N8s=R<Rj"jj&"RR_N8s5CodFR8IFM0R;j2
RRRR8CMRMoCC0sNCdRz;z
ScRS:H5VRNs88I0H8ERR=6o2RCsMCN
0CSFSDI8_N8<sR=jR"j&"RR_N8s5CocFR8IFM0R;j2
MSC8CRoMNCs0zCRcS;
z:6SRRHV58N8s8IH0=ERRRn2oCCMsCN0
DSSFNI_8R8s<'=Rj&'RR_N8s5Co6FR8IFM0R;j2
RRRR8CMRMoCC0sNC6Rz;R
RRnRzRRR:H5VRNs88I0H8ERR>no2RCsMCN
0CRRRRRRRRD_FINs88RR<=Ns8_Cno5RI8FMR0Fj
2;RRRRCRM8oCCMsCN0R;zn
R
RR-R-RRQV5M8H_osC2CRso0H#C7sRQkhR#oHMRiBp
RRRRRz(RH:RV8R5HsM_CRo2oCCMsCN0
RRRRRRRRFbsO#C#Rp5Bi7,RQRh2LHCoMR
RRRRRRRRRRVRHRp5BiRR='R4'NRM8B'piCMPC002RE
CMRRRRRRRRRRRRRRRRHsM_C<oR=QR7hR;
RRRRRRRRRCRRMH8RVR;
RRRRRCRRMb8RsCFO#
#;RRRRCRM8oCCMsCN0R;z(
RRRRRzURH:RVMR5F80RHsM_CRo2oCCMsCN0
RRRRRRRRRRRR_HMsRCo<7=RQ
h;RRRRCRM8oCCMsCN0R;zU
R
RR-R-RRQV5k8F0C_sos2RC#oH0RCs7amzRHk#MmoRB
piRRRRzRgR:VRHRF58ks0_CRo2oCCMsCN0
RRRRRRRRFbsO#C#RB5mpRi,F_k0s2CoRoLCHRM
RRRRRRRRRHRRVmR5BRpi=4R''MRN8BRmpCi'P0CM2ER0CRM
RRRRRRRRRRRRR7RRmRza<F=Rks0_C
o;RRRRRRRRRRRRCRM8H
V;RRRRRRRRCRM8bOsFC;##
RRRR8CMRMoCC0sNCgRz;R
RR4Rzj:RRRRHV50MFRk8F0C_soo2RCsMCN
0CRRRRRRRRRRRR7amzRR<=F_k0s;Co
RRRR8CMRMoCC0sNC4Rzj
;
RRRR-Q-RVNR58_8ss2CoRosCHC#0s7Rq7k)R#oHMRiBp
RRRR4z4RRR:H5VRNs88_osC2CRoMNCs0RC
RRRRRbRRsCFO#5#RB,piR7q7)L2RCMoH
RRRRRRRRRRRRRHV5iBpR'=R4N'RMB8RpCi'P0CM2ER0CRM
RRRRRRRRRRRRRNRR8C_so=R<R7q7)85N8HsI8-0E4FR8IFM0R;j2
RRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMRFbsO#C#;R
RRMRC8CRoMNCs0zCR4
4;RRRRzR4.:VRHRF5M08RN8ss_CRo2oCCMsCN0
RRRRRRRRRRRR_N8sRCo<q=R7;7)
RRRR8CMRMoCC0sNC4Rz.R;
RRRRR
RRRRRR-t-RCsMCNR0C0REC)RqvODCD#MRN8CR#D0CORoDFHRO
RzRR4:dRRsVFRHHRMMR5kOl_C_DD4R.U-2R4RI8FMR0FjCRoMNCs0RC
R-RR-VRQR85N8HsI8R0E>2R6RCMC8FR0RCOsNR0CI0sHCMRCNCLDR8NMR0FkbRk0CLMND#CRCODC0FRDo
HORRRRRRRRzR4c:VRHR85N8HsI8R0E>2R(RMoCC0sNCR
RRRRRRRRRRRRRRkRF0M_C5RH2<'=R4I'RERCM5_N8s5CoNs88I0H8ER-48MFI0(FR2RR=HC2RDR#C';j'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RWRCIEMNR58C_so85N8HsI8-0E4FR8IFM0RR(2=2RHR#CDCjR''R;
RRRRRCRRMo8RCsMCNR0Cz;4c
RRRRR--Q5VRNs88I0H8E=R<RR62MIFRsCH0RNCMLRDCFFsRkk0b0MRCNCLDRD#CCRO0DHFoOCRMC88C
RRRRRRRR6z4RH:RVNR58I8sHE80RR<=(o2RCsMCN
0CRRRRRRRRRRRRRRRRF_k0CHM52=R<R''4;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R R;
RRRRRCRRMo8RCsMCNR0Cz;46
RRRRR--tCCMsCN0RC0ERv)qRDOCDN#RM08Rs#H-0CN0#R
RRRRRR4RznRR:VRFs[MRHRH5I8R0E-2R4RI8FMR0FjCRoMNCs0RC
RRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)Rzq.v4URR:DCNLD#RHR1"1a&"RR0HMCsoC'NHloIC5HE802RR&"R7"&MRH0CCosl'HN5oCH.*4U&2RR""WRH&RMo0CCHs'lCNo5R[2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50E54H+2.*4U8,RCEb02&2RR""XRH&RMo0CCHs'lCNo54[+2R;
RRRRRRRRRLRRCMoH
RRRRRRRRRRRRqz)vU4.RX:R)4qv.4UX1RR
RRRRRRRRRRRRRbRRFRs0lRNb5=7R>MRH_osC5,[2RRqj=D>RFNI_858sjR2,q=4R>FRDI8_N84s52q,R.>R=RIDF_8N8s25.,R
RRRRRRRRRRRRRRRRRRRRRRRRRq=dR>FRDI8_N8ds52q,Rc>R=RIDF_8N8s25c,6RqRR=>D_FINs885,62RRqn=D>RFNI_858sn
2,SSSSSRSRW= R>sRI0M_C5,H2RpWBi>R=RiBp,RRm=F>RkL0_k4#_.HU5,2[2;R
RRRRRRRRRRRRRRkRF0C_so25[RR<=F_k0L_k#45.UH2,[RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRMRC8CRoMNCs0zCR4
n;RRRRR8CMRMoCC0sNC4RzdR;RRRRRRRRRRRR
RRRRRR
RR-R-RMtCC0sNCRRN4InRFRs88bCCRv)qRDOCDVRHRbNbssFbHCN0RRRRRRRRRRRRR
RRRRRRzR4(:VRHRk5MlC_ODnD_cRR=4o2RCsMCN
0CRRRR-Q-RVNR58I8sHE80R(>R2CRMC08RFsROCCN0RHIs0CCRMDNLCMRN8kRF00bkRNCMLRDC#CCDOD0RFOoH
RRRRRRRRUz4NRR:H5VRNs88I0H8ERR>(o2RCsMCN
0CRRRRRRRRRRRRRRRRF_k0CnM_c=R<R''4RCIEM5R5Ns8_CNo58I8sHE80-84RF0IMF2R(RM=RkOl_C_DD42.UR8NMR85N_osC5Rn2=jR''R22CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C_Rnc<W=R ERIC5MR5_N8s5CoNs88I0H8ER-48MFI0(FR2RR=M_klODCD_U4.2MRN8NR58C_so25nR'=Rj2'2R#CDCjR''R;
RRRRRCRRMo8RCsMCNR0CzN4U;R
RRRRRR4RzU:LRRRHV58N8s8IH0=ERRN(RMM8RkOl_C_DD4R.U=2RjRMoCC0sNCR
RRRRRRRRRRRRRRkRF0M_C_Rnc<'=R4I'RERCM585N_osC5Rn2=jR''R22CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C_Rnc<W=R ERIC5MR5_N8s5Con=2RR''j2C2RDR#C';j'
RRRRRRRR8CMRMoCC0sNC4RzU
L;RRRR-Q-RVNR58I8sHE80RR<=6M2RFsRIHR0CCLMNDFCRskRF00bkRNCMLRDC#CCDOD0RFOoHRCMC8
C8RRRRRRRRzR4g:VRHR85N8HsI8R0E<n=R2CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_Mc_nRR<=';4'
RRRRRRRRRRRRRRRR0Is__CMn<cR= RW;R
RRRRRRMRC8CRoMNCs0zCR4
g;RRRR-t-RCsMCNR0C0REC)RqvODCDR8NMRH0s-N#00SC
RRRRz	OE_:.RRRHV58IH0NE_s$sN_5nc4>2RRRj2oCCMsCN0
RRRRRRRRjz.RV:RF[sRRRHM58IH0NE_s$sN_5nc4-2RRR428MFI0jFRRMoCC0sNCR
RRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqz)vRnc:NRDLRCDH"#R1"1aRH&RMo0CCHs'lCNo58IH0RE2&7R""RR&HCM0o'CsHolNCk5MlC_OD4D_.4U*.RU2&WR""RR&HCM0o'CsHolNCH5I8R0E-*R.[RR-.&2RR"" RH&RMo0CCHs'lCNo50oC_8CM_b8C0ME5kOl_C_DD4*.U4R.U+cRn,CR8b20E2RR&"RX"&MRH0CCosl'HN5oCI0H8ERR-.2*[;R
RRRRRRRRRRCRLo
HMRRRRRRRRRRRRzv)qn:cRRqX)vXnc.
1RRRRRRRRRRRRRRRRRb0FsRblNR457RR=>HsM_CIo5HE80-[.*-,42RR7j=H>RMC_soH5I8-0E.-*[.R2,q=jR>FRDI8_N8js52q,R4>R=RIDF_8N8s254,.RqRR=>D_FINs885,.2
RRRRRRRRRRRRRRRRRRRRRRRRqRRd>R=RIDF_8N8s25d,cRqRR=>D_FINs885,c2RRq6=D>RFNI_858s6
2,SSSSSRSRW= R>sRI0M_C_,ncRpWBi>R=RiBp,4RmRR=>F_k0L_k#nMc5kOl_C_DDnIc,HE80-[.*-,42RRmj=F>RkL0_kn#_ck5MlC_ODnD_cH,I8-0E.-*[.;22
RRRRRRRRRRRRRRRR0Fk_osC58IH0.E-*4[-2=R<R0Fk_#Lk_5ncM_klODCD_,ncI0H8E*-.[2-4RCIEMFR5kC0_Mc_nR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soH5I8-0E.-*[.<2R=kRF0k_L#c_n5lMk_DOCDc_n,8IH0.E-*.[-2ERIC5MRF_k0CnM_cRR='24'R#CDCZR''R;
RRRRRRRRCRM8oCCMsCN0Rjz.;S
SR8CMRMoCC0sNCORzE.	_;S
SREzO	R_4:VRHRH5I8_0ENNss$c_n5Rj2>2RjRMoCC0sNCR
RRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqz)vRnc:NRDLRCDH"#R1"1aRH&RMo0CCHs'lCNo58IH0RE2&7R""RR&HCM0o'CsHolNCk5MlC_OD4D_.4U*.RU2&WR""RR&HCM0o'CsHolNCH5I8R0E-*R.I0H8Es_Ns_N$n4c52RR-4&2RR"" RH&RMo0CCHs'lCNo50oC_8CM_b8C0ME5kOl_C_DD4*.U4R.U+cRn,CR8b20E2RR&"RX"&MRH0CCosl'HN5oCI0H8ERR-.H*I8_0ENNss$c_n5242;R
RRRRRRRRRRCRLo
HMRRRRRRRRRRRRzv)qn:cRRv)qn4cX1RR
RRRRRRRRRRRRRbRRFRs0lRNb5=7R>MRH_osC58IH0.E-*8IH0NE_s$sN_5nc442-2q,Rj>R=RIDF_8N8s25j,4RqRR=>D_FINs885,42RRq.=D>RFNI_858s.
2,RRRRRRRRRRRRRRRRRRRRRRRRRdRqRR=>D_FINs885,d2RRqc=D>RFNI_858scR2,q=6R>FRDI8_N86s52S,
SSSSSWRR >R=R0Is__CMnRc,WiBpRR=>B,piR=mR>kRF0k_L#c_n5lMk_DOCDc_n,8IH0.E-*8IH0NE_s$sN_5nc442-2
2;RRRRRRRRRRRRRRRRF_k0s5CoI0H8E*-.I0H8Es_Ns_N$n4c522-4RR<=F_k0L_k#nMc5kOl_C_DDnIc,HE80-I.*HE80_sNsNn$_c254-R42IMECRk5F0M_C_Rnc=4R''C2RDR#C';Z'
RRRRRRRRMRC8CRoMNCs0zCRO_E	4R;
RRRRSMRC8CRoMNCs0zCR4R(;RRRRRRRRRR

R-RR-CRtMNCs0NCRRR4nI8FsRC8CbqR)vCRODHDRVbRNbbsFs0HNCRRRRRRRRRRRRRRR
RRRR4z.RH:RVMR5kOl_C_DDd=.RRR42oCCMsCN0
RRRRR--Q5VRNs88I0H8ERR>6M2RCRC80OFRs0CNCsRIHR0CCLMNDNCRMF8Rkk0b0MRCNCLDRD#CCRO0DHFoOR
RRRRRR.Rz.:NRRRHV58N8s8IH0>ERRN(RMM8RkOl_C_DDn=cRRR42oCCMsCN0
RRRRRRRRRRRRRRRR0Fk__CMd<.R=4R''ERIC5MR5_N8s5CoNs88I0H8ER-48MFI0(FR2RR=M_klODCD_U4.2MRN8NR58C_so25nR'=R4R'2NRM85_N8s5Co6=2RR''j2C2RDR#C';j'
RRRRRRRRRRRRRRRR0Is__CMd<.R= RWRCIEM5R5Ns8_CNo58I8sHE80-84RF0IMF2R(RM=RkOl_C_DD42.UR8NMR85N_osC5Rn2=4R''N2RM58RNs8_C6o52RR='2j'2DRC#'CRj
';RRRRRRRRCRM8oCCMsCN0R.z.NR;
RRRRRzRR.R.L:VRHR85N8HsI8R0E>RR(NRM8M_klODCD_Rnc/4=R2CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_M._dRR<='R4'IMECRN558C_so85N8HsI8-0E4FR8IFM0RR(2=kRMlC_OD4D_.RU2NRM85_N8s5Con=2RR''j2MRN8NR58C_so256R'=Rj2'2R#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_M._dRR<=WI RERCM585N_osC58N8s8IH04E-RI8FMR0F(=2RRlMk_DOCD._4UN2RM58RNs8_Cno52RR='2j'R8NMR85N_osC5R62=jR''R22CCD#R''j;R
RRRRRRMRC8CRoMNCs0zCR.;.L
RRRRRRRR.z.ORR:H5VRNs88I0H8ERR=(MRN8kRMlC_ODnD_cRR=4o2RCsMCN
0CRRRRRRRRRRRRRRRRF_k0CdM_.=R<R''4RCIEM5R5Ns8_Cno52RR='24'R8NMR85N_osC5R62=jR''R22CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C_Rd.<W=R ERIC5MR5_N8s5Con=2RR''42MRN8NR58C_so256R'=Rj2'2R#CDCjR''R;
RRRRRCRRMo8RCsMCNR0CzO..;R
RRRRRR.Rz.:8RRRHV58N8s8IH0=ERRNnRMM8RkOl_C_DDn/cR=2R4RMoCC0sNCR
RRRRRRRRRRRRRRkRF0M_C_Rd.<'=R4I'RERCM585N_osC58N8s8IH04E-RI8FMR0F6=2RRlMk_DOCDc_n2C2RDR#C';j'
RRRRRRRRRRRRRRRR0Is__CMd<.R= RWRCIEM5R5Ns8_CNo58I8sHE80-84RF0IMF2R6RM=RkOl_C_DDn2c2R#CDCjR''R;
RRRRRCRRMo8RCsMCNR0Cz8..;R
RR-R-RRQV58N8s8IH0<ER=2R6RRMFI0sHCMRCNCLDRRFsFbk0kC0RMDNLCCR#D0CORoDFHMORCCC88R
RRRRRR.RzdRR:H5VRNs88I0H8E=R<RR62oCCMsCN0
RRRRRRRRRRRRRRRR0Fk__CMd<.R=4R''R;
RRRRRRRRRRRRRIRRsC0_M._dRR<=W
 ;RRRRRRRRCRM8oCCMsCN0Rdz.;R
RR-R-RMtCC0sNCER0CqR)vCRODNDRM08Rs#H-0CN0
RSRRORzEU	_RH:RVIR5HE80_sNsNd$52RR>jo2RCsMCN
0CSOSzED	_C:6RRRHV58IH0>ER=*RUI0H8Es_Ns5N$dN2RMI8RHE80RR>=Uo2RCsMCN
0CRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FzVR)dqv.RR:DCNLD#RHR1"1a&"RR0HMCsoC'NHloIC5HE802RR&"R7"&MRH0CCosl'HN5oCM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*c&2RR""WRH&RMo0CCHs'lCNo58IH0-ERRLD#_8IH0RE2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50EM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*cRR+dR.,80CbER22&XR""RR&HCM0o'CsHolNCH5I8R0E-#RDLH_I8R0E+2RU;R
RRRRRRRRRRCRLo
HMSRSRR)Rzq.vdRX:R)dqv.1XU
SSSRRRRb0FsRblNRR57=b>RNH85MC_soH5I8-0E4FR8IFM0R8IH0DE-#IL_HE802U,R,#RDLH_I8-0E4R2,q=jR>FRDI8_N8js52S,
SSSSSqRR4>R=RIDF_8N8s254,.RqRR=>D_FINs885,.2RRqd=D>RFNI_858sdR2,q=cR>FRDI8_N8cs52W,R >R=R0Is__CMdR.,WiBpRR=>B,pi
SSSSRSSR=mR>lR0b__Udj.52
2;SSSSNH##o:MRRsVFRRH[HIMRHE80-84RF0IMFHRI8-0ED_#LI0H8ECRoMNCs0SC
SRSSR0Fk_#Lk_5d.M_klODCD_,d.HR[2<0=RlUb__5d.jH25[H-I8+0ED_#LI0H8E
2;RRRRRRRRRRRRRRRRRkRF0C_so[5H2=R<R0Fk_#Lk_5d.M_klODCD_,d.HR[2IMECRk5F0M_C_Rd.=4R''C2RDR#C';Z'
SSSS8CMRMoCC0sNC#RN#MHo;R
RRRRRRRRRR.RzURR:VRFs[MRHR8IH0NE_s$sN5-d24FR8IFM0Ro4RCsMCN
0CRRRRRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqz)vRd.:NRDLRCDH"#R1"1aRH&RMo0CCHs'lCNo58IH0RE2&7R""RR&HCM0o'CsHolNCk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*2ncR"&RW&"RR0HMCsoC'NHloIC5HE80RD-R#IL_HE80R[-R*RU2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50EM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*cRR+dR.,80CbER22&XR""RR&HCM0o'CsHolNCH5I8R0E-#RDLH_I8R0E-[R5-*42U
2;RRRRRRRRRRRRRCRLo
HMRRRRRRRRRRRRR)Rzq.vdRX:R)dqv.1XURR
RRRRRRRRRRRRRRFRbsl0RN5bR7>R=R_HMs5CoI0H8E#-DLH_I8-0EU+*[(FR8IFM0R8IH0DE-#IL_HE80-[U*2q,Rj>R=RIDF_8N8s25j,4RqRR=>D_FINs885,42RRq.=D>RFNI_858s.
2,RRRRRRRRRRRRRRRRRRRRRRRRRdRqRR=>D_FINs885,d2RRqc=D>RFNI_858scR2,W= R>sRI0M_C_,d.RpWBi>R=RiBp,RRm=0>RlUb__5d.[;22
SSSRRRRNH##o:MRRsVFRRH[H(MRRI8FMR0FjCRoMNCs0SC
SRSSR0Fk_#Lk_5d.M_klODCD_,d.I0H8E#-DLH_I8-0EU+*[HR[2<0=RlUb__5d.[H25[
2;RRRRRRRRRRRRRRRRRkRF0C_soH5I8-0ED_#LI0H8E*-U[[+H2=R<R0Fk_#Lk_5d.M_klODCD_,d.I0H8E#-DLH_I8-0EU+*[HR[2IMECRk5F0M_C_Rd.=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR8CMRMoCC0sNC#RN#MHo;R
RRRRRRRRRRMRC8CRoMNCs0zCR.
U;SMSC8CRoMNCs0zCRO_E	D;C6
zSSO_E	oR06:VRHRH5I8R0E>U=RR8NMR8IH0lERFU8RRR>=6o2RCsMCN
0CRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FzVR)dqv.RR:DCNLD#RHR1"1a&"RR0HMCsoC'NHloIC5HE802RR&"R7"&MRH0CCosl'HN5oCM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*c&2RR""WRH&RMo0CCHs'lCNo58IH0-ERRLD#_8IH0RE2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50EM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*cRR+dR.,80CbER22&XR""RR&HCM0o'CsHolNCH5I8R0E-#RDLH_I8R0E+2RU;R
RRRRRRRRRRCRLo
HMSRSRR)Rzq.vdRX:R)dqv.1XU
SSSRRRRb0FsRblNRR57=b>RNH85MC_soH5I8-0E4FR8IFM0R8IH0DE-#IL_HE802U,R,#RDLH_I8-0E4R2,q=jR>FRDI8_N8js52S,
SSSSSqRR4>R=RIDF_8N8s254,.RqRR=>D_FINs885,.2RRqd=D>RFNI_858sdR2,q=cR>FRDI8_N8cs52W,R >R=R0Is__CMdR.,WiBpRR=>B,pi
SSSSRSSR=mR>lR0b__UdI.5HE80_sNsNd$522-42S;
SNSS#o#HMRR:VRFsHH[RMHRI8-0E4FR8IFM0R8IH0DE-#IL_HE80RMoCC0sNCS
SSRSRF_k0L_k#dM.5kOl_C_DDdH.,[<2R=lR0b__UdI.5HE80_sNsNd$522-45-H[I0H8E#+DLH_I820E;R
RRRRRRRRRRRRRRRRRF_k0s5CoHR[2<F=RkL0_kd#_.k5MlC_ODdD_.[,H2ERIC5MRF_k0CdM_.RR='24'R#CDCZR''S;
SCSSMo8RCsMCNR0CNH##o
M;RRRRRRRRRRRRzR.U:FRVsRR[HIMRHE80_sNsNd$52R-.8MFI0jFRRMoCC0sNCR
RRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqz)vRd.:NRDLRCDH"#R1"1aRH&RMo0CCHs'lCNo58IH0RE2&7R""RR&HCM0o'CsHolNCk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*2ncR"&RW&"RR0HMCsoC'NHlo[C5*RU2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50EM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*cRR+dR.,80CbER22&XR""RR&HCM0o'CsHolNC[55+*42U
2;RRRRRRRRRRRRRCRLo
HMRRRRRRRRRRRRR)Rzq.vdRX:R)dqv.1XURR
RRRRRRRRRRRRRRFRbsl0RN5bR7>R=R_HMs5CoU+*[(FR8IFM0R[U*2q,Rj>R=RIDF_8N8s25j,4RqRR=>D_FINs885,42RRq.=D>RFNI_858s.
2,RRRRRRRRRRRRRRRRRRRRRRRRRdRqRR=>D_FINs885,d2RRqc=D>RFNI_858scR2,W= R>sRI0M_C_,d.RpWBi>R=RiBp,RRm=0>RlUb__5d.[;22
SSSS#N#HRoM:FRVs[RHRRHM(FR8IFM0RojRCsMCN
0CSSSSRkRF0k_L#._d5lMk_DOCD._d,[U*+2H[RR<=0_lbU._d55[2H;[2
RRRRRRRRRRRRRRRRFRRks0_CUo5*H[+[<2R=kRF0k_L#._d5lMk_DOCD._d,[U*+2H[RCIEMFR5kC0_M._dR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRMRC8CRoMNCs0NCR#o#HMR;
RRRRRRRRRCRRMo8RCsMCNR0Cz;.U
CSSMo8RCsMCNR0Cz	OE_6o0;S
Sz	OE_:MRRRHV58IH0<ERRRU2oCCMsCN0
RRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVzv)qd:.RRLDNCHDR#1R"1Ra"&MRH0CCosl'HN5oCI0H8E&2RR""7RH&RMo0CCHs'lCNo5lMk_DOCD._4U.*4URR+M_klODCD_*ncnRc2&WR""RR&HCM0o'CsHolNC25jR"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05lMk_DOCD._4U.*4URR+M_klODCD_*ncn+cRR,d.Rb8C02E2R"&RX&"RR0HMCsoC'NHloUC52R;
RRRRRRRRRLRRCMoH
RSSRzRR)dqv.RR:Xv)qdU.X1S
SSRRRRsbF0NRlb7R5RR=>b5N8HsM_CIo5HE80-84RF0IMFHRI8-0ED_#LI0H8ER2,UD,R#IL_HE80-,42RRqj=D>RFNI_858sj
2,SSSSSRSRq=4R>FRDI8_N84s52q,R.>R=RIDF_8N8s25.,dRqRR=>D_FINs885,d2RRqc=D>RFNI_858scR2,W= R>sRI0M_C_,d.RpWBi>R=RiBp,S
SSSSSRRRm=0>RlUb__5d.j;22
SSSS#N#HRoM:FRVs[RHRRHMI0H8ER-48MFI0jFRRMoCC0sNCS
SSRSRF_k0L_k#dM.5kOl_C_DDdH.,[<2R=lR0b__Udj.52[5H2R;
RRRRRRRRRRRRRRRRR0Fk_osC52H[RR<=F_k0L_k#dM.5kOl_C_DDdH.,[I2RERCM50Fk__CMd=.RR''42DRC#'CRZ
';SSSSCRM8oCCMsCN0R#N#H;oM
CSSMo8RCsMCNR0Cz	OE_
M;SMSC8CRoMNCs0zCRO_E	US;
SEzO	R_c:VRHRH5I8_0ENNss$25.Rj>R2CRoMNCs0RC
RRRRRzRR.cc_RH:RVIR5HE80RR>=co2RCsMCN
0CRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FzVR)dqv.RR:DCNLD#RHR1"1a&"RR0HMCsoC'NHloIC5HE802RR&"R7"&MRH0CCosl'HN5oCM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*c&2RR""WRH&RMo0CCHs'lCNo5Rj2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50EM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*cRR+dR.,80CbER22&XR""RR&HCM0o'CsHolNC25c;R
RRRRRRRRRRCRLo
HMRRRRRRRRRRRRzv)qd:.RRqX)vXd.c
1RRRRRRRRRRRRRRRRRb0FsRblNRd57RR=>HsM_Cdo527,R.>R=R_HMs5Co.R2,7=4R>MRH_osC5,42RR7j=H>RMC_so25j,S
SSRRRRRRRRRRRRqRRj>R=RIDF_8N8s25j,4RqRR=>D_FINs885,42RRq.=D>RFNI_858s.
2,RRRRRRRRRRRRRRRRRRRRRRRRRdRqRR=>D_FINs885,d2RRqc=D>RFNI_858scR2,W= R>sRI0M_C_,d.RpWBi>R=RiBp,SR
SSSSSmRRd>R=R0Fk_#Lk_5d.M_klODCD_,d.dR2,m=.R>kRF0k_L#._d5lMk_DOCD._d,,.2
SSSSRSSRRm4=F>RkL0_kd#_.k5MlC_ODdD_.2,4,jRmRR=>F_k0L_k#dM.5kOl_C_DDdj.,2
2;RRRRRRRRRRRRRRRRF_k0s5Cod<2R=kRF0k_L#._d5lMk_DOCD._d,Rd2IMECRk5F0M_C_Rd.=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5R.2<F=RkL0_kd#_.k5MlC_ODdD_.2,.RCIEMFR5kC0_M._dR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so254RR<=F_k0L_k#dM.5kOl_C_DDd4.,2ERIC5MRF_k0CdM_.RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cjo52=R<R0Fk_#Lk_5d.M_klODCD_,d.jI2RERCM50Fk__CMd=.RR''42DRC#'CRZ
';RRRRRRRRCRM8oCCMsCN0Rcz._
c;RRRRRRRRz_.cdRR:H5VRI0H8ERR=do2RCsMCN
0CRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FzVR)dqv.RR:DCNLD#RHR1"1a&"RR0HMCsoC'NHloIC5HE802RR&"R7"&MRH0CCosl'HN5oCM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*c&2RR""WRH&RMo0CCHs'lCNo5Rj2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50EM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*cRR+dR.,80CbER22&XR""RR&HCM0o'CsHolNC25c;R
RRRRRRRRRRCRLo
HMRRRRRRRRRRRRzv)qd:.RRqX)vXd.c
1RRRRRRRRRRRRRRRRRb0FsRblNRd57RR=>',j'RR7.=H>RMC_so25.,4R7RR=>HsM_C4o527,Rj>R=R_HMs5Coj
2,SRSSRRRRRRRRRRRRRRqj=D>RFNI_858sjR2,q=4R>FRDI8_N84s52q,R.>R=RIDF_8N8s25.,R
RRRRRRRRRRRRRRRRRRRRRRRRRq=dR>FRDI8_N8ds52q,Rc>R=RIDF_8N8s25c, RWRR=>I_s0CdM_.W,RBRpi=B>RpRi,
SSSSRSSRRmd=F>Rb,CMRRm.=F>RkL0_kd#_.k5MlC_ODdD_.2,.,S
SSSSSR4RmRR=>F_k0L_k#dM.5kOl_C_DDd4.,2m,Rj>R=R0Fk_#Lk_5d.M_klODCD_,d.j;22
RRRRRRRRRRRRRRRR0Fk_osC5R.2<F=RkL0_kd#_.k5MlC_ODdD_.2,.RCIEMFR5kC0_M._dR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so254RR<=F_k0L_k#dM.5kOl_C_DDd4.,2ERIC5MRF_k0CdM_.RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cjo52=R<R0Fk_#Lk_5d.M_klODCD_,d.jI2RERCM50Fk__CMd=.RR''42DRC#'CRZ
';RRRRRRRRCRM8oCCMsCN0Rcz._
d;SMSC8CRoMNCs0zCRO_E	cS;
SEzO	R_.:VRHRH5I8_0ENNss$254Rj>R2CRoMNCs0RC
RRRRRzRR.:cRRsVFRH[RMIR5HE80_sNsN4$52RR-482RF0IMFRRjoCCMsCN0
RRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVzv)qd:.RRLDNCHDR#1R"1Ra"&MRH0CCosl'HN5oCI0H8E&2RR""7RH&RMo0CCHs'lCNo5lMk_DOCD._4U.*4URR+M_klODCD_*ncnRc2&WR""RR&HCM0o'CsHolNCH5I8-0EUH*I8_0ENNss$25d-[.*-R.2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50EM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*cRR+dR.,80CbER22&XR""RR&HCM0o'CsHolNCH5I8-0EUH*I8_0ENNss$25d-[.*2R;
RRRRRRRRRLRRCMoH
RRRRRRRRRRRRqz)vRd.:qR)vXd..
1RRRRRRRRRRRRRRRRRb0FsRblNRj57RR=>HsM_CIo5HE80-IU*HE80_sNsNd$52*-.[2-.,4R7RR=>HsM_CIo5HE80-IU*HE80_sNsNd$52*-.[2-4,jRqRR=>D_FINs885,j2RRq4=D>RFNI_858s4R2,q=.R>FRDI8_N8.s52R,
RRRRRRRRRRRRRRRRRRRRRRRRRRqd=D>RFNI_858sdR2,q=cR>FRDI8_N8cs52W,R >R=R0Is__CMdR.,WiBpRR=>B,piRRmj=F>RkL0_kd#_.k5MlC_ODdD_.H,I8-0EUH*I8_0ENNss$25d-[.*-,.2
SSSSRSSRRm4=F>RkL0_kd#_.k5MlC_ODdD_.H,I8-0EUH*I8_0ENNss$25d-[.*-242;R
RRRRRRRRRRRRRRkRF0C_soH5I8-0EUH*I8_0ENNss$25d-[.*-R42<F=RkL0_kd#_.k5MlC_ODdD_.H,I8-0EUH*I8_0ENNss$25d-[.*-R42IMECRk5F0M_C_Rd.=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC58IH0UE-*8IH0NE_s$sN5-d2.-*[.<2R=kRF0k_L#._d5lMk_DOCD._d,8IH0UE-*8IH0NE_s$sN5-d2.-*[.I2RERCM50Fk__CMd=.RR''42DRC#'CRZ
';RRRRRRRRCRM8oCCMsCN0Rcz.;S
SCRM8oCCMsCN0REzO	;_.
zSSO_E	4RR:H5VRI0H8Es_Ns5N$j>2RRRj2oCCMsCN0
RRRRRRRRcz.RH:RVIR5HE80R8lFR=URRR42oCCMsCN0
RRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVzv)qd:.RRLDNCHDR#1R"1Ra"&MRH0CCosl'HN5oCI0H8E&2RR""7RH&RMo0CCHs'lCNo5lMk_DOCD._4U.*4URR+M_klODCD_*ncnRc2&WR""RR&HCM0o'CsHolNC25jR"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05lMk_DOCD._4U.*4URR+M_klODCD_*ncn+cRR,d.Rb8C02E2R"&RX&"RR0HMCsoC'NHlo4C52R;
RRRRRRRRRLRRCMoH
RRRRRRRRRRRRqz)vRd.:qR)vXd.4
1RRRRRRRRRRRRRRRRRb0FsRblNRR57=H>RMC_so25j,jRqRR=>D_FINs885,j2RRq4=D>RFNI_858s4R2,q=.R>FRDI8_N8.s52R,
RRRRRRRRRRRRRRRRRRRRRRRRRRqd=D>RFNI_858sdR2,q=cR>FRDI8_N8cs52W,R >R=R0Is__CMdR.,WiBpRR=>B,piR=mR>kRF0k_L#._d5lMk_DOCD._d,2j2;R
RRRRRRRRRRRRRRkRF0C_so25jRR<=F_k0L_k#dM.5kOl_C_DDdj.,2ERIC5MRF_k0CdM_.RR='24'R#CDCZR''R;
RRRRRCRRMo8RCsMCNR0Cz;.c
CSSMo8RCsMCNR0Cz	OE_
4;RRRRCRM8oCCMsCN0R4z.;RRRRRRRR
RR
RRRRR--tCCMsCN0R4NRnFRIs88RCRCb)RqvODCDRRHVNsbbFHbsNR0CRRRRRRRRRRRRRRR
RzRR.:6RRRHV5lMk_DOCDn_4R4=R2CRoMNCs0RC
R-RR-VRQR85N8HsI8R0E>2R6RCMC8FR0RCOsNR0CI0sHCMRCNCLDR8NMR0FkbRk0CLMND#CRCODC0FRDo
HORRRRRRRRzN.nRH:RVNR58I8sHE80R(>RR8NMRlMk_DOCDc_nR4=RR8NMRlMk_DOCD._dR4=R2CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_Mn_4RR<='R4'IMECRN558C_so85N8HsI8-0E4FR8IFM0RR(2=kRMlC_OD4D_.RU2NRM85_N8s5Con=2RR''42MRN8NR58C_so256R'=R4R'2NRM85_N8s5Coc=2RR''j2C2RDR#C';j'
RRRRRRRRRRRRRRRR0Is__CM4<nR= RWRCIEM5R5Ns8_CNo58I8sHE80-84RF0IMF2R(RM=RkOl_C_DD42.UR8NMR85N_osC5Rn2=4R''N2RM58RNs8_C6o52RR='24'R8NMR85N_osC5Rc2=jR''R22CCD#R''j;R
RRRRRRMRC8CRoMNCs0zCR.;nN
RRRRRRRRnz.LRR:H5VRNs88I0H8ERR>(MRN8kRMlC_ODnD_cRR=4MRN8kRMlC_ODdD_.RR=jo2RCsMCN
0CRRRRRRRRRRRRRRRRF_k0C4M_n=R<R''4RCIEM5R5Ns8_CNo58I8sHE80-84RF0IMF2R(RM=RkOl_C_DD42.UR8NMR85N_osC5Rn2=4R''N2RM58RNs8_C6o52RR='2j'R8NMR85N_osC5Rc2=jR''R22CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C_R4n<W=R ERIC5MR5_N8s5CoNs88I0H8ER-48MFI0(FR2RR=M_klODCD_U4.2MRN8NR58C_so25nR'=R4R'2NRM85_N8s5Co6=2RR''j2MRN8NR58C_so25cR'=Rj2'2R#CDCjR''R;
RRRRRCRRMo8RCsMCNR0CzL.n;R
RRRRRR.Rzn:ORRRHV58N8s8IH0>ERRN(RMM8RkOl_C_DDn=cRRNjRMM8RkOl_C_DDd=.RRR42oCCMsCN0
RRRRRRRRRRRRRRRR0Fk__CM4<nR=4R''ERIC5MR5_N8s5CoNs88I0H8ER-48MFI0(FR2RR=M_klODCD_U4.2MRN8NR58C_so25nR'=RjR'2NRM85_N8s5Co6=2RR''42MRN8NR58C_so25cR'=Rj2'2R#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_Mn_4RR<=WI RERCM585N_osC58N8s8IH04E-RI8FMR0F(=2RRlMk_DOCD._4UN2RM58RNs8_Cno52RR='2j'R8NMR85N_osC5R62=4R''N2RM58RNs8_Cco52RR='2j'2DRC#'CRj
';RRRRRRRRCRM8oCCMsCN0Rnz.OR;
RRRRRzRR.Rn8:VRHR85N8HsI8R0E>RR(NRM8M_klODCD_Rnc=RRjNRM8M_klODCD_Rd.=2RjRMoCC0sNCR
RRRRRRRRRRRRRRkRF0M_C_R4n<'=R4I'RERCM585N_osC58N8s8IH04E-RI8FMR0F(=2RRlMk_DOCD._4UN2RM58RNs8_Cno52RR='2j'R8NMR85N_osC5R62=jR''N2RM58RNs8_Cco52RR='2j'2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0C4M_n=R<RRW IMECRN558C_so85N8HsI8-0E4FR8IFM0RR(2=kRMlC_OD4D_.RU2NRM85_N8s5Con=2RR''j2MRN8NR58C_so256R'=RjR'2NRM85_N8s5Coc=2RR''j2C2RDR#C';j'
RRRRRRRR8CMRMoCC0sNC.Rzn
8;RRRRRRRRzC.nRH:RVNR58I8sHE80R(=RR8NMRlMk_DOCDc_nR4=RR8NMRlMk_DOCD._dR4=R2CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_Mn_4RR<='R4'IMECRN558C_so25nR'=R4R'2NRM85_N8s5Co6=2RR''42MRN8NR58C_so25cR'=Rj2'2R#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_Mn_4RR<=WI RERCM585N_osC5Rn2=4R''N2RM58RNs8_C6o52RR='24'R8NMRNR58C_so25cR'=Rj2'2R#CDCjR''R;
RRRRRCRRMo8RCsMCNR0CzC.n;R
RRRRRR.Rzn:VRRRHV58N8s8IH0=ERRN(RMM8RkOl_C_DDn=cRRN4RMM8RkOl_C_DDd=.RRRj2oCCMsCN0
RRRRRRRRRRRRRRRR0Fk__CM4<nR=4R''ERIC5MR5_N8s5Con=2RR''42MRN8NR58C_so256R'=RjR'2NRM85_N8s5Coc=2RR''j2C2RDR#C';j'
RRRRRRRRRRRRRRRR0Is__CM4<nR= RWRCIEM5R5Ns8_Cno52RR='24'R8NMR85N_osC5R62=jR''N2RM58RNs8_Cco52RR='2j'2DRC#'CRj
';RRRRRRRRCRM8oCCMsCN0Rnz.VR;
RRRRRzRR.Rno:VRHR85N8HsI8R0E=RRnNRM8M_klODCD_Rnc=RRjNRM8M_klODCD_Rd.=2R4RMoCC0sNCR
RRRRRRRRRRRRRRkRF0M_C_R4n<'=R4I'RERCM585N_osC5R62=4R''N2RM58RNs8_Cco52RR='2j'2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0C4M_n=R<RRW IMECRN558C_so256R'=R4R'2NRM85_N8s5Coc=2RR''j2C2RDR#C';j'
RRRRRRRR8CMRMoCC0sNC.Rzn
o;RRRRRRRRzE.nRH:RVNR58I8sHE80R6=RR8NMRlMk_DOCD._dRR/=4o2RCsMCN
0CRRRRRRRRRRRRRRRRF_k0C4M_n=R<R''4RCIEM5R5Ns8_CNo58I8sHE80-84RF0IMF2RcRM=RkOl_C_DDd2.2R#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_Mn_4RR<=WI RERCM585N_osC58N8s8IH04E-RI8FMR0Fc=2RRlMk_DOCD._d2C2RDR#C';j'
RRRRRRRR8CMRMoCC0sNC.Rzn
E;RRRR-Q-RVNR58I8sHE80RR<=6M2RFsRIHR0CCLMNDFCRskRF00bkRNCMLRDC#CCDOD0RFOoHRCMC8
C8RRRRRRRRzR.(:VRHR85N8HsI8R0E<c=R2CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_Mn_4RR<=';4'
RRRRRRRRRRRRRRRR0Is__CM4<nR= RW;R
RRRRRRMRC8CRoMNCs0zCR.
(;RRRR-t-RCsMCNR0C0REC)RqvODCDR8NMRH0s-N#00SC
RRRRz	OE_:URRRHV58IH0NE_s$sN5Rd2>2RjRMoCC0sNCS
Sz	OE_6DCRH:RVIR5HE80RR>=UH*I8_0ENNss$25dR8NMR8IH0>ER=2RURMoCC0sNCR
RRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqz)vR4n:NRDLRCDH"#R1"1aRH&RMo0CCHs'lCNo58IH0RE2&7R""RR&HCM0o'CsHolNCk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*Rnc+kRMlC_ODdD_..*d2RR&"RW"&MRH0CCosl'HN5oCI0H8ERR-D_#LI0H8E&2RR"" RH&RMo0CCHs'lCNo50oC_8CM_b8C0ME5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*nRM+RkOl_C_DDdd.*.RR+4Rn,80CbER22&XR""RR&HCM0o'CsHolNCH5I8R0E-#RDLH_I8R0E+2RU;R
RRRRRRRRRRCRLo
HMSRSRR)Rzqnv4RX:R)4qvn1XU
SSSRRRRb0FsRblNRR57=b>RNH85MC_soH5I8-0E4FR8IFM0R8IH0DE-#IL_HE802U,R,#RDLH_I8-0E4R2,q=jR>FRDI8_N8js52S,
SSSSSqRR4>R=RIDF_8N8s254,.RqRR=>D_FINs885,.2RRqd=D>RFNI_858sdR2,W= R>sRI0M_C_,4nRpWBi>R=RiBp,S
SSSSSRRRm=0>RlUb__54nj;22
SSSS#N#HRoM:FRVs[RHRRHMI0H8ER-48MFI0IFRHE80-LD#_8IH0oERCsMCN
0CSSSSRkRF0k_L#n_45lMk_DOCDn_4,2H[RR<=0_lbUn_455j2HI[-HE80+LD#_8IH0;E2
RRRRRRRRRRRRRRRRFRRks0_CHo5[<2R=kRF0k_L#n_45lMk_DOCDn_4,2H[RCIEMFR5kC0_Mn_4R'=R4R'2CCD#R''Z;S
SSMSC8CRoMNCs0NCR#o#HMR;
RRRRRRRRRzRR.:URRsVFRH[RMHRI8_0ENNss$25d-84RF0IMFRR4oCCMsCN0
RRRRRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)Rzqnv4RD:RNDLCRRH#"a11"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloMC5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*nRM+RkOl_C_DDdd.*.&2RR""WRH&RMo0CCHs'lCNo58IH0-ERRLD#_8IH0-ERRU[*2RR&"R "&MRH0CCosl'HN5oCo_C0C_M880CbEk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*Rnc+kRMlC_ODdD_..*dR4+Rn8,RCEb02&2RR""XRH&RMo0CCHs'lCNo58IH0-ERRLD#_8IH0-ERR-5[4U2*2R;
RRRRRRRRRRRRRoLCHRM
RRRRRRRRRRRRRqz)vR4n:)RXqnv4XRU1
RRRRRRRRRRRRRRRRsbF0NRlb7R5RR=>HsM_CIo5HE80-LD#_8IH0UE-*([+RI8FMR0FI0H8E#-DLH_I8-0EU2*[,jRqRR=>D_FINs885,j2RRq4=D>RFNI_858s4R2,q=.R>FRDI8_N8.s52R,
RRRRRRRRRRRRRRRRRRRRRRRRRRqd=D>RFNI_858sdR2,W= R>sRI0M_C_,4nRpWBi>R=RiBp,RRm=0>RlUb__54n[;22
SSSRRRRNH##o:MRRsVFRRH[H(MRRI8FMR0FjCRoMNCs0SC
SRSSR0Fk_#Lk_54nM_klODCD_,4nI0H8E#-DLH_I8-0EU+*[HR[2<0=RlUb__54n[H25[
2;RRRRRRRRRRRRRRRRRkRF0C_soH5I8-0ED_#LI0H8E*-U[[+H2=R<R0Fk_#Lk_54nM_klODCD_,4nI0H8E#-DLH_I8-0EU+*[HR[2IMECRk5F0M_C_R4n=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR8CMRMoCC0sNC#RN#MHo;R
RRRRRRRRRRMRC8CRoMNCs0zCR.
U;SMSC8CRoMNCs0zCRO_E	D;C6
zSSO_E	oR06:VRHRH5I8R0E>U=RR8NMR8IH0lERFU8RRR>=6o2RCsMCN
0CRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FzVR)4qvnRR:DCNLD#RHR1"1a&"RR0HMCsoC'NHloIC5HE802RR&"R7"&MRH0CCosl'HN5oCM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*cRR+M_klODCD_*d.dR.2&WR""RR&HCM0o'CsHolNCH5I8R0E-#RDLH_I820ER"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05lMk_DOCD._4U.*4URR+M_klODCD_*ncn+cRRlMk_DOCD._d*Rd.+nR4,CR8b20E2RR&"RX"&MRH0CCosl'HN5oCI0H8ERR-D_#LI0H8ERR+U
2;RRRRRRRRRRRRLHCoMS
SRRRRzv)q4:nRRqX)vX4nUS1
SRSRRFRbsl0RN5bR7>R=R8bN5_HMs5CoI0H8ER-48MFI0IFRHE80-LD#_8IH0,E2RRU,D_#LI0H8E2-4,jRqRR=>D_FINs885,j2
SSSSRSSRRq4=D>RFNI_858s4R2,q=.R>FRDI8_N8.s52q,Rd>R=RIDF_8N8s25d, RWRR=>I_s0C4M_nW,RBRpi=B>Rp
i,SSSSSRSRm>R=Rb0l_4U_nH5I8_0ENNss$25d-242;S
SS#SN#MHoRV:RFHsR[MRHR8IH04E-RI8FMR0FI0H8E#-DLH_I8R0EoCCMsCN0
SSSSFRRkL0_k4#_nk5MlC_OD4D_n[,H2=R<Rb0l_4U_nH5I8_0ENNss$25d-542HI[-HE80+LD#_8IH0;E2
RRRRRRRRRRRRRRRRFRRks0_CHo5[<2R=kRF0k_L#n_45lMk_DOCDn_4,2H[RCIEMFR5kC0_Mn_4R'=R4R'2CCD#R''Z;S
SSMSC8CRoMNCs0NCR#o#HMR;
RRRRRRRRRzRR.:URRsVFRH[RMHRI8_0ENNss$25d-8.RF0IMFRRjoCCMsCN0
RRRRRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)Rzqnv4RD:RNDLCRRH#"a11"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloMC5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*nRM+RkOl_C_DDdd.*.&2RR""WRH&RMo0CCHs'lCNo5U[*2RR&"R "&MRH0CCosl'HN5oCo_C0C_M880CbEk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*Rnc+kRMlC_ODdD_..*dR4+Rn8,RCEb02&2RR""XRH&RMo0CCHs'lCNo5+5[4U2*2R;
RRRRRRRRRRRRRoLCHRM
RRRRRRRRRRRRRqz)vR4n:)RXqnv4XRU1
RRRRRRRRRRRRRRRRsbF0NRlb7R5RR=>HsM_CUo5*([+RI8FMR0FU2*[,jRqRR=>D_FINs885,j2RRq4=D>RFNI_858s4R2,q=.R>FRDI8_N8.s52R,
RRRRRRRRRRRRRRRRRRRRRRRRRRqd=D>RFNI_858sdR2,W= R>sRI0M_C_,4nRpWBi>R=RiBp,RRm=0>RlUb__54n[;22
SSSS#N#HRoM:FRVs[RHRRHM(FR8IFM0RojRCsMCN
0CSSSSRkRF0k_L#n_45lMk_DOCDn_4,[U*+2H[RR<=0_lbUn_455[2H;[2
RRRRRRRRRRRRRRRRFRRks0_CUo5*H[+[<2R=kRF0k_L#n_45lMk_DOCDn_4,[U*+2H[RCIEMFR5kC0_Mn_4R'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRMRC8CRoMNCs0NCR#o#HMR;
RRRRRRRRRCRRMo8RCsMCNR0Cz;.U
CSSMo8RCsMCNR0Cz	OE_6o0;S
Sz	OE_:MRRRHV58IH0<ERRRU2oCCMsCN0
RRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVzv)q4:nRRLDNCHDR#1R"1Ra"&MRH0CCosl'HN5oCI0H8E&2RR""7RH&RMo0CCHs'lCNo5lMk_DOCD._4U.*4URR+M_klODCD_*ncn+cRRlMk_DOCD._d*2d.R"&RW&"RR0HMCsoC'NHlojC52RR&"R "&MRH0CCosl'HN5oCo_C0C_M880CbEk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*Rnc+kRMlC_ODdD_..*dR4+Rn8,RCEb02&2RR""XRH&RMo0CCHs'lCNo5;U2
RRRRRRRRRRRRoLCHSM
SRRRRqz)vR4n:)RXqnv4X
U1SRSSRbRRFRs0lRNb5=7R>NRb8M5H_osC58IH04E-RI8FMR0FI0H8E#-DLH_I820E,,RURLD#_8IH04E-2q,Rj>R=RIDF_8N8s25j,S
SSSSSR4RqRR=>D_FINs885,42RRq.=D>RFNI_858s.R2,q=dR>FRDI8_N8ds52W,R >R=R0Is__CM4Rn,WiBpRR=>B,pi
SSSSRSSR=mR>lR0b__U4jn52
2;SSSSNH##o:MRRsVFRRH[HIMRHE80-84RF0IMFRRjoCCMsCN0
SSSSFRRkL0_k4#_nk5MlC_OD4D_n[,H2=R<Rb0l_4U_n25j52H[;R
RRRRRRRRRRRRRRRRRF_k0s5CoHR[2<F=RkL0_k4#_nk5MlC_OD4D_n[,H2ERIC5MRF_k0C4M_nRR='24'R#CDCZR''S;
SCSSMo8RCsMCNR0CNH##o
M;SMSC8CRoMNCs0zCRO_E	MS;
S8CMRMoCC0sNCORzEU	_;S
Sz	OE_:cRRRHV58IH0NE_s$sN5R.2>2RjRMoCC0sNCR
RRRRRR.RzgR_c:VRHRH5I8R0E>c=R2CRoMNCs0RC
RRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)Rzqnv4RD:RNDLCRRH#"a11"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloMC5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*nRM+RkOl_C_DDdd.*.&2RR""WRH&RMo0CCHs'lCNo5Rj2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50EM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*cRR+M_klODCD_*d.d+.RR,4nRb8C02E2R"&RX&"RR0HMCsoC'NHlocC52R;
RRRRRRRRRLRRCMoH
RRRRRRRRRRRRqz)vR4n:qR)vX4nc
1RRRRRRRRRRRRRRRRRb0FsRblNRd57RR=>HsM_Cdo527,R.>R=R_HMs5Co.R2,7=4R>MRH_osC5,42RR7j=H>RMC_so25j,S
SSRRRRRRRRRRRRqRRj>R=RIDF_8N8s25j,4RqRR=>D_FINs885,42RRq.=D>RFNI_858s.
2,RRRRRRRRRRRRRRRRRRRRRRRRRdRqRR=>D_FINs885,d2RRW =I>RsC0_Mn_4,BRWp=iR>pRBi
,RSSSSSRSRm=dR>kRF0k_L#n_45lMk_DOCDn_4,,d2RRm.=F>RkL0_k4#_nk5MlC_OD4D_n2,.,S
SSSSSR4RmRR=>F_k0L_k#4Mn5kOl_C_DD44n,2m,Rj>R=R0Fk_#Lk_54nM_klODCD_,4nj;22
RRRRRRRRRRRRRRRR0Fk_osC5Rd2<F=RkL0_k4#_nk5MlC_OD4D_n2,dRCIEMFR5kC0_Mn_4R'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so25.RR<=F_k0L_k#4Mn5kOl_C_DD4.n,2ERIC5MRF_k0C4M_nRR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o52=R<R0Fk_#Lk_54nM_klODCD_,4n4I2RERCM50Fk__CM4=nRR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Coj<2R=kRF0k_L#n_45lMk_DOCDn_4,Rj2IMECRk5F0M_C_R4n=4R''C2RDR#C';Z'
RRRRRRRR8CMRMoCC0sNC.Rzg;_c
RRRRRRRRgz._:dRRRHV58IH0=ERRRd2oCCMsCN0
RRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVzv)q4:nRRLDNCHDR#1R"1Ra"&MRH0CCosl'HN5oCI0H8E&2RR""7RH&RMo0CCHs'lCNo5lMk_DOCD._4U.*4URR+M_klODCD_*ncn+cRRlMk_DOCD._d*2d.R"&RW&"RR0HMCsoC'NHlojC52RR&"R "&MRH0CCosl'HN5oCo_C0C_M880CbEk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*Rnc+kRMlC_ODdD_..*dR4+Rn8,RCEb02&2RR""XRH&RMo0CCHs'lCNo5;c2
RRRRRRRRRRRRoLCHRM
RRRRRRRRRzRR)4qvnRR:)4qvn1XcRR
RRRRRRRRRRRRRRFRbsl0RN5bR7=dR>jR''7,R.>R=R_HMs5Co.R2,7=4R>MRH_osC5,42RR7j=H>RMC_so25j,S
SSRRRRRRRRRRRRqRRj>R=RIDF_8N8s25j,4RqRR=>D_FINs885,42RRq.=D>RFNI_858s.
2,RRRRRRRRRRRRRRRRRRRRRRRRRdRqRR=>D_FINs885,d2RRW =I>RsC0_Mn_4,BRWp=iR>pRBi
,RSSSSSRSRm=dR>bRFCRM,m=.R>kRF0k_L#n_45lMk_DOCDn_4,,.2
SSSSRSSRRm4=F>RkL0_k4#_nk5MlC_OD4D_n2,4,jRmRR=>F_k0L_k#4Mn5kOl_C_DD4jn,2
2;RRRRRRRRRRRRRRRRF_k0s5Co.<2R=kRF0k_L#n_45lMk_DOCDn_4,R.2IMECRk5F0M_C_R4n=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5R42<F=RkL0_k4#_nk5MlC_OD4D_n2,4RCIEMFR5kC0_Mn_4R'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so25jRR<=F_k0L_k#4Mn5kOl_C_DD4jn,2ERIC5MRF_k0C4M_nRR='24'R#CDCZR''R;
RRRRRCRRMo8RCsMCNR0Cz_.gdS;
S8CMRMoCC0sNCORzEc	_;S
Sz	OE_:.RRRHV58IH0NE_s$sN5R42>2RjRMoCC0sNCR
RRRRRRdRzjRR:VRFs[MRHRH5I8_0ENNss$254R4-R2FR8IFM0RojRCsMCN
0CRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FzVR)4qvnRR:DCNLD#RHR1"1a&"RR0HMCsoC'NHloIC5HE802RR&"R7"&MRH0CCosl'HN5oCM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*cRR+M_klODCD_*d.dR.2&WR""RR&HCM0o'CsHolNCH5I8-0EUH*I8_0ENNss$25d-[.*-R.2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50EM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*cRR+M_klODCD_*d.d+.RR,4nRb8C02E2R"&RX&"RR0HMCsoC'NHloIC5HE80-IU*HE80_sNsNd$52*-.[
2;RRRRRRRRRRRRLHCoMR
RRRRRRRRRR)Rzqnv4R):Rqnv4XR.1
RRRRRRRRRRRRRRRRsbF0NRlb7R5j>R=R_HMs5CoI0H8E*-UI0H8Es_Ns5N$d.2-*.[-27,R4>R=R_HMs5CoI0H8E*-UI0H8Es_Ns5N$d.2-*4[-2q,Rj>R=RIDF_8N8s25j,4RqRR=>D_FINs885,42RRq.=D>RFNI_858s.
2,RRRRRRRRRRRRRRRRRRRRRRRRRdRqRR=>D_FINs885,d2RRW =I>RsC0_Mn_4,BRWp=iR>pRBim,Rj>R=R0Fk_#Lk_54nM_klODCD_,4nI0H8E*-UI0H8Es_Ns5N$d.2-*.[-2S,
SSSSSmRR4>R=R0Fk_#Lk_54nM_klODCD_,4nI0H8E*-UI0H8Es_Ns5N$d.2-*4[-2
2;RRRRRRRRRRRRRRRRF_k0s5CoI0H8E*-UI0H8Es_Ns5N$d.2-*4[-2=R<R0Fk_#Lk_54nM_klODCD_,4nI0H8E*-UI0H8Es_Ns5N$d.2-*4[-2ERIC5MRF_k0C4M_nRR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_CIo5HE80-IU*HE80_sNsNd$52*-.[2-.RR<=F_k0L_k#4Mn5kOl_C_DD4In,HE80-IU*HE80_sNsNd$52*-.[2-.RCIEMFR5kC0_Mn_4R'=R4R'2CCD#R''Z;R
RRRRRRMRC8CRoMNCs0zCRd
j;SMSC8CRoMNCs0zCRO_E	.S;
SEzO	R_4:VRHRH5I8_0ENNss$25jRj>R2CRoMNCs0RC
RRRRRzRRd:4RRRHV58IH0lERFU8RR4=R2CRoMNCs0RC
RRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)Rzqnv4RD:RNDLCRRH#"a11"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloMC5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*nRM+RkOl_C_DDdd.*.&2RR""WRH&RMo0CCHs'lCNo5Rj2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50EM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*cRR+M_klODCD_*d.d+.RR,4nRb8C02E2R"&RX&"RR0HMCsoC'NHlo4C52R;
RRRRRRRRRLRRCMoH
RRRRRRRRRRRRqz)vR4n:qR)vX4n4
1RRRRRRRRRRRRRRRRRb0FsRblNRR57=H>RMC_so25j,jRqRR=>D_FINs885,j2RRq4=D>RFNI_858s4R2,q=.R>FRDI8_N8.s52R,
RRRRRRRRRRRRRRRRRRRRRRRRRRqd=D>RFNI_858sdR2,W= R>sRI0M_C_,4nRpWBi>R=RiBp,RRm=F>RkL0_k4#_nk5MlC_OD4D_n2,j2R;
RRRRRRRRRRRRRFRRks0_Cjo52=R<R0Fk_#Lk_54nM_klODCD_,4njI2RERCM50Fk__CM4=nRR''42DRC#'CRZ
';RRRRRRRRCRM8oCCMsCN0R4zd;S
SCRM8oCCMsCN0REzO	;_4
RRRRMRC8CRoMNCs0zCR.R6;RRRRRRRRRC

MN8RsHOE00COkRsC#CCDOs0_N
l;
