// --------------------------------------------------------------------
// >>>>>>>>>>>>>>>>>>>>>>>>> COPYRIGHT NOTICE <<<<<<<<<<<<<<<<<<<<<<<<<
// --------------------------------------------------------------------
// Copyright (c) 2005 by Lattice Semiconductor Corporation
// --------------------------------------------------------------------
//
//
//                     Lattice Semiconductor Corporation
//                     5555 NE Moore Court
//                     Hillsboro, OR 97214
//                     U.S.A.
//
//                     TEL: 1-800-Lattice  (USA and Canada)
//                          1-408-826-6000 (other locations)
//
//                     web: http://www.latticesemi.com/
//                     email: techsupport@latticesemi.com
//
// --------------------------------------------------------------------
//
// Simulation Library File for MACHXO2
//
// $Header: 
//
`timescale 1ns / 1ps
module PDPW8KC (DI17, DI16, DI15, DI14, DI13, DI12, DI11, DI10, DI9,
         DI8, DI7, DI6, DI5, DI4, DI3, DI2, DI1, DI0,
         ADW8, ADW7, ADW6, ADW5, ADW4, ADW3, ADW2, ADW1, ADW0,
         BE1, BE0,
         CEW, CLKW, CSW2, CSW1, CSW0,
         ADR12, ADR11, ADR10, ADR9, ADR8, ADR7, ADR6, ADR5,
         ADR4,  ADR3,  ADR2, ADR1, ADR0,
         CER, OCER, CLKR, CSR2, CSR1, CSR0, RST,
         DO17, DO16, DO15, DO14, DO13, DO12, DO11, DO10, DO9,
         DO8, DO7, DO6, DO5, DO4, DO3, DO2, DO1, DO0);

   parameter  DATA_WIDTH_W = 18;
   parameter  DATA_WIDTH_R = 9;
   parameter  REGMODE = "NOREG";
   parameter  CSDECODE_W = "0b000";
   parameter  CSDECODE_R = "0b000";
   parameter  GSR = "ENABLED";
   parameter  RESETMODE = "SYNC";
   parameter  ASYNC_RESET_RELEASE = "SYNC";
   parameter  INIT_DATA = "STATIC";

parameter INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
parameter INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
parameter INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
parameter INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
parameter INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
parameter INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
parameter INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
parameter INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
parameter INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
parameter INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
parameter INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
parameter INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
parameter INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
parameter INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
parameter INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
parameter INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
parameter INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
parameter INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
parameter INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
parameter INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
parameter INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
parameter INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
parameter INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
parameter INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
parameter INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
parameter INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
parameter INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
parameter INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
parameter INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
parameter INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
parameter INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
parameter INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";

input    DI17, DI16, DI15, DI14, DI13, DI12, DI11, DI10, DI9,
         DI8, DI7, DI6, DI5, DI4, DI3, DI2, DI1, DI0,
         ADW8, ADW7, ADW6, ADW5, ADW4, ADW3, ADW2, ADW1, ADW0,
         BE1, BE0,
         CEW, CLKW, CSW2, CSW1, CSW0,
         ADR12, ADR11, ADR10, ADR9, ADR8, ADR7, ADR6, ADR5,
         ADR4,  ADR3,  ADR2, ADR1, ADR0,
         CER, OCER, CLKR, CSR2, CSR1, CSR0, RST;

output   DO17, DO16, DO15, DO14, DO13, DO12, DO11, DO10, DO9,
         DO8, DO7, DO6, DO5, DO4, DO3, DO2, DO1, DO0;

reg lo;
reg hi;

initial
begin
   lo = 1'b0;
   hi = 1'b1;
end

DP8KC EBR_INST (.DIA0(DI0), .DIA1(DI1), .DIA2(DI2), .DIA3(DI3), .DIA4(DI4),
       .DIA5(DI5), .DIA6(DI6), .DIA7(DI7), .DIA8(DI8), .DIB0(DI9), .DIB1(DI10), 
       .DIB2(DI11), .DIB3(DI12), .DIB4(DI13), .DIB5(DI14), .DIB6(DI15),
       .DIB7(DI16), .DIB8(DI17), 
       .CEA(CEW), .CLKA(CLKW), .WEA(hi), .CSA0(CSW0), .CSA1(CSW1),
       .CSA2(CSW2), .RSTA(RST), .ADA0(BE0), .ADA1(BE1), .ADA2(lo), .ADA3(lo), 
       .ADA4(ADW0), .ADA5(ADW1), .ADA6(ADW2), .ADA7(ADW3), .ADA8(ADW4), .ADA9(ADW5),
       .ADA10(ADW6), .ADA11(ADW7), .ADA12(ADW8), .CEB(CER), .CLKB(CLKR), .WEB(lo),
       .CSB0(CSR0), .CSB1(CSR1), .CSB2(CSR2), .RSTB(RST), .ADB0(ADR0), .ADB1(ADR1), 
       .ADB2(ADR2), .ADB3(ADR3), .ADB4(ADR4), .ADB5(ADR5), .ADB6(ADR6), .ADB7(ADR7), 
       .ADB8(ADR8), .ADB9(ADR9), .ADB10(ADR10), .ADB11(ADR11), .ADB12(ADR12), 
       .OCEA(lo), .OCEB(OCER),
       .DOB0(DO0), .DOB1(DO1), .DOB2(DO2), .DOB3(DO3), .DOB4(DO4), .DOB5(DO5), .DOB6(DO6), 
       .DOB7(DO7), .DOB8(DO8), .DOA0(DO9), .DOA1(DO10), .DOA2(DO11), .DOA3(DO12),
       .DOA4(DO13), .DOA5(DO14), .DOA6(DO15), .DOA7(DO16), .DOA8(DO17)); 

defparam EBR_INST.DATA_WIDTH_A = 18;
defparam EBR_INST.DATA_WIDTH_B = DATA_WIDTH_R;
defparam EBR_INST.REGMODE_A = REGMODE;
defparam EBR_INST.REGMODE_B = REGMODE;
defparam EBR_INST.CSDECODE_A = CSDECODE_W;
defparam EBR_INST.CSDECODE_B = CSDECODE_R;
defparam EBR_INST.GSR = GSR;
defparam EBR_INST.RESETMODE = RESETMODE;
defparam EBR_INST.ASYNC_RESET_RELEASE = ASYNC_RESET_RELEASE;
defparam EBR_INST.INITVAL_00 = INITVAL_00;
defparam EBR_INST.INITVAL_01 = INITVAL_01;
defparam EBR_INST.INITVAL_02 = INITVAL_02;
defparam EBR_INST.INITVAL_03 = INITVAL_03;
defparam EBR_INST.INITVAL_04 = INITVAL_04;
defparam EBR_INST.INITVAL_05 = INITVAL_05;
defparam EBR_INST.INITVAL_06 = INITVAL_06;
defparam EBR_INST.INITVAL_07 = INITVAL_07;
defparam EBR_INST.INITVAL_08 = INITVAL_08;
defparam EBR_INST.INITVAL_09 = INITVAL_09;
defparam EBR_INST.INITVAL_0A = INITVAL_0A;
defparam EBR_INST.INITVAL_0B = INITVAL_0B;
defparam EBR_INST.INITVAL_0C = INITVAL_0C;
defparam EBR_INST.INITVAL_0D = INITVAL_0D;
defparam EBR_INST.INITVAL_0E = INITVAL_0E;
defparam EBR_INST.INITVAL_0F = INITVAL_0F;
defparam EBR_INST.INITVAL_10 = INITVAL_10;
defparam EBR_INST.INITVAL_11 = INITVAL_11;
defparam EBR_INST.INITVAL_12 = INITVAL_12;
defparam EBR_INST.INITVAL_13 = INITVAL_13;
defparam EBR_INST.INITVAL_14 = INITVAL_14;
defparam EBR_INST.INITVAL_15 = INITVAL_15;
defparam EBR_INST.INITVAL_16 = INITVAL_16;
defparam EBR_INST.INITVAL_17 = INITVAL_17;
defparam EBR_INST.INITVAL_18 = INITVAL_18;
defparam EBR_INST.INITVAL_19 = INITVAL_19;
defparam EBR_INST.INITVAL_1A = INITVAL_1A;
defparam EBR_INST.INITVAL_1B = INITVAL_1B;
defparam EBR_INST.INITVAL_1C = INITVAL_1C;
defparam EBR_INST.INITVAL_1D = INITVAL_1D;
defparam EBR_INST.INITVAL_1E = INITVAL_1E;
defparam EBR_INST.INITVAL_1F = INITVAL_1F;

endmodule
