-- $Header: //synplicity/maplat2018q2p1/mappers/xilinx/lib/generic/gen_generic/seq_srl.vhd#1 $
@EH
DLssN$ RQ 
 ;kR#CQ   38#0_oDFH4O_43ncN;DD
Ck#R Q  03#8F_Do_HOkHM#o8MC3DND;#
kC RQ # 30D8_FOoH_HNs0NE3D
D;DsHLNRs$k#MHH
l;kR#Ck#MHHPl3ObFlFMMC0N#3D
D;
0CMHR0$1_ T1R)pHR#
RMoCCOsH5R
RRRRRNs88_8IH0:ERR0HMCsoCRR:=(R;
RRRRR8N8sH_#x:CRR0HMCsoCRR:=n
6;RRRRR_R8I0H8ERR:HCM0oRCs:U=R;R
RRRRRHH#_M0bkRL:RFCFDN:MR=sR0k
C;RRRRR#RH_0FkbRk0:FRLFNDCM=R:Rk0sC
2;RFRbs
05RRRRRqR)7R7):MRHR8#0_oDFHPO_CFO0s85N8Is_HE80-84RF0IMF2Rj;R
RRRRR7qqaRRRR:MRHR8#0_oDFHPO_CFO0s_58I0H8ER-48MFI0jFR2R;
RRRRRRW RRR:H#MR0D8_FOoH;R
RRRRRBRpiRH:RM0R#8F_Do;HO
RRRRqRR_a)1RRR:H#MR0D8_FOoH;R
RRRRR11_)a:RRRRHM#_08DHFoOR;
RRRRRz7maRRRRF:Rk#0R0D8_FOoH_OPC05Fs8H_I8-0E4FR8IFM0R2j2;M
C8 R1T)_1p
;
NEsOHO0C0CksRosCHC#0sF#RV R1T)_1p#RH
b0$CsR#Ds_NsRN$HN#Rs$sNRR5j08FR_8IH04E-2VRFR8#0_oDFHPO_CFO0s85N8#s_H-xC4FR8IFM0R;j2
o#HMRNDJM_H0RR:#_sDNNss$L;
CMoH
zRR4RR:VRFsHMRHR0jRF_R8I0H8E4R-RMoCC0sNCR
RRsRbF#OC#p5BiR2
RLRRCMoH
RSRH5VRsHH#MCo_85oCB2pi2ER0CSM
RHRRVWR5 RR='24'RC0EMS
SH5VRNs88_x#HCRR>402RE
CMSJSS_0HM5RH2<5=RJM_H025H58N8sH_#x.C-RI8FMR0Fj&2RRa7qq25H2S;
S#CDCS
SSHJ_MH05225jRR<=7qqa5;H2
CSSMH8RVS;
RCRRMH8RVS;
RMRC8VRH;C
SMb8RsCFO#
#;Sz7ma25HRR<=JM_H025H5MOFPM_H0CCosq5)727)2R;
R8CMRMoCC0sNC4Rz;C

Ms8RC#oH0#Cs;



ONsECH0Os0kC0R#NO0H_D#sRRFV1_ T1R)pHV#
k0MOHRFMM_klODCD5:MRR0HMCsoC;#RH_bHMkR0,HF#_kk0b0RR:LDFFC2NMskC0sHMRMo0CCHsR#RRRRPR
NNsHLRDCPkNDCRR:HCM0o;Cs
sPNHDNLCkRMlC_so:#RR0HMCsoC;C
Lo
HMRkRMlC_so:#R=;Rj
HRRV#5H_bHMkR020MECRR
RRRRRM_kls#CoRR:=M_kls#CoR4+R;R
RCRM8H
V;RVRH5_H#Fbk0kR020MECRR
RRRRRRlMk_osC#=R:RlMk_osC#RR+4R;
R8CMR;HV
PRRNCDkRR:=5-MRRlMk_osC#42/nR;
R0sCkRsMPkNDCC;
MM8RkOl_C;DD
k
VMHO0FsMRCHlNMoHM_osC5RM:HCM0o;CsR_H#HkMb0H,R#k_F00bkRL:RFCFDNsM2Cs0kMMRH0CCos#RHRRRRRN
PsLHNDPCRNCDkRH:RMo0CC
s;PHNsNCLDRlMk_osC#RR:HCM0o;Cs
oLCHRM
RlMk_osC#=R:R
j;RNRPDRkC:j=R;R
RHHV5#M_Hb2k0RC0EMRR
RRRRRlMk_osC#=R:RlMk_osC#RR+4R;
R8CMR;HV
HRRV#5H_0Fkb2k0RC0EMRR
RRRRRkRMlC_so:#R=kRMlC_so+#RR
4;RMRC8VRH;R
RPkNDC=R:RR5M-kRMlC_soR#2sRCl4
n;RCRs0MksRDPNk
C;CRM8sNClHMMHoC_so
;
VOkM0MHFRN#0sM0HoC_so#5H_bHMk:0RRFLFDMCN2CRs0MksR0HMCsoCR
H#LHCoMR
RHHV5#M_Hb2k0RC0EMR
RRRRRskC0s4MR;R
RCRM8H
V;RCRs0MksR
j;CRM8#s0N0oHM_osC;V

k0MOHRFMbVsCHoG_CHM5#k_F00bkRL:RFCFDNRM2skC0s#MR0MsHo#RH
oLCHRM
R5HVHF#_kk0b002RE
CMRRRRRCRs0MksRa"pa
";RMRC8VRH;R
RskC0s"MRp"wa;M
C8sRbCGVH_MoC;O

F0M#NRM0M_kl#_sDODCD#RR:HCM0oRCs:M=RkOl_C5DDNs88_x#HCH,R#M_Hb,k0R_H#Fbk0k;02
MOF#M0N0kRMl	_#Hsb_CRo#:MRH0CCos=R:RlsCNHHMMso_CNo58_8s#CHx,#RH_bHMkR0,HF#_kk0b0
2;O#FM00NMRlMk_N#0ss0_C:oRR0HMCsoCRR:=#s0N0oHM_osC5_H#HkMb0
2;O#FM00NMRD#s_CbsVRHG:0R#soHMRR:=bVsCHoG_CHM5#k_F00bk2
;
#MHoNDDR#:LRR8#0_oDFHPO_CFO0sR5d8MFI0jFR2=R:Rj"jj;j"
b0$C#RRs0D_lNb_s$sNRRH#NNss$jR5RR0F5lMk_D#s_DOCD+#RR242RRFV#_08DHFoOC_POs0F5I8_HE80R4-RRI8FMR0Fj
2;
o#HMRND0_lbNNss$RR:#_sD0_lbNNss$#;
HNoMDlR0b__8NNss$RR:#_sD0_lbNNss$#;
HNoMDlR0b8_N8:sRR8#0_oDFHPO_CFO0s85N8Is_HE80-84RF0IMF2Rj;H
#oDMNRb0l_0Fk_8N8sRR:#_08DHFoOC_POs0F5I8_HE80-84RF0IMF2Rj;N

0H0sLCk0R#\3sFD_VCV#0:\RRs#0H;Mo
C
Lo
HM
Rzj:VRHR_H#HkMb0CRoMNCs0
CRRsRbF#OC#p5BiR2
RoLCHRM
RHRRVsR5HM#Ho8_CoBC5p2i2RC0EMR
RRRRRH5VRW= RR''42ER0CRM
RRRRR0RRlNb_s$sN5Rj2<7=Rq;aq
RRRRCRRMH8RVR;
RCRRMH8RVR;
R8CMRFbsO#C#;CR
Mo8RCsMCN;0C
j
z4RR:HMVRFH05#M_Hb2k0RMoCC0sNCRR
RRRRR0RRlNb_s$sN5Rj2<7=Rq;aq
8CMRMoCC0sNC
;

4
z:VRHR8N8sH_I8R0E<c=RRMoCC0sNCR
RRCRLo
HMS#SDL=R<RhBmea_17m_pt_QBea BmM)5k#l_	_Hbs#CoR4-R,2Rc;R
RRRRRR4Rz4RR:VRFsHMRHR0jRF8R5_8IH0-ER4o2RCsMCN
0CSNSS0H0sLCk0R#\3sFD_VCV#0F\RV4Rz4:4RRLDNCHDR#sR#Ds_bCGVHRH&RMo0CCHs'lCNo5I8_HE802RR&"R7"&MRH0CCosl'HN5oCM_kl#s0N0C_so&2RR""WRH&RMo0CCHs'lCNo5RH2& R""RR&HCM0o'CsHolNCk5Ml0_#N_s0sRCo+kRMl	_#Hsb_C2o#R"&RX&"RR0HMCsoC'NHloHC5R4+R2S;
SCSLo
HMRRRRRRRRRRRRz444:)R1p 4n
RRRRRRRRRRRRsbF0NRlbR5
RRRRRRRRRRRRRqRRj>R=RLD#5,j2
RRRRRRRRRRRRRRRRRq4=D>R#4L52R,
RRRRRRRRRRRRRqRR.>R=RLD#5,.2
RRRRRRRRRRRRRRRRRqd=D>R#dL52R,
RRRRRRRRRRRRRBRR >R=R,W 
RRRRRRRRRRRRRRRRiBpRR=>B,pi
RRRRRRRRRRRRRRRR=7R>lR0bs_Ns5N$jH252R,
RRRRRRRRRRRRRTRRRR=>0_lb8s_Ns5N$jH252R
RRRRRRRRRR;R2
RRRRRRRR8CMRMoCC0sNC4Rz4R;
RRRRRzRR4:.RRRHVHF#_kk0b0CRoMNCs0
CRRRRRRRRRbOsFC5##O2D	
RRRRRRRRRRRRoLCHRM
RRRRRRRRRRRRRHRRVsR5HM#Ho8_CoBC5p2i2RC0EMR
RRRRRRRRRRRRRRRRRRVRHR 5WR'=R4R'20MEC
RRRRRRRRRRRRRRRRRRRRRRRRz7ma=R<Rb0l_N8_s$sN5;j2
RRRRRRRRRRRRRRRRRRRR8CMR;HV
RRRRRRRRRRRRRRRR8CMR;HV
RRRRRRRRRRRR8CMRFbsO#C#;RR
RRRRRCRRMo8RCsMCN;0C
RRRRRRRRdz4RH:RVFRM0#5H_0Fkb2k0RMoCC0sNCS
SRRRR7amzRR<=0_lb8s_Ns5N$j
2;RRRRRRRRCRM8oCCMsCN0Rdz4;M
C8CRoMNCs0zCR4
;
zR.:HNVR8_8sI0H8ERR>cCRoMNCs0RC
RLRRCMoH
RRRRRRRRR
RRRRRR.Rz.RR:VRFsHMRHR04RFMR5k#l_sOD_C#DD2CRoMNCs0
CRRRRRRRRRRRRRz4..:FRVsRR[HjMRRR0F5I8_HE80R2-4RMoCC0sNCS
SS0N0skHL0\CR3D#s_VFV#\C0RRFVz...RD:RNDLCRRH#"apw"RR&HCM0o'CsHolNC_58I0H8E&2RR""7RH&RMo0CCHs'lCNo5lMk_N#0ss0_C+oRRR5H-2R4*24nR"&RW&"RR0HMCsoC'NHlo[C52RR&"R "&MRH0CCosl'HN5oCM_kl#s0N0C_soRR+Hn*42RR&"RX"&MRH0CCosl'HN5oC[RR+4
2;RRRRRRRRRRRRLHCoMR
RRRRRRRRRRRRRR.Rz.R.:1B)p4
n RRRRRRRRRRRRRRRRb0FsRblN5R
RRRRRRRRRRRRRRjRqR'=>4
',RRRRRRRRRRRRRRRRq=4R>4R''R,
RRRRRRRRRRRRRqRR.>R=R''4,R
RRRRRRRRRRRRRRdRqRR=>',4'
RRRRRRRRRRRRRRRRRB =W>R R,
RRRRRRRRRRRRRBRRp=iR>pRBiR,
RRRRRRRRRRRRR7RRRR=>0_lbNNss$R5H-2R45,[2
RRRRRRRRRRRRRRRR6T4RR=>0_lbNNss$25H5,[2
SSSS=TR>lR0b__8NNss$R5H-2R45
[2RRRRRRRRRRRR2S;
SRS
RRRRRRRRRRRRRRRRR
RRRRRRRRRRRRRRCRM8oCCMsCN0R.Rz.
4;SzSS6H:RVk5Ml	_#Hsb_CRo#=2RjRMoCC0sNCSR
S0SSlFb_kN0_8R8s<0=Rl8b__sNsNM$5k#l_sOD_C#DDR4-R2S;
SMSC8CRoMNCs0zCR6R;
RRRRRCRRMo8RCsMCNR0Cz;..
RRRRRRRRR
RRRRRR.Rz.:dRR5HVM_kl#b	H_osC#=R/RRj2oCCMsCN0RS
SSLD#RR<=Bemh_71a_tpmQeB_ mBa)k5Ml	_#Hsb_CRo#-,R4R;c2
RRRRRRRRRRRR.z.cV:RF[sRRRHMjFR0R_58I0H8E4R-2CRoMNCs0SC
S0SN0LsHkR0C\s3#DV_FV0#C\VRFR.z..RR:DCNLD#RHRD#s_CbsVRHG&MRH0CCosl'HN5oC8H_I820ER"&R7&"RR0HMCsoC'NHloMC5k#l_00Ns_osCRM+Rk#l_sOD_C#DD*24nR"&RW&"RR0HMCsoC'NHlo[C52RR&"R "&MRH0CCosl'HN5oCM_kl#s0N0C_soRR+M_kl#_sDODCD#n*4RM+Rk#l_	_Hbs#Co2RR&"RX"&MRH0CCosl'HN5oC[RR+4
2;RRRRRRRRRRRRLHCoMR
RRRRRRRRRRRRRR.Rz.R.:1B)p4
n RRRRRRRRRRRRRRRRb0FsRblN5R
RRRRRRRRRRRRRRjRqRR=>D5#Lj
2,RRRRRRRRRRRRRRRRq=4R>#RDL254,R
RRRRRRRRRRRRRR.RqRR=>D5#L.
2,RRRRRRRRRRRRRRRRq=dR>#RDL25d,R
RRRRRRRRRRRRRR RBRR=>W
 ,RRRRRRRRRRRRRRRRBRpi=B>Rp
i,RRRRRRRRRRRRRRRR7>R=Rb0l_sNsNM$5k#l_sOD_C#DD225[,R
RRRRRRRRRRRRRR4RT6>R=Rb0l_sNsNM$5k#l_sOD_C#DDR4+R225[,S
SSRST=0>Rl8b__sNsNM$5k#l_sOD_C#DD225[
RRRRRRRRRRRR
2;S
SSRRRRRRRRRRRRCRM8oCCMsCN0R.Rz.
c;S0SSlFb_kN0_8R8s<0=Rl8b__sNsNM$5k#l_sOD_C#DD2R;
RRRRRCRRMo8RCsMCNR0Czd..;R
RRRRRR.RzdRR:HHVR#k_F00bkRMoCC0sNCRR
RRRRRbRRsCFO#O#5D
	2RRRRRRRRRRRRLHCoMR
RRRRRRRRRRRRRRVRHRH5s#oHM_oC8Cp5BiR220MEC
RRRRRRRRRRRRRRRRRRRRRHV5RW =4R''02RE
CMRRRRRRRRRRRRRRRRRRRRRRRR7amzRR<=0_lbF_k0Ns88;R
RRRRRRRRRRRRRRRRRRMRC8VRH;R
RRRRRRRRRRRRRRMRC8VRH;R
RRRRRRRRRRMRC8sRbF#OC#
;RRRRRRRRRCRM8oCCMsCN0;R
RRRRRR.RzcRR:HMVRFH05#k_F00bk2CRoMNCs0SC
SRRRRz7ma=R<Rb0l_0Fk_8N8sR;
RRRRRCRRMo8RCsMCNR0Cz;.c
8CMRMoCC0sNC.Rz;C

MN8RsHOE00COkRsC#00NH#O_s
D;
s
NO0EHCkO0s#CRCODC0s_#DVRFRT1 _p1)R
H#VOkM0MHFRlMk_DOCDR5M:MRH0CCosH;R#M_Hb,k0R_H#Fbk0k:0RRFLFDMCN20sCkRsMHCM0oRCsHR#RR
RRPHNsNCLDRDPNk:CRR0HMCsoC;N
PsLHNDMCRksl_CRo#:MRH0CCosL;
CMoH
MRRksl_CRo#:M=R;R
RPkNDC=R:RlMk_osC#n/4;R
RH5VRMCRslnR4RR/=j02RE
CMRRRRPkNDC=R:RDPNk+CRR
4;RMRC8VRH;R
RskC0sPMRNCDk;M
C8kRMlC_OD
D;VOkM0MHFR0oC_8CM_b8C0#E5HRxC:MRH0CCosRR;80CbERR:HCM0o2CsR0sCkRsMHCM0oRCsHP#
NNsHLRDCl_HM#CHxRH:RMo0CC:sR=;Rj
oLCHRM
RMlH_x#HC=R:Rb8C0
E;RVRHRH5#x<CRRb8C0RE20MEC
RRRRMlH_x#HC=R:Rx#HCR;
R8CMR;HV
sRRCs0kMHRlMH_#x
C;CRM8o_C0C_M880CbE
;
O#FM00NMRlMk_D#s_DOCD:#RR0HMCsoCRR:=M_klODCD58N8sH_#xRC,HH#_M0bk,#RH_0Fkb2k0;#

HNoMD#RDLRR:#_08DHFoOC_POs0F58dRF0IMF2RjRR:="jjjj
";0C$bRsR#Dl_0bs_NsRN$HN#Rs$sNRR5j0MFRk#l_sOD_C#DD2VRFR8#0_oDFHPO_CFO0s_58I0H8ERR-4FR8IFM0R;j2
H
#oDMNRb0l_sNsN:$RRD#s_b0l_sNsN
$;#MHoN0DRl8b__sNsN:$RRD#s_b0l_sNsN
$;
0N0skHL0\CR3D#s_VFV#\C0R#:R0MsHo
;
LHCoM0

lNb_s$sN5Rj2<7=Rq;aq
4
z:VRHR8N8sH_I8R0E<c=RRMoCC0sNCR
RRCRLo
HMRRRRRRRRD5#LNs88_8IH0-ERR84RF0IMF2RjRR<=)7q7)R;
RRRRRzRR4:4RRsVFRHHRMRRj05FR8H_I8R0E-R42oCCMsCN0
SSSNs00H0LkC3R\#_sDF#VVCR0\FzVR4R44:NRDLRCDH"#R)"waRH&RMo0CCHs'lCNo5I8_HE802RR&"R7"&MRH0CCosl'HN5oCj&2RR""WRH&RMo0CCHs'lCNo5RH2& R""RR&HCM0o'CsHolNC85N8#s_H2xCR"&RX&"RR0HMCsoC'NHloHC5R4+R2S;
SCSLo
HMRRRRRRRRRRRRz444:)R1p 4n
RRRRRRRRRRRRsbF0NRlbR5
RRRRRRRRRRRRRqRRj>R=RLD#5,j2
RRRRRRRRRRRRRRRRRq4=D>R#4L52R,
RRRRRRRRRRRRRqRR.>R=RLD#5,.2
RRRRRRRRRRRRRRRRRqd=D>R#dL52R,
RRRRRRRRRRRRRBRR >R=R,W 
RRRRRRRRRRRRRRRRiBpRR=>B,pi
RRRRRRRRRRRRRRRR=7R>lR0bs_Ns5N$jH252R,
RRRRRRRRRRRRRTRRRR=>0_lb8s_Ns5N$jH252R
RRRRRRRRRR;R2
RRRRRRRR8CMRMoCC0sNC4Rz4S;
Sz7ma=R<Rb0l_N8_s$sN5;j2
8CMRMoCC0sNC4Rz;z

.H:RV8RN8Is_HE80Rc>RRMoCC0sNCR
RRCRLo
HMRRRRRRRRDR#L<)=Rq)7758dRF0IMF2Rj;R
RRRRRR.Rz.RR:VRFsHMRHR04RFMR5k#l_sOD_C#DD2CRoMNCs0
CRRRRRRRRRRRRRz4..:FRVsRR[HjMRRR0F5I8_HE80R2-4RMoCC0sNCS
SS0N0skHL0\CR3D#s_VFV#\C0RRFVz...RD:RNDLCRRH#"a)w"RR&HCM0o'CsHolNC_58I0H8E&2RR""7RH&RMo0CCHs'lCNo5R5H-2R4*24nR"&RW&"RR0HMCsoC'NHlo[C52RR&"R "&MRH0CCosl'HN5oCo_C0C_M880CbE85N8#s_H,xCR4H*nR22&XR""RR&HCM0o'CsHolNCR5[+2R4;R
RRRRRRRRRRCRLo
HMRRRRRRRRRRRRRRRRz...:)R1pnB4 R
RRRRRRRRRRRRRRFRbsl0RN
b5RRRRRRRRRRRRRRRRq=jR>#RDL25j,R
RRRRRRRRRRRRRR4RqRR=>D5#L4
2,RRRRRRRRRRRRRRRRq=.R>#RDL25.,R
RRRRRRRRRRRRRRdRqRR=>D5#Ld
2,RRRRRRRRRRRRRRRRB= R> RW,R
RRRRRRRRRRRRRRpRBi>R=RiBp,R
RRRRRRRRRRRRRRRR7=0>RlNb_s$sN5-HRR542[
2,RRRRRRRRRRRRRRRRTR46=0>RlNb_s$sN55H2[
2,SSSST>R=Rb0l_N8_s$sN5-HRR542[R2
RRRRRRRRR2RR;R
RRRRRRRRRRRRRRRRRRRR
RRRRRRRRRCRRMo8RCsMCNR0CR.z.4R;
RRRRRCRRMo8RCsMCNR0Cz;..
7SSmRza<0=Rl8b__sNsNO$5F_MPHCM0o5Cs)7q7)85N8Is_HE80R4-RRI8FMR0Fc222;C

Mo8RCsMCNR0Cz
.;
8CMRONsECH0Os0kCCR#D0CO_D#s;



