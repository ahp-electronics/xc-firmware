--
@ER--B$FbsEHo0OR52gR4g-cRRj.jd$R1MHbDO$H0ROQM
R--fN]C8:CsR#//$DMbH0OH$N/lb0DN.Uj4J4.b/blNb#Cs/0N0/LDH/MoC_OFsN/dOs_Nls3_IPyE84
Rf-
-


-----
--
-RN7kDF-bs)0RqIvRHR0E#CCbsCN0R7q7)1 1RsVFRNsC8MRN8sRIH
0C-a-RNCso0RR:pCkOM-0RRBm)qBRd

--DsHLNRs$HCCC;#
kCCRHC#C30D8_FOoH_n44cD3NDk;
#HCRC3CC#_08DHFoOH_#o8MC3DND;#
kCCRHC#C30D8_FOoH_HNs0NE3D
D;DsHLNRs$FNsOdk;
#FCRsdON3OFsNlOFbD3NDC;
M00H$qR)v__)W#RH
RRRRMoCCOsHRR5
RRRRRVRRNDlH$#:R0MsHo=R:RF"MM;C"
RRRRRRRR8IH0:ERR0HMCsoCRR:=(
;RRRRRRRRRNs88I0H8ERR:HCM0oRCs:(=R;RRRRRRRRR--LRHoCkMFoVERF8sRCEb0
RRRRRRRRb8C0:ERR0HMCsoCRR:=RU4.;R
RRRRRRFR8ks0_C:oRRFLFDMCNRR:=V#NDCR;RR-RR-NRE#kRF00bkRosC
RRRRRRRRM8H_osCRL:RFCFDN:MR=NRVD;#CRRRRR-R-R#ENR08NNMRHbRk0s
CoRRRRRRRRs8N8sC_soRR:LDFFCRNM:V=RNCD#;RRRRR--ERN8s8CNR8N8s#C#RosC
RRRRRRRR8IN8ss_C:oRRFLFDMCNRR:=V#NDCRRRR-R-R8ENRHIs0NCR8C8s#s#RCRo
RRRRR2RR;R
RRFRbs50R
RRRRRRRRz7ma:RRR0FkR8#0_oDFHPO_CFO0sH5I8-0E4FR8IFM0R;j2
RRRRRRRR7)q7:)RRRHMR8#0_oDFHPO_CFO0s85N8HsI8-0E4FR8IFM0R;j2
RRRRRRRRh7QR:RRRRHMR8#0_oDFHPO_CFO0sH5I8-0E4FR8IFM0R;j2
RRRRRRRR7Wq7:)RRRHMR8#0_oDFHPO_CFO0s85N8HsI8-0E4FR8IFM0R;j2
RRRRRRRRRW R:RRRRHMR8#0_oDFHRO;RRRRR-R-RHIs0CCRMDNLCFRVsNRslR
RRRRRRpRBiRRR:MRHR0R#8F_Do;HORRRRR-RR-DROFRO	VRFss,NlR8N8s8,RHRM
RRRRRmRRBRpiRH:RM#RR0D8_FOoHRRRRRRRR-F-RbO0RD	FORsVFRk8F0R
RRRRRR;R2
8CMR0CMHR0$)_qv);_W
-
-
R--w#Hs0lRHblDCCNM00MHFR#lk0CRLRDONDRC8NEsOj-
-
ONsECH0Os0kCsRNOREjF)VRq)v__HWR#F
OMN#0MM0RkOl_C#DD_C8CbRR:HCM0oRCs:5=R5b8C0-ERR/42d;.2RRRRRRRRRR--yVRFRIsF#VRFR 7Bdc.XRDOCDM#RCCC88F
OMN#0MM0RkOl_C#DD_8IHCRR:HCM0oRCs:5=R58IH0-ERR/42cR2;RRRRRRRRRR--yVRFRDOFk#lMRRFV7dB .RXcODCD#CRMC88C
b0$CkRF0k_L#$_0bHCR#sRNsRN$5lMk_DOCD8#_CRCb8MFI0jFR,MR5kOl_C#DD_8IHC2*c+8dRF0IMF2RjRRFV#_08DHFoO#;
HNoMDkRF0k_L#RR:F_k0L_k#0C$b;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFRk8F0HR5M0bkRR0F0-sH#00NC
#2#MHoNFDRkC0_MRRRR#:R0D8_FOoH_OPC05FsM_klODCD#C_8C8bRF0IMF2Rj;-RR-MRCNCLD#FRVssR0H0-#N#0C
o#HMRNDIjbC_RCMRRR:#_08DHFoOC_POs0F5lMk_DOCD8#_CRCb8MFI0jFR2R;R-I-RsCH0RNCML#DCRsVFROCNEFRsIVRFRv)qRDOCD##
HNoMDbRICC4_MRRR:0R#8F_Do_HOP0COFMs5kOl_C#DD_C8CbFR8IFM0R;j2R-R-RHIs0CCRMDNLCV#RFCsRNROEsRFIF)VRqOvRC#DD
o#HMRNDHsM_CRoRRRR:#_08DHFoOC_POs0F58IH0dE+RI8FMR0FjR2;RRRRRRRR-k-R#RC80sFRC#oH0RCs7RQh
o#HMRNDW) _ Rt4RRR:#_08DHFoO#;
HNoMDMRH_osC4RRR:0R#8F_Do_HOP0COFIs5HE80+8dRF0IMF2Rj;RRRRH
#oDMNR0Fk_osCR:RRR8#0_oDFHPO_CFO0sH5I8+0EdFR8IFM0R;j2RRRRRRRRRR--k8#CRR0FsHCo#s0CRz7maH
#oDMNR8sN_osCR:RRR8#0_oDFHPO_CFO0s85N8HsI8-0E4FR8IFM0R;j2RRRRRR--k8#CRR0FsHCo#s0CR7)q7#)
HNoMDNRI8C_soRRR:0R#8F_Do_HOP0COFNs58I8sHE80-84RF0IMF2Rj;RRRR-R-RCk#8FR0RosCHC#0sqRW7
7)#MHoNDDRFsI_Ns88R#:R0D8_FOoH_OPC05FscFR8IFM0R;j2RRRRRRRRRRRRR-RR-NRs8R8sL#H0RbHMk00RFqR)vCRODRD#5L6RHR0#skCJH8sC2H
#oDMNRIDF_8IN8:sRR8#0_oDFHPO_CFO0sR5c8MFI0jFR2R;RRRRRRRRRRRRRRR--I8N8sHRL0H#RM0bkRR0F)RqvODCD#6R5R0LH#CRsJskHC
820C$bRb0l_8N8s$_0bHCR#sRNsRN$5lMk_DOCD8#_CRCb8MFI0jFR2VRFR8#0_oDFHPO_CFO0sgR5RI8FMR0Fj
2;#MHoN0DRlNb_8R8sR0:RlNb_8_8s0C$b;L

CMoH
R
RR-R-RRQVNs88I0H8ERR<6#RN#MHoR''jRR0Fk#MkCL8RH
0#RRRRzR4R:VRHR85N8HsI8R0E=2R4RMoCC0sNCR
RRRRRRFRDIN_s8R8s<"=Rjjjj"RR&s_N8s5Coj
2;RRRRRRRRD_FII8N8s=R<Rj"jjRj"&NRI8C_so25j;R
RRMRC8CRoMNCs0zCR4R;
RzRR.:RRRRHV58N8s8IH0=ERRR.2oCCMsCN0
RRRRRRRRIDF_8sN8<sR=jR"jRj"&NRs8C_soR548MFI0jFR2R;
RRRRRDRRFII_Ns88RR<="jjj"RR&I_N8s5Co4FR8IFM0R;j2
RRRR8CMRMoCC0sNC.Rz;R
RRdRzRRR:H5VRNs88I0H8ERR=do2RCsMCN
0CRRRRRRRRD_FIs8N8s=R<Rj"j"RR&s_N8s5Co.FR8IFM0R;j2
RRRRRRRRIDF_8IN8<sR=jR"j&"RR8IN_osC58.RF0IMF2Rj;R
RRMRC8CRoMNCs0zCRdR;
RzRRc:RRRRHV58N8s8IH0=ERRRc2oCCMsCN0
RRRRRRRRIDF_8sN8<sR=jR''RR&s_N8s5CodFR8IFM0R;j2
RRRRRRRRIDF_8IN8<sR=jR''RR&I_N8s5CodFR8IFM0R;j2
RRRR8CMRMoCC0sNCcRz;R
RR6RzRRR:H5VRNs88I0H8ERR>co2RCsMCN
0CRRRRRRRRD_FIs8N8s=R<R8sN_osC58cRF0IMF2Rj;R
RRRRRRFRDIN_I8R8s<I=RNs8_Cco5RI8FMR0Fj
2;RRRRCRM8oCCMsCN0R;z6
R
RR-R-RRQV5M8H_osC2CRso0H#C7sRQkhR#oHMRiBp
RRRRRznRH:RV8R5HsM_CRo2oCCMsCN0
RRRRRRRRFbsO#C#Rp5Bi7,RQRh2LHCoMR
RRRRRRRRRRVRHRp5BiRR='R4'NRM8B'piCMPC002RE
CMRRRRRRRRRRRRRRRRHsM_C<oR="R5jjjj"RR&72Qh;R
RRRRRRRRRRMRC8VRH;R
RRRRRRMRC8sRbF#OC#R;
RCRRMo8RCsMCNR0Cz
n;RRRRzR(R:VRHRF5M0HR8MC_soo2RCsMCN
0CRRRRRRRRRRRRHsM_C<oR="R5jjjj"RR&72Qh;R
RRMRC8CRoMNCs0zCR(
;
RRRR-Q-RVsR5Ns88_osC2CRso0H#C)sRq)77RHk#MBoRpRi
RzRR4RjR:VRHRN5s8_8ss2CoRMoCC0sNCR
RRRRRRsRbF#OC#mR5B,piR7)q7R)2LHCoMR
RRRRRRRRRRVRHRB5mp=iRR''4R8NMRpmBiP'CC2M0RC0EMR
RRRRRRRRRRRRRRNRs8C_so=R<R7)q7N)58I8sHE80-84RF0IMF2Rj;R
RRRRRRRRRRMRC8VRH;R
RRRRRRMRC8sRbF#OC#R;
RCRRMo8RCsMCNR0Cz;4j
RRRR4z4RH:RVMR5Fs0RNs88_osC2CRoMNCs0RC
RRRRRRRRRsRRNs8_C<oR=qR)757)Ns88I0H8ER-48MFI0jFR2R;
RCRRMo8RCsMCNR0Cz;44
RRRRRRRRR
RR-R-RRQV58IN8ss_CRo2sHCo#s0CR7Wq7k)R#oHMRiBp
RRRR.z4RRR:H5VRI8N8sC_soo2RCsMCN
0CRRRRRRRRbOsFCR##5iBp,qRW727)RoLCHRM
RRRRRRRRRHRRVBR5p=iRR''4R8NMRiBp'CCPMR020MEC
RRRRRRRRRRRRRRRR8IN_osCRR<=W7q7)85N8HsI8-0E4FR8IFM0R;j2
RRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMRFbsO#C#;R
RRMRC8CRoMNCs0zCR4
.;RRRRzR4d:VRHRF5M0NRI8_8ss2CoRMoCC0sNCR
RRRRRRRRRRNRI8C_so=R<R7Wq7
);RRRRCRM8oCCMsCN0Rdz4;R

R-RR-CRtMNCs00CRE)CRqOvRC#DDR8NMRD#CCRO0DHFoOR
RR4RzcRR:VRFsHMRHRlMk_DOCD8#_CRCb8MFI0jFRRMoCC0sNCR
RR-R-RHAkDF8Rkk0b0MRCNCLDRD#CCRO0DHFoOR
RRRRRR-R-RRQV58N8s8IH0>ERR246RMON'k0R#NCRRQ1pBCRODRD
RRRRRmRR R4n:VRHR85N8HsI8R0E>6R42CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_M25HRR<='R4'IMECRN5s8C_so85N8HsI8-0E4FR8IFM0RR62=2RHR#CDCjR''R;
RRRRRCRRMo8RCsMCNR0Cmn 4;R
RRRRRR-R-RRQV58N8s8IH0>ERRR62qRh758N8s8IH0<ER=6R42#RkNRRN1BpQRDOCDR
RRRRRR Rm4:6RRRHV58N8s8IH0=ERR246RMoCC0sNCR
RRRRRRRRRRRRRRlR0b8_N8Hs52R5g8MFI0jFR2=R<Rahm5MOFP0_#8F_Do_HOP0COFHs5,jR42X2Rms)RNs8_CNo58I8sHE80-84RF0IMF2R6;R
RRRRRRRRRRRRRRqR1h47_6RR:17qh4bjRFRs0lRNb5=qR>lR0b8_N8Hs5225j,RRA=0>RlNb_858sH4252B,RRR=>0_lbNs8855H2.R2,7>R=Rb0l_8N8s25H5,d2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR >R=Rb0l_8N8s25H5,c2R=wR>lR0b8_N8Hs52256,RRt=0>RlNb_858sHn252],RRR=>0_lbNs8855H2(R2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRQ>R=Rb0l_8N8s25H5,U2R=KR>lR0b8_N8Hs5225g,RRZ=F>RkC0_M25H2R;
RRRRRCRRMo8RCsMCNR0Cm6 4;R
RRRRRR Rm4:cRRRHV58N8s8IH0=ERR24cRMoCC0sNCR
RRRRRRRRRRRRRRlR0b8_N8Hs52R5U8MFI0jFR2=R<Rahm5MOFP0_#8F_Do_HOP0COFHs5,2Rg2mRX)NRs8C_so85N8HsI8-0E4FR8IFM0R;62
RRRRRRRRRRRRRRRRh1q7c_4R1:Rq4h7jFRbsl0RN5bRq>R=Rb0l_8N8s25H5,j2R=AR>lR0b8_N8Hs52254,RRB=0>RlNb_858sH.2527,RRR=>0_lbNs8855H2d
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR RRRR=>0_lbNs8855H2cR2,w>R=Rb0l_8N8s25H5,62R=tR>lR0b8_N8Hs5225n,RR]=0>RlNb_858sH(252
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRQRRRR=>0_lbNs8855H2UR2,K>R=R''4,RRZ=F>RkC0_M25H2R;
RRRRRCRRMo8RCsMCNR0Cmc 4;R
RRRRRR Rm4:dRRRHV58N8s8IH0=ERR24dRMoCC0sNCR
RRRRRRRRRRRRRRlR0b8_N8Hs52R5(8MFI0jFR2=R<Rahm5MOFP0_#8F_Do_HOP0COFHs5,2RU2mRX)NRs8C_so85N8HsI8-0E4FR8IFM0R;62
RRRRRRRRRRRRRRRRh1q7d_4R1:RqUh7RFRbsl0RN5bRq>R=Rb0l_8N8s25H5,j2R=AR>lR0b8_N8Hs52254,RRB=0>RlNb_858sH.2527,RRR=>0_lbNs8855H2d
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR RRRR=>0_lbNs8855H2cR2,w>R=Rb0l_8N8s25H5,62R=tR>lR0b8_N8Hs5225n,RR]=0>RlNb_858sH(252
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRZRRRR=>F_k0CHM52
2;RRRRRRRRCRM8oCCMsCN0R4m dR;
RRRRRmRR R4.:VRHR85N8HsI8R0E=.R42CRoMNCs0RC
RRRRRRRRRRRRR0RRlNb_858sHn25RI8FMR0Fj<2R=mRhaF5OM#P_0D8_FOoH_OPC05FsH(,R2X2Rms)RNs8_CNo58I8sHE80-84RF0IMF2R6;R
RRRRRRRRRRRRRRqR1h47_.RR:17qhUbRRFRs0lRNb5=qR>lR0b8_N8Hs5225j,RRA=0>RlNb_858sH4252B,RRR=>0_lbNs8855H2.R2,7>R=Rb0l_8N8s25H5,d2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR >R=Rb0l_8N8s25H5,c2R=wR>lR0b8_N8Hs52256,RRt=0>RlNb_858sHn252],RRR=>',4'RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR=ZR>kRF0M_C52H2;R
RRRRRRMRC8CRoMNCs0mCR ;4.
RRRRRRRR4m 4RR:H5VRNs88I0H8ERR=4R42oCCMsCN0
RRRRRRRRRRRRRRRRb0l_8N8s25H586RF0IMF2RjRR<=h5maOPFM_8#0_oDFHPO_CFO0s,5HR2n2R)XmR8sN_osC58N8s8IH04E-RI8FMR0F6
2;RRRRRRRRRRRRRRRR17qh_R44:qR1hR7nRsbF0NRlbqR5RR=>0_lbNs8855H2jR2,A>R=Rb0l_8N8s25H5,42R=BR>lR0b8_N8Hs5225.,RR7=0>RlNb_858sHd252R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR =0>RlNb_858sHc252w,RRR=>0_lbNs8855H26R2,Z>R=R0Fk_5CMH;22
RRRRRRRR8CMRMoCC0sNC Rm4
4;RRRRRRRRmj 4RH:RVNR58I8sHE80R4=Rjo2RCsMCN
0CRRRRRRRRRRRRRRRR0_lbNs8855H2cFR8IFM0RRj2<h=RmOa5F_MP#_08DHFoOC_POs0F5RH,6R22XRm)s_N8s5CoNs88I0H8ER-48MFI06FR2R;
RRRRRRRRRRRRR1RRq_h74:jRRh1q7RnRb0FsRblNRR5q=0>RlNb_858sHj252A,RRR=>0_lbNs8855H24R2,B>R=Rb0l_8N8s25H5,.2R=7R>lR0b8_N8Hs5225d,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR= R>lR0b8_N8Hs5225c,RRw='>R4R',Z>R=R0Fk_5CMH;22
RRRRRRRR8CMRMoCC0sNC Rm4
j;RRRRRRRRmR gRH:RVNR58I8sHE80Rg=R2CRoMNCs0RC
RRRRRRRRRRRRR0RRlNb_858sHd25RI8FMR0Fj<2R=mRhaF5OM#P_0D8_FOoH_OPC05FsHc,R2X2Rms)RNs8_CNo58I8sHE80-84RF0IMF2R6;R
RRRRRRRRRRRRRRqR1hg7_R1:Rqch7RbRRFRs0lRNb5=qR>lR0b8_N8Hs5225j,RRA=0>RlNb_858sH4252B,RRR=>0_lbNs8855H2.R2,7>R=Rb0l_8N8s25H5,d2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRZ>R=R0Fk_5CMH;22
RRRRRRRR8CMRMoCC0sNC RmgR;
RRRRRmRR RUR:VRHR85N8HsI8R0E=2RURMoCC0sNCR
RRRRRRRRRRRRRRlR0b8_N8Hs52R5.8MFI0jFR2=R<Rahm5MOFP0_#8F_Do_HOP0COFHs5,2Rd2mRX)NRs8C_so85N8HsI8-0E4FR8IFM0R;62
RRRRRRRRRRRRRRRRh1q7R_U:qR1hR7cRFRbsl0RN5bRq>R=Rb0l_8N8s25H5,j2R=AR>lR0b8_N8Hs52254,RRB=0>RlNb_858sH.2527,RRR=>',4'
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRZ>R=R0Fk_5CMH;22
RRRRRRRR8CMRMoCC0sNC RmUR;
RRRRRmRR R(R:VRHR85N8HsI8R0E=2R(RMoCC0sNCR
RRRRRRRRRRRRRRlR0b8_N8Hs52R548MFI0jFR2=R<Rahm5MOFP0_#8F_Do_HOP0COFHs5,2R.2mRX)NRs8C_so85N8HsI8-0E4FR8IFM0R;62
RRRRRRRRRRRRRRRRh1q7R_(:qR1hR7.RFRbsl0RN5bRq>R=Rb0l_8N8s25H5,j2R=AR>lR0b8_N8Hs52254,RRZ=F>RkC0_M25H2R;
RRRRRCRRMo8RCsMCNR0Cm; (
RRRRRRRRnm RRR:H5VRNs88I0H8ERR=no2RCsMCN
0CRRRRRRRRRRRRRRRRF_k0CHM52=R<R''4RCIEMsR5Ns8_C6o52RR=OPFM_8#0_oDFHPO_CFO0s,5H4j252C2RDR#C';j'
RRRRRRRR8CMRMoCC0sNC RmnR;
R-RR-VRQR85N8HsI8R0E<6=R2FRMR0FkbRk0CLMND#CRCODC0FRDoRHOM8CCCR8
RRRRRmRR :6RRRHV58N8s8IH0<ER=2R6RMoCC0sNCR
RRRRRRRRRRRRRRkRF0M_C5RH2<'=R4
';RRRRRRRRCRM8oCCMsCN0R6m ;R

R-RR-VRQR85N8HsI8R0E>2RgRCk#R WujFR0RO8CFR8CNs88CR##L#H0R0nREksFogERR8NMR Wu4FR0RO8CFR8CL#H0RR4j+R
RRRRRR RW4:jRRRHV58N8s8IH0>ERRRg2oCCMsCN0
RRRRRRRRRRRRRRRRCIbjM_C5RH2<'=R4I'RERCM58IN_osC58URF0IMF2R6RO=RF_MP#_08DHFoOC_POs0F5.H,jd25RI8FMR0FjR22CCD#R''j;R
RRRRRRRRRRRRRRbRICC4_M25HRR<='R4'IMECRN5I8C_so85N8HsI8-0E4FR8IFM0RRg2=FROM#P_0D8_FOoH_OPC05FsHj,.285N8HsI8-0EnFR8IFM0R2c2R#CDCjR''R;
RRRRRRRRRCRRMo8RCsMCNR0CWj 4;R
RR-R-RRQV58N8s8IH0=ERRFURs2RgRCk#R WujFR0RO8CFR8CNs88CR##L#H0R0nREksFogER
RRRRRRRRgW RRR:H5VR58N8s8IH0=ERRRU2m5)RNs88I0H8ERR=gR22oCCMsCN0
RRRRRRRRRRRRRRRRCIbjM_C5RH2<'=R4I'RERCM58IN_osC58N8s8IH04E-RI8FMR0F6=2RRRH2CCD#R''j;R
RRRRRRRRRRRRRRbRICC4_M25HRR<=';4'
RRRRRRRRRRRR8CMRMoCC0sNC RWgR;
R-RR-VRQR85N8HsI8R0E=2R(RCk#R WujFR0RO8CFR8C0RECnR0ENs88CR##LRH0&uRW 04RFCR8OCF8RC0ERE(0R8N8s#C#R0LH
RRRRRRRR(W RRR:H5VRNs88I0H8ERR=(o2RCsMCN
0CRRRRRRRRRRRRRRRRIjbC_5CMH<2R=4R''ERIC5MRI_N8s5Co6=2RRMOFP0_#8F_Do_HOP0COFHs5,5.2jR22CCD#R''j;R
RRRRRRRRRRRRRRbRICC4_M25HRR<='R4'IMECRN5I8C_so25nRO=RF_MP#_08DHFoOC_POs0F5.H,22542DRC#'CRj
';RRRRRRRRCRM8oCCMsCN0R(W ;R
RR-R-RRQV58N8s8IH0=ERRRn2kR#CWju RR0F8FCO80CREnCR0NER8C8s#L#RHR0
RRRRRWRR RnR:VRHR85N8HsI8R0E=2RnRMoCC0sNCR
RRRRRRRRRRRRRRbRICCj_M25HRR<='R4'IMECRN5I8C_so256RO=RF_MP#_08DHFoOC_POs0F54H,225j2DRC#'CRj
';RRRRRRRRRRRRRRRRI4bC_5CMH<2R=4R''R;
RRRRRCRRMo8RCsMCNR0CW; n
RRRRR--Q5VRNs88I0H8E=R<RR62MIFRsCH0RNCMLRDC#CCDOD0RFOoHRCMC8
C8RRRRRRRRWR 6RH:RVNR58I8sHE80RR<=6o2RCsMCN
0CRRRRRRRRRRRRRRRRIjbC_5CMH<2R=4R''R;
RRRRRRRRRRRRRIRRb_C4CHM52=R<R''4;R
RRRRRRMRC8CRoMNCs0WCR 
6;
RRRR8CMRMoCC0sNC4Rzc
;
RRRRbOsFCR##5iBp,QR7hL2RCMoH
RRRRRRRH5VRBRpi=4R''MRN8pRBiP'CC2M0RC0EMR
RRRRRRRRRR_HMs4CoRR<=HsM_C
o;RRRRRRRRRWRR  _)t<4R= RW;R
RRRRRR8CMR;HV
RRRR8CMRFbsO#C#;R

RzRR.:6RRRHV50MFRk8F0C_soo2RCsMCN
0CRRRRRRRRz44(:sRbF#OC#WR5  _)tR4,)7q7)W,Rq)77,MRH_osC4F,Rks0_C
o2RRRRRRRRLHCoMR
RRRRRRRRRRVRHRW55  _)t=4RR''42MRN8)R5q)77RW=Rq)77202RE
CMRRRRRRRRRRRRRRRR7amzRR<=HsM_C5o4I0H8ER-48MFI0jFR2R;
RRRRRRRRRCRRD
#CRRRRRRRRRRRRRRRR7amzRR<=F_k0s5CoI0H8ER-48MFI0jFR2R;
RRRRRRRRRCRRMH8RVR;
RRRRRCRRMb8RsCFO#z#R4;(4
RRRR8CMRMoCC0sNC.Rz6
;
RRRRzRdjRH:RV8R5F_k0s2CoRMoCC0sNCR
RRRRRRsRbF#OC#mR5B,piR0Fk_osC2CRLo
HMRRRRRRRRRRRRH5VRmiBpR'=R4N'RMm8RB'piCMPC002RE
CMRRRRRRRRRRRRRRRR7amzRR<=F_k0s5CoI0H8ER-48MFI0jFR2R;
RRRRRRRRRCRRMH8RVR;
RRRRRCRRMb8RsCFO#
#;RRRRCRM8oCCMsCN0Rjzd;R

R-RR-MRtC0sNCER0CqR)vCRODRD#IEH0RH0s-N#00
C#RRRRzR46:FRVsRRHHMMRkOl_C#DD_C8CbFR8IFM0RojRCsMCN
0CRRRRRRRRzR4(:FRVsRR[HMMRkOl_C#DD_8IHCFR8IFM0RojRCsMCN
0CRRRRRRRRRRRRzv)q:BR7 Xd.cRR
RRRRRRRRRRRRRbRRFRs0lRNb5j7QRR=>HsM_C5o5[2*c27,RQ=4R>MRH_osC5*5[c42+27,RQ=.R>MRH_osC5*5[c.2+27,RQ=dR>MRH_osC5*5[cd2+2R,
RRRRRRRRRRRRRRRRRRRRRRRRR7Wqj>R=RIDF_8IN8js52W,RqR74=D>RFII_Ns885,42R7Wq.>R=RIDF_8IN8.s52W,RqR7d=D>RFII_Ns885,d2R7Wqc>R=RIDF_8IN8cs52R,
RRRRRRRRRRRRRRRRRRRRRRRRR7)qj>R=RIDF_8sN8js52),RqR74=D>RFsI_Ns885,42R7)q.>R=RIDF_8sN8.s52),RqR7d=D>RFsI_Ns885,d2R7)qc>R=RIDF_8sN8cs52-,
-RRRRRRRRRRRRRRRRRRRRRRRRWRR)R h=W>R W,RuR j=I>Rb_CjCHM52W,RuR 4=I>Rb_C4CHM52B,Ri>R=Rahm5iBp2
,RRRRRRRRRRRRRRRRRRRRRRRRRR)RW =hR> RW,uRW =jR>bRICCj_M25H,uRW =4R>bRICC4_M25H,iRBRR=>B,piRR
RRRRRRRRRRRRRRRRRRRRRRRRR7Rmj=F>RkL0_kH#5,*5[c,22R47mRR=>F_k0L5k#H[,5*+c24R2,7Rm.=F>RkL0_kH#5,*5[c.2+27,Rm=dR>kRF0k_L#,5H5c[*22+d2R;
RRRRRRRRRRRRRFRRks0_C5o5[2*c2=R<R0Fk_#Lk55H,[2*c2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C5o5[2*c+R42<F=RkL0_kH#5,*5[c42+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C5o5[2*c+R.2<F=RkL0_kH#5,*5[c.2+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C5o5[2*c+Rd2<F=RkL0_kH#5,*5[cd2+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRCRRMo8RCsMCNR0Cz;4(
RRRR8CMRMoCC0sNC4Rz6
;
-R-RzR.U:VRHRF58ks0_CRo2oCCMsCN0
R--RRRRRzRR4:nRRsVFRHHRMkRMlC_OD_D#8bCCRI8FMR0FjCRoMNCs0-C
-RRRRRRRRUz4RV:RF[sRRRHMM_klODCD#H_I88CRF0IMFRRjoCCMsCN0
R--RRRRRRRRRzRR):qvR 7Bdc.XR-
-RRRRRRRRRRRRRRRRb0FsRblNRQ57j>R=R_HMs5Co5c[*2R2,7RQ4=H>RMC_so[55*+c24R2,7RQ.=H>RMC_so[55*+c2.R2,7RQd=H>RMC_so[55*+c2d
2,-R-RRRRRRRRRRRRRRRRRRRRRRRRRWjq7RR=>D_FII8N8s25j,qRW7=4R>FRDIN_I858s4R2,W.q7RR=>D_FII8N8s25.,qRW7=dR>FRDIN_I858sdR2,Wcq7RR=>D_FII8N8s25c,-
-RRRRRRRRRRRRRRRRRRRRRRRRRqR)7=jR>FRDIN_s858sjR2,)4q7RR=>D_FIs8N8s254,qR)7=.R>FRDIN_s858s.R2,)dq7RR=>D_FIs8N8s25d,qR)7=cR>FRDIN_s858sc
2,-R-RRRRRRRRRRRRRRRRRRRRRRRRRWh) RR=>WR ,Wju RR=>IjbC_5CMHR2,W4u RR=>I4bC_5CMHR2,B=iR>mRhap5BiR2,
R--RRRRRRRRRRRRRRRRRRRRRRRRRmT7j>R=R0Fk_#Lk55H,[2*c2T,R7Rm4=F>RkL0_kH#5,*5[c42+2T,R7Rm.=F>RkL0_kH#5,*5[c.2+2T,R7Rmd=F>RkL0_kH#5,*5[cd2+2
2;---
-RRRRRRRRRRRRFRRks0_C5o5[2*c2=R<R0Fk_#Lk55H,[2*c2ERIC5MRF_k0CHM52RR='24'R#CDCZR''-;
-RRRRRRRRRRRRRRRR0Fk_osC5*5[c42+2=R<R0Fk_#Lk55H,[2*c+R42IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
R--RRRRRRRRRRRRRFRRks0_C5o5[2*c+R.2<F=RkL0_kH#5,*5[c.2+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''-;
-RRRRRRRRRRRRRRRR0Fk_osC5*5[cd2+2=R<R0Fk_#Lk55H,[2*c+Rd2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
R--RRRRRRRRRCRRMo8RCsMCNR0Cz;4U
R--RRRRRMRC8CRoMNCs0zCR4
n;-R-RRMRC8CRoMNCs0zCR.
U;
R--RRRRRRkU:VRHRF58ks0_CRo2oCCMsCN0
R--RRRRRz7ma=R<R0Fk_osC58IH04E-RI8FMR0Fj
2;-R-RCRM8oCCMsCN0R;kU
RRRRRRRRM
C8sRNO0EHCkO0sNCRsjOE;



