--
@ER--B$FbsEHo0OR52gR4g-cRRj.jd$R1MHbDO$H0ROQM
R--fN]C8:CsR#//$DMbH0OH$N/lb0DN.Uj4J4.b/blNb#Cs/DGHH/MGD/HLoCCMs/HOo_CMoCCMs/HOs_Nls3_IPyE84
Rf-
-
----- RBpXpR)dqv.7X4R----D-
HNLssH$RC;CC
Ck#RCHCC03#8F_Do_HO4c4n3DND;#
kCCRHC#C30D8_FOoH_o#HM3C8N;DD
LDHs$NsRHkM#;Hl
Ck#RHkM#3HlPlOFbCFMM30#N;DD
M
C0$H0RqX)vXd.4H7R#R
Rb0FsRR5
RRRRR7RRuRmRRF:Rk#0R0k8_DHFoOR;RRRRRRRR
RRRRR1RRuRmRRF:Rk#0R0k8_DHFoO
;
RRRRRRRRqRjRRRR:H#MR0k8_DHFoOR;
RRRRRqRR4RRRRH:RM0R#8D_kFOoH;R
RRRRRR.RqRRRR:MRHR8#0_FkDo;HO
RRRRRRRRRqdR:RRRRHM#_08koDFH
O;RRRRRRRRqRcRRRR:H#MR0k8_DHFoOR;
RRRRR7RRRRRRRH:RM0R#8D_kFOoH;R
RRRRRRuR7)Rqj:MRHR8#0_FkDo;HO
RRRRRRRR)7uq:4RRRHM#_08koDFH
O;RRRRRRRR7qu).RR:H#MR0k8_DHFoOR;
RRRRR7RRud)qRH:RM0R#8D_kFOoH;R
RRRRRRuR7)Rqc:MRHR8#0_FkDo;HO
RRRRRRRRpWBi:RRRRHM#_08koDFHRO;RRRRR
RRRRRRRRRRWR RRRR:H#MR0k8_DHFoOR
RRRRRRR2;RM
C8)RXq.vdX;47
ONsECH0Os0kC)RXq.vdX_47eVRFRqX)vXd.4H7R#R
RSo#HMRNDI,CjR4IC,FR#j#,RFR4,8,FjR48F:0R#8F_Do;HO
oLCHSM
7Rum<8=RFIjRERCM5)7uq=cRR''j2DRC#8CRF
4;Sm1uRR<=#RFjIMECRc5qR'=RjR'2CCD#R4#F;I
SC<jR= RWR8NMRF5M0cRq2S;
IRC4<W=R MRN8cRq;S
Rz:jRRv)q44nX7RR
RRRRRRRRRRRRRbRRFRs0lRNb5=7R>,R7RRqj=q>Rjq,R4>R=R,q4RRq.=q>R.q,Rd>R=R,qd
SRSS)7uq=jR>uR7),qjR)7uq=4R>uR7),q4R)7uq=.R>uR7),q.R)7uq=dR>uR7),qdRS
SSRW =I>RCRj,WiBpRR=>WiBp,uR7m>R=Rj8F,uR1m>R=Rj#F2R;
SRz4:qR)vX4n4
7RRRRRRRRRRRRRRRRRb0FsRblNRR57=7>R,jRqRR=>qRj,q=4R>4Rq,.RqRR=>qR.,q=dR>dRq,S
RSuS7)Rqj=7>Ruj)q,uR7)Rq4=7>Ru4)q,uR7)Rq.=7>Ru.)q,uR7)Rqd=7>Rud)q,SR
S SWRR=>I,C4RpWBi>R=RpWBi7,Ru=mR>FR841,Ru=mR>FR#4
2;CRM8Xv)qd4.X7;_e
-
--R--Bp pRqX)vXnc4-7R----
LDHs$NsRCHCCk;
#HCRC3CC#_08DHFoO4_4nNc3D
D;kR#CHCCC38#0_oDFH#O_HCoM8D3NDD;
HNLssk$RMHH#lk;
#kCRMHH#lO3PFFlbM0CM#D3ND
;
CHM00X$R)nqvc7X4R
H#RFRbs50R
RRRRRRRRm7uR:RRR0FkR8#0_FkDo;HORRRRRRRR
RRRRRRRRm1uR:RRR0FkR8#0_FkDo;HO
R
RRRRRRjRqRRRR:MRHR8#0_FkDo;HO
RRRRRRRRRq4R:RRRRHM#_08koDFH
O;RRRRRRRRqR.RRRR:H#MR0k8_DHFoOR;
RRRRRqRRdRRRRH:RM0R#8D_kFOoH;R
RRRRRRcRqRRRR:MRHR8#0_FkDo;HO
RRRRRRRRRq6R:RRRRHM#_08koDFH
O;RRRRRRRR7RRRRRR:H#MR0k8_DHFoOR;
RRRRR7RRuj)qRH:RM0R#8D_kFOoH;R
RRRRRRuR7)Rq4:MRHR8#0_FkDo;HO
RRRRRRRR)7uq:.RRRHM#_08koDFH
O;RRRRRRRR7qu)dRR:H#MR0k8_DHFoOR;
RRRRR7RRuc)qRH:RM0R#8D_kFOoH;R
RRRRRRuR7)Rq6:MRHR8#0_FkDo;HO
RRRRRRRRpWBi:RRRRHM#_08koDFHRO;RRRRR
RRRRRRRRRRWR RRRR:H#MR0k8_DHFoOR
RRRRRRR2;RM
C8)RXqcvnX;47
ONsECH0Os0kC)RXqcvnX_47eVRFRqX)vXnc4H7R#R
RSo#HMRNDI,CjR4IC,CRI.I,RCRd,#,FjR4#F,FR#.#,RFRd,8,FjR48F,FR8.8,RFRd:#_08DHFoOL;
CMoH
uS7m=R<RFR8jERIC5MR7qu)6RR='Rj'NRM87qu)cRR='2j'R#CDCSR
S48FRCIEM7R5u6)qR'=RjN'RM78Ruc)qR'=R4R'2CCD#RS
S8RF.IMECRu57)Rq6=4R''MRN8uR7)Rqc=jR''C2RDR#C
8SSF
d;Sm1uRR<=Rj#FRCIEMqR56RR='Rj'NRM8q=cRR''j2DRC#
CRSFS#4ERIC5MRq=6RR''jR8NMRRqc=4R''C2RDR#C
#SSFI.RERCM5Rq6=4R''MRN8cRqR'=RjR'2CCD#RS
S#;Fd
CSIj=R<RRW NRM850MFR2q6R8NMRF5M0cRq2S;
IRC4<W=R MRN8MR5Fq0R6N2RMq8RcS;
IRC.<W=R MRN86RqR8NMRF5M0cRq2S;
IRCd<W=R MRN86RqR8NMR;qc
zRSjRR:)4qvn7X4RR
RRRRRRRRRRRRRRFRbsl0RN5bR7>R=RR7,q=jR>jRq,4RqRR=>qR4,q=.R>.Rq,dRqRR=>q
d,RSSS7qu)j>R=R)7uqRj,7qu)4>R=R)7uqR4,7qu).>R=R)7uqR.,7qu)d>R=R)7uqRd,
SSSW= R>CRIjW,RBRpi=W>RB,piRm7uRR=>8,FjRm1uRR=>#2Fj;S
Rz:4RRv)q44nX7RR
RRRRRRRRRRRRRbRRFRs0lRNb5=7R>,R7RRqj=q>Rjq,R4>R=R,q4RRq.=q>R.q,Rd>R=R,qd
SRSS)7uq=jR>uR7),qjR)7uq=4R>uR7),q4R)7uq=.R>uR7),q.R)7uq=dR>uR7),qdRS
SSRW =I>RCR4,WiBpRR=>WiBp,uR7m>R=R48F,uR1m>R=R4#F2R;
SRz.:qR)vX4n4
7RRRRRRRRRRRRRRRRRb0FsRblNRR57=7>R,jRqRR=>qRj,q=4R>4Rq,.RqRR=>qR.,q=dR>dRq,S
RSuS7)Rqj=7>Ruj)q,uR7)Rq4=7>Ru4)q,uR7)Rq.=7>Ru.)q,uR7)Rqd=7>Rud)q,SR
S SWRR=>I,C.RpWBi>R=RpWBi7,Ru=mR>FR8.1,Ru=mR>FR#.
2;RdSzR):Rqnv4XR47
RRRRRRRRRRRRRRRRsbF0NRlb7R5RR=>7q,Rj>R=R,qjRRq4=q>R4q,R.>R=R,q.RRqd=q>RdR,
S7SSuj)qRR=>7qu)j7,Ru4)qRR=>7qu)47,Ru.)qRR=>7qu).7,Rud)qRR=>7qu)d
,RSWSS >R=RdIC,BRWp=iR>BRWpRi,7Rum=8>RFRd,1Rum=#>RF;d2
8CMRqX)vXnc4e7_;-

--
-
R--1bHlD)CRqIvRHR0E#oHMDqCR7 7)1V1RFLsRFR0Es8CNR8NMRHIs0-C
-NRas0oCRX:RHMDHG-
-
H
DLssN$CRHC
C;kR#CHCCC38#0_oDFH4O_43ncN;DD
Ck#RCHCC03#8F_Do_HO#MHoCN83D
D;DsHLNRs$k#MHH
l;kR#Ck#MHHPl3ObFlFMMC0N#3D
D;CHM00)$Rq)v__HWR#o
SCsMCH5OR
RSRRNRVl$HDR#:R0MsHo=R:RF"MM;C"
ISSHE80RH:RMo0CC:sR=;R4RS
SNs88I0H8ERR:HCM0oRCs:n=R;RRRRRRRRR--LRHoCkMFoVERF8sRCEb0
8SSCEb0RH:RMo0CC:sR=URc;S
S80Fk_osCRL:RFCFDN:MR=NRVD;#CRRRRR-R-R#ENR0FkbRk0s
CoSHS8MC_soRR:LDFFCRNM:V=RNCD#;RRRRRRRRR--ERN#8NN0RbHMks0RCSo
S8sN8ss_C:oRRFLFDMCNRR:=V#NDCR;RRRRR-E-RNs#RCRN8Ns88CR##s
CoSNSI8_8ssRCo:FRLFNDCM:RR=NRVDR#CRRRRRR--ERN#I0sHC8RN8#sC#CRsoS
S2S;
b0FsRS5
Sz7maF:Rk#0R0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2S;
S7)q7:)RRRHM#_08DHFoOC_POs0F58N8s8IH04E-RI8FMR0Fj
2;SQS7h:RRRRHM#_08DHFoOC_POs0F58IH04E-RI8FMR0Fj
2;SqSW7R7):MRHR8#0_oDFHPO_CFO0s85N8HsI8-0E4FR8IFM0R;j2
WSS :RRRRHM#_08DHFoOR;RRRRRRR--I0sHCMRCNCLDRsVFRlsN
BSSp:iRRRHM#_08DHFoOR;RRRRRRR--OODF	FRVsNRslN,R8,8sRM8H
mSSBRpi:MRHR8#0_oDFHRORRRRRRR--FRb0OODF	FRVs_RI80Fk
2SS;M
C8MRC0$H0Rv)q_W)_;-

--
-RswH#H0RlCbDl0CMNF0HMkRl#L0RCNROD8DCRONsE-j
-s
NO0EHCkO0sLCRD	FO_lsNRRFV)_qv)R_WHO#
FFlbM0CMRqX)vXd.4R7RRsbF0
R5RRRRRRRR7RumRRR:FRk0#_08koDFHRO;RRRRR
RRRRRRRRRR1RumRRR:FRk0#_08koDFH
O;
RRRRRRRRRqjR:RRRRHM#_08koDFH
O;RRRRRRRRqR4RRRR:H#MR0k8_DHFoOR;
RRRRRqRR.RRRRH:RM0R#8D_kFOoH;R
RRRRRRdRqRRRR:MRHR8#0_FkDo;HO
RRRRRRRRRqcR:RRRRHM#_08koDFH
O;RRRRRRRR7RRRRRR:H#MR0k8_DHFoOR;
RRRRR7RRuj)qRH:RM0R#8D_kFOoH;R
RRRRRRuR7)Rq4:MRHR8#0_FkDo;HO
RRRRRRRR)7uq:.RRRHM#_08koDFH
O;RRRRRRRR7qu)dRR:H#MR0k8_DHFoOR;
RRRRR7RRuc)qRH:RM0R#8D_kFOoH;R
RRRRRRBRWpRiR:MRHR8#0_FkDo;HORRRRRRRR
RRRRRRRRRW R:RRRRHM#_08koDFHRO
RRRRR;R2RCR
MO8RFFlbM0CM;F
OlMbFCRM0Xv)qn4cX7RRRb0FsRR5
RRRRR7RRuRmRRF:Rk#0R0k8_DHFoOR;RRRRRRRR
RRRRR1RRuRmRRF:Rk#0R0k8_DHFoO
;
RRRRRRRRqRjRRRR:H#MR0k8_DHFoOR;
RRRRRqRR4RRRRH:RM0R#8D_kFOoH;R
RRRRRR.RqRRRR:MRHR8#0_FkDo;HO
RRRRRRRRRqdR:RRRRHM#_08koDFH
O;RRRRRRRRqRcRRRR:H#MR0k8_DHFoOR;
RRRRRqRR6RRRRH:RM0R#8D_kFOoH;R
RRRRRRRR7RRRR:MRHR8#0_FkDo;HO
RRRRRRRR)7uq:jRRRHM#_08koDFH
O;RRRRRRRR7qu)4RR:H#MR0k8_DHFoOR;
RRRRR7RRu.)qRH:RM0R#8D_kFOoH;R
RRRRRRuR7)Rqd:MRHR8#0_FkDo;HO
RRRRRRRR)7uq:cRRRHM#_08koDFH
O;RRRRRRRR7qu)6RR:H#MR0k8_DHFoOR;
RRRRRWRRBRpiRH:RM0R#8D_kFOoH;RRRRRRRRR
RRRRRR RWRRRR:MRHR8#0_FkDo
HORRRRR2RR;
RRCRM8ObFlFMMC0V;
k0MOHRFMVOkM_HHM0R5L:FRLFNDCMs2RCs0kM0R#soHMR
H#LHCoMR
RH5VRL02RE
CMRRRRskC0s"M5"
2;RDRC#RC
RsRRCs0kMB5"F8kDR0MFRbHlDCClMA0RD	FORv)q3#RQRC0ERNsC88RN8#sC#CRso0H#C8sCRHk#M0oRE#CRNRlCOODF	#RNRC0ERv)q?;"2
CRRMH8RVC;
MV8Rk_MOH0MH;k
VMHO0FoMRCC0_M88_CEb05x#HCRR:HCM0oRCs;CR8bR0E:MRH0CCoss2RCs0kMMRH0CCos#RH
sPNHDNLCHRlMH_#x:CRR0HMCsoCRR:=jL;
CMoH
lRRH#M_HRxC:8=RCEb0;R
RH5VR#CHxR8<RCEb02ER0CRM
RlRRH#M_HRxC:#=RH;xC
CRRMH8RVR;
R0sCkRsMl_HM#CHx;M
C8CRo0M_C8C_8b;0E
0N0skHL0oCRCsMCNs0F_bsCFRs0:0R#soHM;0
N0LsHkR0CoCCMsFN0sC_sb0FsRRFVLODF	N_slRR:NEsOHO0C0CksRRH#VOkM_HHM0N5s8_8ss2Co;-
-RoLCHLMRD	FORlsNRbHlDCClM00NHRFM#MHoN
D#0C$bR0HM_sNsNH$R#sRNsRN$50jRF2R6RRFVHCM0o;Cs
MOF#M0N0HRI8_0ENNss$RR:H_M0NNss$=R:R,54RR.,cg,R,UR4,nRd2O;
F0M#NRM080CbEs_NsRN$:MRH0s_NsRN$:5=R4UndcU,R4,g.Rgcjn.,Rj,cUR.4jc6,R4;.2
MOF#M0N0HR8PRd.:MRH0CCos=R:RH5I8-0E4d2/nO;
F0M#NRM084HPnRR:HCM0oRCs:5=RI0H8E2-4/;4U
MOF#M0N0HR8P:URR0HMCsoCRR:=58IH04E-2;/g
MOF#M0N0HR8P:cRR0HMCsoCRR:=58IH04E-2;/c
MOF#M0N0HR8P:.RR0HMCsoCRR:=58IH04E-2;/.
MOF#M0N0HR8P:4RR0HMCsoCRR:=58IH04E-2;/4
F
OMN#0ML0RF4FDRL:RFCFDN:MR=8R5HRP4>2Rj;F
OMN#0ML0RF.FDRL:RFCFDN:MR=8R5HRP.>2Rj;F
OMN#0ML0RFcFDRL:RFCFDN:MR=8R5HRPc>2Rj;F
OMN#0ML0RFUFDRL:RFCFDN:MR=8R5HRPU>2Rj;F
OMN#0ML0RF4FDnRR:LDFFCRNM:5=R84HPnRR>j
2;O#FM00NMRFLFDRd.:FRLFNDCM=R:RH58PRd.>2Rj;O

F0M#NRM084HPncdURH:RMo0CC:sR=8R5CEb0-/424UndcO;
F0M#NRM08UHP4Rg.:MRH0CCos=R:RC58b-0E4U2/4;g.
MOF#M0N0HR8PgcjnRR:HCM0oRCs:5=R80CbE2-4/gcjnO;
F0M#NRM08.HPjRcU:MRH0CCos=R:RC58b-0E4.2/j;cU
MOF#M0N0HR8P.4jcRR:HCM0oRCs:5=R80CbE2-4/.4jcO;
F0M#NRM086HP4:.RR0HMCsoCRR:=5b8C04E-24/6.
;
O#FM00NMRFLFD.64RL:RFCFDN:MR=8R5H4P6.RR>j
2;O#FM00NMRFLFD.4jcRR:LDFFCRNM:5=R84HPjR.c>2Rj;F
OMN#0ML0RF.FDjRcU:FRLFNDCM=R:RH58Pc.jURR>j
2;O#FM00NMRFLFDgcjnRR:LDFFCRNM:5=R8cHPjRgn>2Rj;F
OMN#0ML0RFUFD4Rg.:FRLFNDCM=R:RH58PgU4.RR>j
2;O#FM00NMRFLFDd4nU:cRRFLFDMCNRR:=5P8H4UndcRR>j
2;
MOF#M0N0kR#lH_I8R0E:MRH0CCos=R:RmAmph q'#bF5FLFDR42+mRAmqp hF'b#F5LF2D.RA+Rm mpqbh'FL#5FcFD2RR+Apmm 'qhb5F#LDFFU+2RRmAmph q'#bF5FLFD24n;F
OMN#0M#0Rk8l_CEb0RH:RMo0CC:sR=RR6-AR5m mpqbh'FL#5F6FD4R.2+mRAmqp hF'b#F5LFjD4.Rc2+mRAmqp hF'b#F5LFjD.cRU2+mRAmqp hF'b#F5LFjDcgRn2+mRAmqp hF'b#F5LF4DUg2.2;O

F0M#NRM0IE_OFCHO_8IH0:ERR0HMCsoCRR:=I0H8Es_Ns5N$#_klI0H8E
2;O#FM00NMROI_EOFHCC_8bR0E:MRH0CCos=R:Rb8C0NE_s$sN5l#k_8IH0;E2
MOF#M0N0_R8OHEFOIC_HE80RH:RMo0CC:sR=HRI8_0ENNss$k5#lC_8b20E;F
OMN#0M80R_FOEH_OC80CbERR:HCM0oRCs:8=RCEb0_sNsN#$5k8l_CEb02
;
O#FM00NMRII_HE80_lMk_DOCD:#RR0HMCsoCRR:=58IH04E-2_/IOHEFOIC_HE80R4+R;F
OMN#0MI0R_b8C0ME_kOl_C#DDRH:RMo0CC:sR=8R5CEb0-/42IE_OFCHO_b8C0+ERR
4;
MOF#M0N0_R8I0H8Ek_MlC_ODRD#:MRH0CCos=R:RH5I8-0E482/_FOEH_OCI0H8ERR+4O;
F0M#NRM08C_8b_0EM_klODCD#RR:HCM0oRCs:5=R80CbE2-4/O8_EOFHCC_8bR0E+;R4
F
OMN#0MI0R_x#HCRR:HCM0oRCs:I=R_8IH0ME_kOl_C#DDRI*R_b8C0ME_kOl_C#DD;F
OMN#0M80R_x#HCRR:HCM0oRCs:8=R_8IH0ME_kOl_C#DDR8*R_b8C0ME_kOl_C#DD;O

F0M#NRM0LDFF_:8RRFLFDMCNRR:=5#8_HRxC-_RI#CHxRR<=j
2;O#FM00NMRFLFDR_I:FRLFNDCM=R:R0MF5FLFD2_8;O

F0M#NRM0OHEFOIC_HE80RH:RMo0CC:sR=AR5m mpqbh'FL#5F_FD8*2RRO8_EOFHCH_I820ER5+RApmm 'qhb5F#LDFF_RI2*_RIOHEFOIC_HE802O;
F0M#NRM0OHEFO8C_CEb0RH:RMo0CC:sR=AR5m mpqbh'FL#5F_FD8*2RRO8_EOFHCC_8b20ER5+RApmm 'qhb5F#LDFF_RI2*_RIOHEFO8C_CEb02O;
F0M#NRM0I0H8Ek_MlC_ODRD#:MRH0CCos=R:Rm5Amqp hF'b#F5LF8D_25R*I0H8E2-4/O8_EOFHCH_I820ER5+RApmm 'qhb5F#LDFF_RI2*IR5HE80-/42IE_OFCHO_8IH0RE2+;R4
MOF#M0N0CR8b_0EM_klODCD#RR:HCM0oRCs:5=RApmm 'qhb5F#LDFF_R82*C58b-0E482/_FOEH_OC80CbE+2RRm5Amqp hF'b#F5LFID_2RR*5b8C04E-2_/IOHEFO8C_CEb02RR+40;
$RbCF_k0L4k#_b0$C#RHRsNsN5$R80CbEk_MlC_OD-D#4FR8IFM0RRj,I0H8Ek_MlC_OD-D#4FR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNR0Fk_#Lk4RR:F_k0L4k#_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFR8s_FRk05bHMk00RFsR0H0-#N#0C2$
0bFCRkL0_k_#.0C$bRRH#NNss$8R5CEb0_lMk_DOCD4#-RI8FMR0Fj.,R*8IH0ME_kOl_C#DD+84RF0IMF2RjRRFV#_08DHFoO#;
HNoMDkRF0k_L#:.RR0Fk_#Lk.$_0bRC;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RV_Rs80FkRM5HbRk000FRs#H-0CN0#02
$RbCF_k0Lck#_b0$C#RHRsNsN5$R80CbEk_MlC_OD-D#4FR8IFM0RRj,cH*I8_0EM_klODCD#R+d8MFI0jFR2VRFR8#0_oDFH
O;#MHoNFDRkL0_kR#c:kRF0k_L#0c_$;bCRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$FsVR_k8F0HR5M0bkRR0F0-sH#00NC
#20C$bR0Fk_#LkU$_0bHCR#sRNsRN$5b8C0ME_kOl_C#DD-84RF0IMF,RjRIU*HE80_lMk_DOCD(#+RI8FMR0FjF2RV0R#8F_Do;HO
o#HMRNDF_k0LUk#RF:RkL0_k_#U0C$b;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFVsF_8k50RHkMb0FR0RH0s-N#002C#
b0$CNRbs$H0_#LkU$_0bHCR#sRNsRN$5b8C0ME_kOl_C#DD-84RF0IMF,RjR8IH0ME_kOl_C#DD-84RF0IMF2RjRRFV#_08DHFoO#;
HNoMDNRbs$H0_#LkURR:bHNs0L$_k_#U0C$b;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RV_Rs80FkRM5HbRk000FRs#H-0CN0#02
$RbCF_k0L4k#n$_0bHCR#sRNsRN$5b8C0ME_kOl_C#DD-84RF0IMF,RjR*4nI0H8Ek_MlC_OD+D#486RF0IMF2RjRRFV#_08DHFoO#;
HNoMDkRF0k_L#R4n:kRF0k_L#_4n0C$b;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RV_Rs80FkRM5HbRk000FRs#H-0CN0#02
$RbCbHNs0L$_kn#4_b0$C#RHRsNsN5$R80CbEk_MlC_OD-D#4FR8IFM0RRj,.H*I8_0EM_klODCD#R+48MFI0jFR2VRFR8#0_oDFH
O;#MHoNbDRN0sH$k_L#R4n:NRbs$H0_#Lk40n_$;bCRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$FsVR_k8F0HR5M0bkRR0F0-sH#00NC
#20C$bR0Fk_#Lkd0._$RbCHN#Rs$sNRC58b_0EM_klODCD#R-48MFI0jFR,.Rd*8IH0ME_kOl_C#DD+Rd48MFI0jFR2VRFR8#0_oDFH
O;#MHoNFDRkL0_k.#dRF:RkL0_k.#d_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$FsVR_k8F0HR5M0bkRR0F0-sH#00NC
#20C$bRsbNH_0$Ldk#.$_0bHCR#sRNsRN$5b8C0ME_kOl_C#DD-84RF0IMF,RjRIc*HE80_lMk_DOCDd#+RI8FMR0FjF2RV0R#8F_Do;HO
o#HMRNDbHNs0L$_k.#dRb:RN0sH$k_L#_d.0C$b;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFVsF_8k50RHkMb0FR0RH0s-N#002C#
o#HMRNDF_k0C:MRR8#0_oDFHPO_CFO0sC58b_0EM_klODCD#R-48MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-MRCNCLD#FRVssR0H0-#N#0C
o#HMRNDI_s0C:MRR8#0_oDFHPO_CFO0sC58b_0EM_klODCD#R-48MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-sRIHR0CCLMNDRC#VRFsCENORIsFRRFV)RqvODCD#H
#oDMNR_HMsRCo:0R#8F_Do_HOP0COFIs5HE80+Rd68MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--k8#CRR0FsHCo#s0CRh7QRH
#oDMNR0Fk_osCR#:R0D8_FOoH_OPC05FsI0H8E6+dRI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--k8#CRR0FsHCo#s0CRz7maH
#oDMNR0Fk_osC4RR:#_08DHFoOC_POs0F58IH04E-RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-k-R#RC80OFRE#FFCCRL0CICMQR7hMRN8kRF00bkRRFVAODF	qR)vH
#oDMNR8sN_osCR#:R0D8_FOoH_OPC05FsNs88I0H8ER-48MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--k8#CRR0FsHCo#s0CR7)q7#)
HNoMDNRI8C_soRR:#_08DHFoOC_POs0F58N8s8IH04E-RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RCk#8FR0RosCHC#0sqRW7
7)#MHoNDDRFsI_Ns88R#:R0D8_FOoH_OPC05Fs48dRF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-s-RNs88R0LH#MRHbRk00)FRqOvRC#DDRR5cL#H0RJsCkCHs8#2
HNoMDFRDIN_I8R8s:0R#8F_Do_HOP0COF4s5dFR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-NRI8R8sL#H0RbHMk00RFqR)vCRODRD#5LcRHR0#skCJH8sC2H
#oDMNR7)q70)_l:bRR8#0_oDFHPO_CFO0s85N8HsI8-0E4FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-#RkC08RFHRbbHCDM)CRq)77
o#HMRNDW7q7)l_0bRR:#_08DHFoOC_POs0F58N8s8IH04E-RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RCk#8FR0RbbHCMDHCqRW7
7)#MHoN7DRQ0h_l:bRR8#0_oDFHPO_CFO0sH5I8-0E4FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--k8#CRR0FbCHbDCHMRh7Q
o#HMRNDW0 _l:bRR8#0_oDFHRO;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RCk#8FR0RbbHCMDHC RW
R--CRM8LODF	NRsllRHblDCCNM00MHFRo#HM#ND
R--LHCoMCR#D0CORlsNRbHlDCClM00NHRFM#MHoN
D#VOkM0MHFR0oC_lMk_5nc80CbEH:RMo0CCRs2skC0sHMRMo0CCHsR#N
PsLHNDPCRN:DRR0HMCsoCRR:=jL;
CMoH
PRRN:DR=CR8b/0En
c;RVRHR855CEb0R8lFR2ncRc>RU02RE
CMRRRRPRND:P=RN+DRR
4;RMRC8VRH;R
RskC0sPMRN
D;CRM8o_C0M_kln
c;VOkM0MHFR0oC_VDC0CFPs._d5b8C0:ERR0HMCsoC2CRs0MksR0HMCsoCR
H#LHCoMR
RskC0s8M5CEb0R8lFR2nc;M
C8CRo0C_DVP0FCds_.V;
k0MOHRFMo_C0D0CVFsPC5b8C0:ERR0HMCsoC;NRlGRR:HCM0o2CsR0sCkRsMHCM0oRCsHP#
NNsHLRDCPRND:MRH0CCos=R:R
j;LHCoMR
RH5VR80CbERR-lRNG>j=R2ER0CRM
RPRRN:DR=CR8bR0E-NRlGR;
R#CDCR
RRNRPD=R:Rb8C0
E;RMRC8VRH;R
RskC0sPM5N;D2
8CMR0oC_VDC0CFPsV;
k0MOHRFMo_C0M_kld8.5CEb0RH:RMo0CCRs2skC0sHMRMo0CCHsR#N
PsLHNDPCRN:DRR0HMCsoCRR:=jL;
CMoH
HRRV8R5CEb0RR<=cNURM88RCEb0R4>Rn02RE
CMRRRRRDPNRR:=4R;
R8CMR;HV
sRRCs0kMNRPDC;
Mo8RCM0_kdl_.V;
k0MOHRFMo_C0M_kl48n5CEb0RH:RMo0CCRs2skC0sHMRMo0CCHsR#N
PsLHNDPCRN:DRR0HMCsoCRR:=jL;
CMoH
HRRV8R5CEb0RR<=4NnRM88RCEb0Rj>R2ER0CRM
RRRRPRND:4=R;R
RCRM8H
V;RCRs0MksRDPN;M
C8CRo0k_Mln_4;F
OMN#0MM0RkOl_C_DDn:cRR0HMCsoCRR:=o_C0M_kln8c5CEb02O;
F0M#NRM0D0CVFsPC_Rd.:MRH0CCos=R:R0oC_VDC0CFPs._d5b8C0;E2
MOF#M0N0kRMlC_ODdD_.RR:HCM0oRCs:o=RCM0_kdl_.C5DVP0FCds_.
2;O#FM00NMRVDC0CFPsn_4RH:RMo0CC:sR=CRo0C_DVP0FCDs5CFV0P_CsdR.,d;.2
MOF#M0N0kRMlC_OD4D_nRR:HCM0oRCs:o=RCM0_k4l_nC5DVP0FC4s_n
2;
b0$CkRF0k_L#$_0bnC_cH#R#sRNsRN$5lMk_DOCDc_nRI8FMR0FjI,RHE80-84RF0IMF2RjRRFV#_08DHFoO0;
$RbCF_k0L_k#0C$b_#d.RRH#NNss$MR5kOl_C_DDd8.RF0IMF,RjR8IH04E-RI8FMR0FjF2RV0R#8F_Do;HO
b0$CkRF0k_L#$_0b4C_nH#R#sRNsRN$5lMk_DOCDn_4RI8FMR0FjI,RHE80-84RF0IMF2RjRRFV#_08DHFoO#;
HNoMDkRF0k_L#c_n#RR:F_k0L_k#0C$b_#nc;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFV80FkRM5HbRk000FRs#H-0CN0##2
HNoMDkRF0k_L#._d#RR:F_k0L_k#0C$b_#d.;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFV80FkRM5HbRk000FRs#H-0CN0##2
HNoMDkRF0k_L#n_4#RR:F_k0L_k#0C$b_#4n;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFV80FkRM5HbRk000FRs#H-0CN0##2
HNoMDkRF0M_C_:#RR8#0_oDFHPO_CFO0sk5MlC_ODnD_cFR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--CLMNDRC#VRFs0-sH#00NC##
HNoMDkRF0M_C_Rd.:0R#8F_Do;HO
o#HMRNDF_k0C4M_nRR:#_08DHFoO#;
HNoMDsRI0M_C_:#RR8#0_oDFHPO_CFO0sk5MlC_ODnD_cFR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--I0sHCMRCNCLD#FRVsNRCOsERFFIRVqR)vCROD
D##MHoNIDRsC0_M._dR#:R0D8_FOoH;H
#oDMNR0Is__CM4:nRR8#0_oDFH
O;#MHoNHDRMC_soR_#:0R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-k-R#RC80sFRC#oH0RCs7RQh
o#HMRNDF_k0s_Co#RR:#_08DHFoOC_POs0F58IH04E-RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--k8#CRR0FsHCo#s0CRz7maH
#oDMNR8sN_osC_:#RR8#0_oDFHPO_CFO0s85N8HsI8-0E4FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-#RkC08RFCRso0H#CqsR7
7)#MHoNIDRNs8_C#o_R#:R0D8_FOoH_OPC05FsNs88I0H8ER-48MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--k8#CRR0FsHCo#s0CR7q7)H
#oDMNRIDF_8sN8#s_R#:R0D8_FOoH_OPC05Fs6FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-8RN8LsRHR0#HkMb0FR0Rv)qRDOCD5#RcHRL0s#RCHJks2C8
o#HMRNDD_FII8N8sR_#:0R#8F_Do_HOP0COF6s5RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-R8N8sHRL0H#RM0bkRR0F)RqvODCD#cR5R0LH#CRsJskHC
82-C-RM#8RCODC0NRsllRHblDCCNM00MHFRo#HM#ND
0N0skHL0\CR3lsN_VFV#\C0R#:R0MsHo
;
LHCoMR
Rz:cdRRHV58sN8ss_CRo2oCCMsCN0RR--oCCMsCN0RFLDOs	RNRl
R-RR-VRQR8N8s8IH0<ERRFOEH_OCI0H8E#RN#MHoR''jRR0Fk#MkCL8RH
0#RRRRzRjR:VRHR85N8HsI8R0E=2R4RMoCC0sNCR
SRDRRFsI_Ns88RR<="jjjjjjjjjjjjRj"&NRs8C_so25j;R
SRDRRFII_Ns88RR<="jjjjjjjjjjjjRj"&NRI8C_so25j;C
SMo8RCsMCNR0Cz
j;RRRRzR4R:VRHR85N8HsI8R0E=2R.RMoCC0sNCS
SD_FIs8N8s=R<Rj"jjjjjjjjjjRj"&NRs8C_soR548MFI0jFR2S;
RRRRD_FII8N8s=R<Rj"jjjjjjjjjjRj"&NRI8C_soR548MFI0jFR2S;
CRM8oCCMsCN0R;z4
RRRRRz.RH:RVNR58I8sHE80Rd=R2CRoMNCs0SC
SIDF_8sN8<sR=jR"jjjjjjjjjRj"&NRs8C_soR5.8MFI0jFR2S;
RRRRD_FII8N8s=R<Rj"jjjjjjjjjj&"RR8IN_osC58.RF0IMF2Rj;C
SMo8RCsMCNR0Cz
.;RRRRzRdR:VRHR85N8HsI8R0E=2RcRMoCC0sNCS
SD_FIs8N8s=R<Rj"jjjjjjjjj"RR&s_N8s5CodFR8IFM0R;j2
RSRRFRDIN_I8R8s<"=RjjjjjjjjjRj"&NRI8C_soR5d8MFI0jFR2S;
CRM8oCCMsCN0R;zd
RRRRRzcRH:RVNR58I8sHE80R6=R2CRoMNCs0SC
RRRRD_FIs8N8s=R<Rj"jjjjjj"jjRs&RNs8_Cco5RI8FMR0Fj
2;SRRRRIDF_8IN8<sR=jR"jjjjjjjj"RR&I_N8s5CocFR8IFM0R;j2
MSC8CRoMNCs0zCRcR;
RzRR6:RRRRHV58N8s8IH0=ERRRn2oCCMsCN0
RSRRFRDIN_s8R8s<"=Rjjjjjjjj"RR&s_N8s5Co6FR8IFM0R;j2
DSSFII_Ns88RR<="jjjjjjjj&"RR8IN_osC586RF0IMF2Rj;C
SMo8RCsMCNR0Cz
6;RRRRzRnR:VRHR85N8HsI8R0E=2R(RMoCC0sNCR
SRDRRFsI_Ns88RR<="jjjjjjj"RR&s_N8s5ConFR8IFM0R;j2
DSSFII_Ns88RR<="jjjjjjj"RR&I_N8s5ConFR8IFM0R;j2
MSC8CRoMNCs0zCRnR;
RzRR(:RRRRHV58N8s8IH0=ERRRU2oCCMsCN0
RSRRFRDIN_s8R8s<"=RjjjjjRj"&NRs8C_soR5(8MFI0jFR2S;
SIDF_8IN8<sR=jR"jjjjj&"RR8IN_osC58(RF0IMF2Rj;C
SMo8RCsMCNR0Cz
(;RRRRzRUR:VRHR85N8HsI8R0E=2RgRMoCC0sNCR
SRDRRFsI_Ns88RR<="jjjjRj"&NRs8C_soR5U8MFI0jFR2S;
SIDF_8IN8<sR=jR"jjjj"RR&I_N8s5CoUFR8IFM0R;j2
MSC8CRoMNCs0zCRUR;
RzRRg:RRRRHV58N8s8IH0=ERR24jRMoCC0sNCR
SRDRRFsI_Ns88RR<="jjjj&"RR8sN_osC58gRF0IMF2Rj;S
SD_FII8N8s=R<Rj"jjRj"&NRI8C_soR5g8MFI0jFR2S;
CRM8oCCMsCN0R;zg
RRRRjz4RRR:H5VRNs88I0H8ERR=4R42oCCMsCN0
RSRRFRDIN_s8R8s<"=Rj"jjRs&RNs8_C4o5jFR8IFM0R;j2
DSSFII_Ns88RR<="jjj"RR&I_N8s5Co48jRF0IMF2Rj;C
SMo8RCsMCNR0Cz;4j
RRRR4z4RRR:H5VRNs88I0H8ERR=4R.2oCCMsCN0
RSRRFRDIN_s8R8s<"=RjRj"&NRs8C_so454RI8FMR0Fj
2;SFSDIN_I8R8s<"=RjRj"&NRI8C_so454RI8FMR0Fj
2;S8CMRMoCC0sNC4Rz4R;
RzRR4R.R:VRHR85N8HsI8R0E=dR42CRoMNCs0SC
RRRRD_FIs8N8s=R<R''jRs&RNs8_C4o5.FR8IFM0R;j2
DSSFII_Ns88RR<='Rj'&NRI8C_so.54RI8FMR0Fj
2;S8CMRMoCC0sNC4Rz.R;
RzRR4RdR:VRHR85N8HsI8R0E>dR42CRoMNCs0SC
RRRRD_FIs8N8s=R<R8sN_osC5R4d8MFI0jFR2S;
RRRRD_FII8N8s=R<R8IN_osC5R4d8MFI0jFR2S;
CRM8oCCMsCN0Rdz4;R

R-RR-VRQRH58MC_sos2RC#oH0RCs7RQhkM#HopRBiR
RR4Rzc:RRRRHV5M8H_osC2CRoMNCs0RC
RRRRRbRRsCFO#5#RB,piRh7Q2CRLo
HMRRRRRRRRRRRRH5VRBRpi=4R''MRN8pRBiP'CC2M0RC0EMR
RRRRRRRRRRRRRRMRH_osCRR<=5j"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjRj"&QR7h
2;RRRRRRRRRRRRCRM8H
V;RRRRRRRRCRM8bOsFC;##
MSC8CRoMNCs0zCR4
c;RRRRzR46RH:RVMR5F80RHsM_CRo2oCCMsCN0
RRRRRRRRRRRR_HMsRCo<5=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj&"RRh7Q2S;
CRM8oCCMsCN0R6z4;R

R-RR-VRQR85sF_k0s2CoRosCHC#0s_R)7amzRHk#M)oR_pmBiR
RR4Rzn:RRRRHV5k8F0C_soo2RCsMCN
0CRRRRRRRRbOsFCR##5pmBiF,Rks0_C2o4RoLCHRM
RRRRRRRRRHRRVmR5BRpi=4R''MRN8BRmpCi'P0CM2ER0CRM
RRRRRRRRRRRRR7RRmRza<F=Rks0_C;o4
RRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMRFbsO#C#;R
RRRRRRMRC8CRoMNCs0zCR4
n;RRRRzR4(RH:RVMR5F80RF_k0s2CoRMoCC0sNCR
RRRRRRRRRRmR7z<aR=kRF0C_so
4;S8CMRMoCC0sNC4Rz(
;
RRRR-Q-RVsR5Ns88_osC2CRso0H#C)sRq)77RHk#MmoRB
piRRRRzs4nRRR:H5VRs8N8sC_soo2RCsMCN
0C-R-RRRRRRsRbF#OC#mR5B,piR7)q7R)2LHCoM-
-RRRRRRRRRRRRH5VRmiBpR'=R4N'RMm8RB'piCMPC002RE
CM-R-RRRRRRRRRRRRRRNRs8C_so=R<R7)q7N)58I8sHE80-84RF0IMF2Rj;-
-RRRRRRRRRRRRCRM8H
V;-R-RRRRRRMRC8sRbF#OC#-;
-MSC8CRoMNCs0zCR4;ns
R--RzRR4R(s:VRHRF5M0NRs8_8ss2CoRMoCC0sNCR
RRRRRRRRRRNRs8C_so=R<R7)q7
);S8CMRMoCC0sNC4Rzn
s;
-S-RRQV58IN8ss_CRo2sHCo#s0CR7Wq7k)R#oHMRmW_B
piRRRRzI4nRRR:H5VRI8N8sC_soo2RCsMCN
0CRRRRRRRRbOsFCR##5iBp,qRW727)RoLCHRM
RRRRRRRRRHRRVBR5p=iRR''4R8NMRiBp'CCPMR020MEC
RRRRRRRRRRRRRRRR8IN_osCRR<=W7q7)85N8HsI8-0E4FR8IFM0R;j2
RRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMRFbsO#C#;C
SMo8RCsMCNR0CzI4n;R
RR4Rz(:IRRRHV50MFR8IN8ss_CRo2oCCMsCN0
RRRRRRRRRRRR8IN_osCRR<=W7q7)S;
CRM8oCCMsCN0R(z4I
;
RRRR- -RGN0sRoDFHVORF7sRkRNDb0FsR#ONCz
SsRCo:sRbF#OC#p5BiL2RCMoH
RSRH5VRB'pi he aMRN8pRBiRR='24'RC0EMR
SRQR7hl_0b=R<Rh7Q;R
SRqR)7_7)0Rlb<)=Rq)77;R
SRqRW7_7)0Rlb<W=Rq)77;R
SR RW_b0lRR<=W
 ;SCRRMH8RVS;
CRM8bOsFC;##
-
S-VRQRN)C88Rq8#sC#RR=W0sHC8Rq8#sC#L,R$#bN#QR7hFR0R0FkbRk0HWVR #RHRNCML8DC
lSzk:GRRFbsO#C#5_W 0,lbR7)q70)_lRb,W7q7)l_0b7,RQ0h_lRb,F_k0s2Co
RSRLHCoMR
SRHRRVWR5q)77_b0lR)=Rq)77_b0lR8NMR_W 0Rlb=4R''02RE
CMSRSRF_k0s4CoRR<=7_Qh0;lb
CSSD
#CSRSRF_k0s4CoRR<=F_k0s5CoI0H8ER-48MFI0jFR2S;
S8CMR;HV
MSC8sRbF#OC#S;
RRRR
RRRRR--tCCMsCN0RC0ERv)qRDOCDN#RM#8RCODC0FRDoRHOVRFs)Aqv41n_44_1
4SzURR:H5VROHEFOIC_HE80R4=R2CRoMNCs0RC
RSRRzR4g:FRVsRRHH5MR80CbEk_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0SC
-Q-RVNR58I8sHE80R4>RcM2RCRC80OFRs0CNCsRIHR0CCLMNDNCRMF8Rkk0b0MRCNCLDRD#CCRO0DHFoOR
RRRRRRzRS.:jRRRHV58N8s8IH0>ERR24cRMoCC0sNC-
S-HRVGFRVsNROD4DRd(UU,CR#D0CORRFV0#sH0CN0R0MFRHLCMsoRC#oH0CCs8S
SSkSF0M_C5RH2<'=R4I'RERCM57)q70)_lNb58I8sHE80-84RF0IMFcR42RR=HC2RDR#C';j'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RWRCIEMIR5Ns8_CNo58I8sHE80-84RF0IMFcR42RR=HC2RDR#C';j'
RRRRRRRRMSC8CRoMNCs0zCR.
j;SR--Q5VRNs88I0H8E=R<R24cRRMFI0sHCMRCNCLDRRFsFbk0kC0RMDNLCCR#D0CORoDFHMORCCC88S
RRRRRS4z.RH:RVNR58I8sHE80RR<=4Rc2oCCMsCN0
SSSS0Fk_5CMH<2R=4R''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=W
 ;RRRRRRRRS8CMRMoCC0sNC.Rz4S;
-t-RCsMCNR0C0REC)RqvODCD#MRN8sR0H0-#N#0C
RRRRRRRR.Sz.RR:VRFs[MRHRH5I8_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
RRRRRRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVAv)q_d4nU4cX7RR:DCNLD#RHR""W;R
RRRRRRRRRRRRRRCRLo
HMRRRRRRRRRRRRSqA)vn_4dXUc4:7RRv)qA_4n114_4R
SRRRRRRRRRbRRFRs0lRNb5q7Q5Rj2=H>RMC_so25[,7Rq7R)q=D>RFII_Ns885R4d8MFI0jFR27,RQ=AR>jR""q,R7A7)RR=>D_FIs8N8sd54RI8FMR0Fj
2,SSSS Rhq='>R4R',1q1)RR=>',j'RqW RR=>I_s0CHM52B,RpRiq=B>RpRi, RhA='>R4R',1A1)RR=>',j'RAW RR=>',j'RiBpA>R=RiBp,S
SSRRRRq7mRR=>FMbC,mR7A25jRR=>F_k0L4k#5[H,2
2;
RRRRRRRRRRRRRRRR0Fk_osC5R[2<F=RkL0_k5#4H2,[RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRCRSMo8RCsMCNR0Cz;..
RRRRCRSMo8RCsMCNR0Cz;4g
RRRR8CMRMoCC0sNC4RzUR;RRRR
RRRRRR
RR-R-RMtCC0sNCER0CqR)vCRODRD#NRM8#CCDOD0RFOoHRsVFRv)qA_4n11._.z
S.:dRRRHV5FOEH_OCI0H8ERR=.o2RCsMCN
0CRRRRScz.RV:RFHsRRRHM5b8C0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CSR--Q5VRNs88I0H8ERR>4Rd2M8CCRR0FONsC0ICRsCH0RNCMLRDCNRM8Fbk0kC0RMDNLCCR#D0CORoDFHRO
RRRRRSRRzR.6:VRHR85N8HsI8R0E>dR42CRoMNCs0SC
-V-RHVGRFOsRNRDD4UdU(#,RCODC0VRFRH0s#00NCFRM0CRLHRMosHCo#s0CCR8
RRRRRRRRRRRRRFRRkC0_M25HRR<='R4'IMECRq5)7_7)05lbNs88I0H8ER-48MFI04FRd=2RRRH2CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R ERIC5MRI_N8s5CoNs88I0H8ER-48MFI04FRd=2RRRH2CCD#R''j;R
RRRRRRCRSMo8RCsMCNR0Cz;.6
-S-RRQV58N8s8IH0<ER=dR42FRMRHIs0CCRMDNLCsRFR0FkbRk0CLMND#CRCODC0FRDoRHOM8CCCR8
SRRRR.SznRR:H5VRNs88I0H8E=R<R24dRMoCC0sNCR
SRRRRRRRRRFRRkC0_M25HRR<=';4'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RW;R
RRRRRRCRSMo8RCsMCNR0Cz;.n
-S-RMtCC0sNCER0CqR)vCRODRD#NRM80-sH#00NCR#
RRRRRSRRzR.(:FRVsRR[H5MRI0H8Ek_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0RC
RRRRRRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)RAqUv_4Xg..:7RRLDNCHDR#WR""R;
RRRRRRRRRRRRRLRRCMoH
RRRRRRRRRRRR)SAqUv_4Xg..:7RRv)qA_4n11._.R
SRRRRRRRRRbRRFRs0lRNb5q7QRR=>HsM_C.o5*4[+RI8FMR0F.2*[,7Rq7R)q=D>RFII_Ns885R4.8MFI0jFR27,RQ=AR>jR"jR",q)77A>R=RIDF_8sN84s5.FR8IFM0R,j2
SSSRRRR Rhq='>R4R',1q1)RR=>',j'RqW RR=>I_s0CHM52B,RpRiq=B>RpRi, RhA='>R4R',1A1)RR=>',j'RAW RR=>',j'RiBpA>R=RiBp,S
SSRRRRq7mRR=>FMbC,mR7A254RR=>F_k0L.k#5.H,*4[+27,RmjA52>R=R0Fk_#Lk.,5HR[.*2
2;RRRRRRRRRRRRRRRRF_k0s5Co.2*[RR<=F_k0L.k#5.H,*R[2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5[.*+R42<F=RkL0_k5#.H*,.[2+4RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRCRSMo8RCsMCNR0Cz;.(
RRRRCRSMo8RCsMCNR0Cz;.c
RRRR8CMRMoCC0sNC.RzdR;R
R
SR-RR-CRtMNCs00CRE)CRqOvRC#DDR8NMRD#CCRO0DHFoOFRVsqR)vnA4__1c1Sc
zR.U:VRHRE5OFCHO_8IH0=ERRRc2oCCMsCN0
RRRR.SzgRR:VRFsHMRHRC58b_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
-S-RRQV58N8s8IH0>ERR24.RCMC8FR0RCOsNR0CI0sHCMRCNCLDR8NMR0FkbRk0CLMND#CRCODC0FRDo
HORRRRRRRRSjzdRH:RVNR58I8sHE80R4>R.o2RCsMCN
0CSR--VRHGVRFsODNDRU4dUR(,#CCDOF0RVsR0HN#00MCRFL0RCoHMRosCHC#0s
C8RRRRRRRRRRRRRRRRF_k0CHM52=R<R''4RCIEM)R5q)77_b0l58N8s8IH04E-RI8FMR0F4R.2=2RHR#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=WI RERCM58IN_osC58N8s8IH04E-RI8FMR0F4R.2=2RHR#CDCjR''R;
RRRRRSRRCRM8oCCMsCN0Rjzd;-
S-VRQR85N8HsI8R0E<4=R.M2RFsRIHR0CCLMNDFCRskRF00bkRNCMLRDC#CCDOD0RFOoHRCMC8
C8RRSRRzRSd:4RRRHV58N8s8IH0<ER=.R42CRoMNCs0SC
SFSSkC0_M25HRR<=';4'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RW;R
RRRRRRCRSMo8RCsMCNR0Cz;d4
-S-RMtCC0sNCER0CqR)vCRODRD#NRM80-sH#00NCR#
RRRRRSRRzRd.:FRVsRR[H5MRI0H8Ek_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0RC
RRRRRRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)RAqcv_jXgnc:7RRLDNCHDR#WR""R;
RRRRRRRRRRRRRLRRCMoH
RRRRRRRRRRRR)SAqcv_jXgnc:7RRv)qA_4n11c_cR
SRRRRRRRRRbRRFRs0lRNb5q7QRR=>HsM_Cco5*d[+RI8FMR0Fc2*[,7Rq7R)q=D>RFII_Ns885R448MFI0jFR27,RQ=AR>jR"j"jj,7Rq7R)A=D>RFsI_Ns885R448MFI0jFR2S,
S SSh=qR>4R''1,R1R)q='>RjR',WR q=I>RsC0_M25H,pRBi=qR>pRBi ,Rh=AR>4R''1,R1R)A='>RjR',WR A='>RjR',BApiRR=>B,pi
SSSSq7mRR=>FMbC,mR7A25dRR=>F_k0Lck#5RH,c+*[dR2,75mA.=2R>kRF0k_L#Hc5,[c*+,.2RS
SSmS7A254RR=>F_k0Lck#5cH,*4[+27,RmjA52>R=R0Fk_#Lkc,5HR[c*2
2;RRRRRRRRRRRRRRRRF_k0s5Coc2*[RR<=F_k0Lck#5cH,*R[2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5[c*+R42<F=RkL0_k5#cH*,c[2+4RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so*5c[2+.RR<=F_k0Lck#5cH,*.[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cco5*d[+2=R<R0Fk_#Lkc,5Hc+*[dI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';
RRRRRRRRMSC8CRoMNCs0zCRd
.;RRRRRMSC8CRoMNCs0zCR.
g;RRRRCRM8oCCMsCN0RUz.;S

RRRR-t-RCsMCNR0C0REC)RqvODCD#MRN8CR#D0CORoDFHVORF)sRq4vAng_1_
1gSdzdRH:RVOR5EOFHCH_I8R0E=2RgRMoCC0sNCR
RRzRSd:cRRsVFRHHRM8R5CEb0_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNC-
S-VRQR85N8HsI8R0E>4R42CRMC08RFsROCCN0RHIs0CCRMDNLCMRN8kRF00bkRNCMLRDC#CCDOD0RFOoH
RRRRRRRRdSz6RR:H5VRNs88I0H8ERR>4R42oCCMsCN0
-S-RGVHRsVFRDONDdR4U,U(RD#CCRO0F0VRs0H#NR0CMRF0LMCHoCRso0H#C8sC
RRRRRRRRRRRRRRRR0Fk_5CMH<2R=4R''ERIC5MR)7q7)l_0b85N8HsI8-0E4FR8IFM0R244RH=R2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0CHM52=R<RRW IMECRN5I8C_so85N8HsI8-0E4FR8IFM0R244RH=R2DRC#'CRj
';RRRRRRRRS8CMRMoCC0sNCdRz6S;
-Q-RVNR58I8sHE80RR<=4R42MIFRsCH0RNCMLRDCFFsRkk0b0MRCNCLDRD#CCRO0DHFoOCRMC88C
RRSRSRRzRdn:VRHR85N8HsI8R0E<4=R4o2RCsMCN
0CSRRRRRRRRRRRR0Fk_5CMH<2R=4R''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=W
 ;RRRRRRRRS8CMRMoCC0sNCdRznS;
-t-RCsMCNR0C0REC)RqvODCD#MRN8sR0H0-#N#0C
RRRRRRRRdSz(RR:VRFs[MRHRH5I8_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
RRRRRRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVAv)q_c.jU7XURD:RNDLCRRH#";W"
RRRRRRRRRRRRRRRRoLCHRM
RRRRRRRRRSRRAv)q_c.jU7XUR):Rq4vAng_1_
1gRRRRRRRRRRRRRRRRRFRbsl0RN5bR7RQq=H>RMC_so*5g[R+(8MFI0gFR*,[2R7q7)=qR>FRDIN_I858s48jRF0IMF2Rj,QR7A>R=Rj"jjjjjj,j"R7q7)=AR>FRDIN_s858s48jRF0IMF2Rj,R
RRRRRRRRRRRRRRRRRRRRRRRRRRhR q>R=R''4,1R1)=qR>jR''W,R =qR>sRI0M_C5,H2RiBpq>R=RiBp,hR A>R=R''4,1R1)=AR>jR''W,R =AR>jR''B,RpRiA=B>RpRi,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRq7mRR=>FMbC,mR7A25(RR=>F_k0LUk#5UH,*([+27,RmnA52>R=R0Fk_#LkU,5HU+*[nR2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRA7m5R62=F>RkL0_k5#UH*,U[2+6,mR7A25cRR=>F_k0LUk#5UH,*c[+27,RmdA52>R=R0Fk_#LkU,5HU+*[dR2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRA7m5R.2=F>RkL0_k5#UH*,U[2+.,mR7A254RR=>F_k0LUk#5UH,*4[+27,RmjA52>R=R0Fk_#LkU,5HU2*[,RR
RRRRRRRRRRRRRRRRRRRRRRRRR7RRQ5uqj=2R>MRH_osC5[g*+,U2Ru7QA>R=R""j,mR7u=qR>bRFCRM,7Amu5Rj2=b>RN0sH$k_L#HU5,2[2;R
RRRRRRRRRRRRRRkRF0C_so*5g[<2R=kRF0k_L#HU5,[U*2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cgo5*4[+2=R<R0Fk_#LkU,5HU+*[4I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cog+*[.<2R=kRF0k_L#HU5,[U*+R.2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5[g*+Rd2<F=RkL0_k5#UH*,U[2+dRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so*5g[2+cRR<=F_k0LUk#5UH,*c[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cgo5*6[+2=R<R0Fk_#LkU,5HU+*[6I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cog+*[n<2R=kRF0k_L#HU5,[U*+Rn2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5[g*+R(2<F=RkL0_k5#UH*,U[2+(RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so*5g[2+URR<=bHNs0L$_k5#UH2,[RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRCRSMo8RCsMCNR0Cz;d(
RRRRCRSMo8RCsMCNR0Cz;dc
RRRR8CMRMoCC0sNCdRzd
;
SRRRRR--tCCMsCN0RC0ERv)qRDOCDN#RM#8RCODC0FRDoRHOVRFs)Aqv41n_41U_4SU
zRdU:VRHRE5OFCHO_8IH0=ERR24URMoCC0sNCR
RRzRSd:gRRsVFRHHRM8R5CEb0_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNC-
S-VRQR85N8HsI8R0E>jR42CRMC08RFsROCCN0RHIs0CCRMDNLCMRN8kRF00bkRNCMLRDC#CCDOD0RFOoH
RRRRRRRRcSzjRR:H5VRNs88I0H8ERR>4Rj2oCCMsCN0
-S-RGVHRsVFRDONDdR4U,U(RD#CCRO0F0VRs0H#NR0CMRF0LMCHoCRso0H#C8sC
RRRRRRRRRRRRRRRR0Fk_5CMH<2R=4R''ERIC5MR)7q7)l_0b85N8HsI8-0E4FR8IFM0R24jRH=R2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0CHM52=R<RRW IMECRN5I8C_so85N8HsI8-0E4FR8IFM0R24jRH=R2DRC#'CRj
';RRRRRRRRS8CMRMoCC0sNCcRzjS;
-Q-RVNR58I8sHE80RR<=4Rj2MIFRsCH0RNCMLRDCFFsRkk0b0MRCNCLDRD#CCRO0DHFoOCRMC88C
RRSRSRRzRc4:VRHR85N8HsI8R0E<4=Rjo2RCsMCN
0CSRRRRRRRRRRRR0Fk_5CMH<2R=4R''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=W
 ;RRRRRRRRS8CMRMoCC0sNCcRz4S;
-t-RCsMCNR0C0REC)RqvODCD#MRN8sR0H0-#N#0C
RRRRRRRRcSz.RR:VRFs[MRHRH5I8_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
RRRRRRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVAv)q_.4jcnX47RR:DCNLD#RHR""W;R
RRRRRRRRRRRRRRCRLo
HMRRRRRRRRRRRRSqA)vj_4.4cXn:7RRv)qA_4n1_4U1
4URRRRRRRRRRRRRRRRRFRbsl0RN5bR7RQq=H>RMC_soU54*4[+6FR8IFM0R*4U[R2,q)77q>R=RIDF_8IN8gs5RI8FMR0FjR2,7RQA=">Rjjjjjjjjjjjjjjjj"q,R7A7)RR=>D_FIs8N8sR5g8MFI0jFR2R,
RRRRRRRRRRRRRRRRRRRRRRRRR RRh=qR>4R''1,R1R)q='>RjR',WR q=I>RsC0_M25H,pRBi=qR>pRBi ,Rh=AR>4R''1,R1R)A='>RjR',WR A='>RjR',BApiRR=>B,piRR
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7q>R=RCFbM7,Rm4A56=2R>kRF0k_L#54nHn,4*4[+6R2,75mA4Rc2=F>RkL0_kn#454H,n+*[4,c2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7Ad542>R=R0Fk_#Lk4Hn5,*4n[d+427,Rm4A5.=2R>kRF0k_L#54nHn,4*4[+.R2,75mA4R42=F>RkL0_kn#454H,n+*[4,42RR
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7Aj542>R=R0Fk_#Lk4Hn5,*4n[j+427,RmgA52>R=R0Fk_#Lk4Hn5,*4n[2+g,mR7A25URR=>F_k0L4k#n,5H4[n*+,U2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7A25(RR=>F_k0L4k#n,5H4[n*+,(2RA7m5Rn2=F>RkL0_kn#454H,n+*[nR2,75mA6=2R>kRF0k_L#54nHn,4*6[+2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mAc=2R>kRF0k_L#54nHn,4*c[+27,RmdA52>R=R0Fk_#Lk4Hn5,*4n[2+d,mR7A25.RR=>F_k0L4k#n,5H4[n*+,.2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7A254RR=>F_k0L4k#n,5H4[n*+,42RA7m5Rj2=F>RkL0_kn#454H,n2*[,RR
RRRRRRRRRRRRRRRRRRRRRRRRR7RRQRuq=H>RMC_soU54*4[+(FR8IFM0R*4U[n+427,RQRuA=">Rj,j"Ru7mq>R=RCFbMR,
RRRRRRRRRRRRRRRRRRRRRRRRR7RRm5uA4=2R>NRbs$H0_#Lk4Hn5,[.*+,42Ru7mA25jRR=>bHNs0L$_kn#45.H,*2[2;R
RRRRRRRRRRRRRRkRF0C_soU54*R[2<F=RkL0_kn#454H,n2*[RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*4[+2=R<R0Fk_#Lk4Hn5,*4n[2+4RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*.[+2=R<R0Fk_#Lk4Hn5,*4n[2+.RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*d[+2=R<R0Fk_#Lk4Hn5,*4n[2+dRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*c[+2=R<R0Fk_#Lk4Hn5,*4n[2+cRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*6[+2=R<R0Fk_#Lk4Hn5,*4n[2+6RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*n[+2=R<R0Fk_#Lk4Hn5,*4n[2+nRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*([+2=R<R0Fk_#Lk4Hn5,*4n[2+(RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*U[+2=R<R0Fk_#Lk4Hn5,*4n[2+URCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*g[+2=R<R0Fk_#Lk4Hn5,*4n[2+gRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*4[+j<2R=kRF0k_L#54nHn,4*4[+jI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+244RR<=F_k0L4k#n,5H4[n*+244RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*4[+.<2R=kRF0k_L#54nHn,4*4[+.I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+24dRR<=F_k0L4k#n,5H4[n*+24dRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*4[+c<2R=kRF0k_L#54nHn,4*4[+cI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+246RR<=F_k0L4k#n,5H4[n*+246RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*4[+n<2R=NRbs$H0_#Lk4Hn5,[.*2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[4R(2<b=RN0sH$k_L#54nH*,.[2+4RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRCRSMo8RCsMCNR0Cz;c.
RRRRCRSMo8RCsMCNR0Cz;dg
RRRR8CMRMoCC0sNCdRzU
;
SRRRRR--tCCMsCN0RC0ERv)qRDOCDN#RM#8RCODC0FRDoRHOVRFs)Aqv41n_d1n_dSn
zNdURH:RVOR5EOFHCH_I8R0E=nRd2CRoMNCs0SC
RRRRzNdgRV:RFHsRRRHM5b8C0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CSR--Q5VRNs88I0H8ERR>gM2RCRC80OFRs0CNCsRIHR0CCLMNDNCRMF8Rkk0b0MRCNCLDRD#CCRO0DHFoOS
SSjzcNRR:H5VRNs88I0H8ERR>go2RCsMCN
0CSR--VRHGVRFsODNDRU4dUR(,#CCDOF0RVsR0HN#00MCRFL0RCoHMRosCHC#0s
C8SSSSF_k0CHM52=R<R''4RCIEM)R5q)77_b0l58N8s8IH04E-RI8FMR0Fg=2RRRH2CCD#R''j;S
SSsSI0M_C5RH2<W=R ERIC5MRI_N8s5CoNs88I0H8ER-48MFI0gFR2RR=HC2RDR#C';j'
SSSCRM8oCCMsCN0RjzcNS;
-Q-RVNR58I8sHE80RR<=gM2RFsRIHR0CCLMNDFCRskRF00bkRNCMLRDC#CCDOD0RFOoHRCMC8
C8SzSScR4N:VRHR85N8HsI8R0E<g=R2CRoMNCs0SC
SFSSkC0_M25HRR<=';4'
SSSS0Is_5CMH<2R= RW;S
SS8CMRMoCC0sNCcRz4
N;SR--tCCMsCN0RC0ERv)qRDOCDN#RM08Rs#H-0CN0#S
SS.zcNRR:VRFs[MRHRH5I8_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
RRRRRRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVAv)q_.64X7d.RD:RNDLCRRH#";W"
RRRRRRRRRRRRRRRRoLCHSM
SASS)_qv6X4.dR.7:qR)vnA4_n1d_n1d
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRbRRFRs0lRNb5q7QRR=>HsM_Cdo5n+*[d84RF0IMFnRd*,[2R7q7)=qR>FRDIN_I858sUFR8IFM0R,j2RA7QRR=>"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjR",q)77A>R=RIDF_8sN8Us5RI8FMR0Fj
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR Rhq='>R4R',1q1)RR=>',j'RqW RR=>I_s0CHM52B,RpRiq=B>RpRi, RhA='>R4R',1A1)RR=>',j'RAW RR=>',j'RiBpA>R=RiBp,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7q>R=RCFbM7,RmdA54=2R>kRF0k_L#5d.H.,d*d[+4R2,75mAdRj2=F>RkL0_k.#d5dH,.+*[d,j2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRA7m52.gRR=>F_k0Ldk#.,5Hd[.*+2.g,mR7AU5.2>R=R0Fk_#LkdH.5,*d.[U+.27,Rm.A5(=2R>kRF0k_L#5d.H.,d*.[+(
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mA.Rn2=F>RkL0_k.#d5dH,.+*[.,n2RA7m52.6RR=>F_k0Ldk#.,5Hd[.*+2.6,mR7Ac5.2>R=R0Fk_#LkdH.5,*d.[c+.2R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRm.A5d=2R>kRF0k_L#5d.H.,d*.[+dR2,75mA.R.2=F>RkL0_k.#d5dH,.+*[.,.2RA7m52.4RR=>F_k0Ldk#.,5Hd[.*+2.4,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7Aj5.2>R=R0Fk_#LkdH.5,*d.[j+.27,Rm4A5g=2R>kRF0k_L#5d.H.,d*4[+gR2,75mA4RU2=F>RkL0_k.#d5dH,.+*[4,U2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRA7m524(RR=>F_k0Ldk#.,5Hd[.*+24(,mR7An542>R=R0Fk_#LkdH.5,*d.[n+427,Rm4A56=2R>kRF0k_L#5d.H.,d*4[+6
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mA4Rc2=F>RkL0_k.#d5dH,.+*[4,c2RA7m524dRR=>F_k0Ldk#.,5Hd[.*+24d,mR7A.542>R=R0Fk_#LkdH.5,*d.[.+42R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRm4A54=2R>kRF0k_L#5d.H.,d*4[+4R2,75mA4Rj2=F>RkL0_k.#d5dH,.+*[4,j2RA7m5Rg2=F>RkL0_k.#d5dH,.+*[g
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mAU=2R>kRF0k_L#5d.H.,d*U[+27,Rm(A52>R=R0Fk_#LkdH.5,*d.[2+(,mR7A25nRR=>F_k0Ldk#.,5Hd[.*+,n2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRA7m5R62=F>RkL0_k.#d5dH,.+*[6R2,75mAc=2R>kRF0k_L#5d.H.,d*c[+27,RmdA52>R=R0Fk_#LkdH.5,*d.[2+d,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7A25.RR=>F_k0Ldk#.,5Hd[.*+,.2RA7m5R42=F>RkL0_k.#d5dH,.+*[4R2,75mAj=2R>kRF0k_L#5d.H.,d*,[2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRu7Qq>R=R_HMs5Cod[n*+Rd68MFI0dFRn+*[d,.2Ru7QA>R=Rj"jj,j"Ru7mq>R=RCFbMR,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRm5uAd=2R>NRbs$H0_#LkdH.5,[c*+,d2Ru7mA25.RR=>bHNs0L$_k.#d5cH,*.[+2R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRm5uA4=2R>NRbs$H0_#LkdH.5,[c*+,42Ru7mA25jRR=>bHNs0L$_k.#d5cH,*2[2;S
SSkSF0C_son5d*R[2<F=RkL0_k.#d5dH,.2*[RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;S
SSkSF0C_son5d*4[+2=R<R0Fk_#LkdH.5,*d.[2+4RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;S
SSkSF0C_son5d*.[+2=R<R0Fk_#LkdH.5,*d.[2+.RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;S
SSkSF0C_son5d*d[+2=R<R0Fk_#LkdH.5,*d.[2+dRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;S
SSkSF0C_son5d*c[+2=R<R0Fk_#LkdH.5,*d.[2+cRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;S
SSkSF0C_son5d*6[+2=R<R0Fk_#LkdH.5,*d.[2+6RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;S
SSkSF0C_son5d*n[+2=R<R0Fk_#LkdH.5,*d.[2+nRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;S
SSkSF0C_son5d*([+2=R<R0Fk_#LkdH.5,*d.[2+(RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;S
SSkSF0C_son5d*U[+2=R<R0Fk_#LkdH.5,*d.[2+URCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;S
SSkSF0C_son5d*g[+2=R<R0Fk_#LkdH.5,*d.[2+gRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;S
SSkSF0C_son5d*4[+j<2R=kRF0k_L#5d.H.,d*4[+jI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';SSSSF_k0s5Cod[n*+244RR<=F_k0Ldk#.,5Hd[.*+244RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;S
SSkSF0C_son5d*4[+.<2R=kRF0k_L#5d.H.,d*4[+.I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';SSSSF_k0s5Cod[n*+24dRR<=F_k0Ldk#.,5Hd[.*+24dRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;S
SSkSF0C_son5d*4[+c<2R=kRF0k_L#5d.H.,d*4[+cI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';SSSSF_k0s5Cod[n*+246RR<=F_k0Ldk#.,5Hd[.*+246RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;S
SSkSF0C_son5d*4[+n<2R=kRF0k_L#5d.H.,d*4[+nI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';SSSSF_k0s5Cod[n*+24(RR<=F_k0Ldk#.,5Hd[.*+24(RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;S
SSkSF0C_son5d*4[+U<2R=kRF0k_L#5d.H.,d*4[+UI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';SSSSF_k0s5Cod[n*+24gRR<=F_k0Ldk#.,5Hd[.*+24gRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;S
SSkSF0C_son5d*.[+j<2R=kRF0k_L#5d.H.,d*.[+jI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';SSSSF_k0s5Cod[n*+2.4RR<=F_k0Ldk#.,5Hd[.*+2.4RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;S
SSkSF0C_son5d*.[+.<2R=kRF0k_L#5d.H.,d*.[+.I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';SSSSF_k0s5Cod[n*+2.dRR<=F_k0Ldk#.,5Hd[.*+2.dRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;S
SSkSF0C_son5d*.[+c<2R=kRF0k_L#5d.H.,d*.[+cI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';SSSSF_k0s5Cod[n*+2.6RR<=F_k0Ldk#.,5Hd[.*+2.6RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;S
SSkSF0C_son5d*.[+n<2R=kRF0k_L#5d.H.,d*.[+nI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';SSSSF_k0s5Cod[n*+2.(RR<=F_k0Ldk#.,5Hd[.*+2.(RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;S
SSkSF0C_son5d*.[+U<2R=kRF0k_L#5d.H.,d*.[+UI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';SSSSF_k0s5Cod[n*+2.gRR<=F_k0Ldk#.,5Hd[.*+2.gRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;S
SSkSF0C_son5d*d[+j<2R=kRF0k_L#5d.H.,d*d[+jI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';SSSSF_k0s5Cod[n*+2d4RR<=F_k0Ldk#.,5Hd[.*+2d4RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;S
SSkSF0C_son5d*d[+.<2R=NRbs$H0_#LkdH.5,[c*2ERIC5MRF_k0CHM52RR='24'R#CDCZR''S;
SFSSks0_Cdo5n+*[dRd2<b=RN0sH$k_L#5d.H*,c[2+4RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;S
SSkSF0C_son5d*d[+c<2R=NRbs$H0_#LkdH.5,[c*+R.2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
SSSS0Fk_osC5*dn[6+d2=R<RsbNH_0$Ldk#.,5Hc+*[dI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';SCSSMo8RCsMCNR0CzNc.;S
SCRM8oCCMsCN0RgzdNS;
CRM8oCCMsCN0RUzdNR;
R8CMRMoCC0sNCcRzd
;
RcRzcRR:H5VRMRF0s8N8sC_soo2RCsMCNR0C-o-RCsMCNR0C#CCDOs0RNRl
R-RR-VRQR8N8s8IH0<ERRN6R#o#HMjR''FR0RkkM#RC8L#H0
RRRRRzjRH:RVNR58I8sHE80R4=R2CRoMNCs0RC
RRRRRDRRFsI_Ns88_<#R=jR"jjjj"RR&s_N8s_Co#25j;R
RRRRRRFRDIN_I8_8s#=R<Rj"jj"jjRI&RNs8_C#o_5;j2
RRRR8CMRMoCC0sNCjRz;R
RR4RzRRR:H5VRNs88I0H8ERR=.o2RCsMCN
0CRRRRRRRRD_FIs8N8sR_#<"=Rjjjj"RR&s_N8s_Co#R548MFI0jFR2R;
RRRRRDRRFII_Ns88_<#R=jR"j"jjRI&RNs8_C#o_584RF0IMF2Rj;R
RRMRC8CRoMNCs0zCR4R;
RzRR.:RRRRHV58N8s8IH0=ERRRd2oCCMsCN0
RRRRRRRRIDF_8sN8#s_RR<="jjj"RR&s_N8s_Co#R5.8MFI0jFR2R;
RRRRRDRRFII_Ns88_<#R=jR"jRj"&NRI8C_so5_#.FR8IFM0R;j2
RRRR8CMRMoCC0sNC.Rz;R
RRdRzRRR:H5VRNs88I0H8ERR=co2RCsMCN
0CRRRRRRRRD_FIs8N8sR_#<"=RjRj"&NRs8C_so5_#dFR8IFM0R;j2
RRRRRRRRIDF_8IN8#s_RR<=""jjRI&RNs8_C#o_58dRF0IMF2Rj;R
RRMRC8CRoMNCs0zCRdS;
z:cSRRHV58N8s8IH0=ERRR62oCCMsCN0
DSSFsI_Ns88_<#R=jR''RR&s_N8s_Co#R5c8MFI0jFR2S;
SIDF_8IN8#s_RR<='Rj'&NRI8C_so5_#cFR8IFM0R;j2
MSC8CRoMNCs0zCRcR;
RzRR6:RRRRHV58N8s8IH0>ERRR62oCCMsCN0
RRRRRRRRIDF_8sN8#s_RR<=s_N8s_Co#R568MFI0jFR2R;
RRRRRDRRFII_Ns88_<#R=NRI8C_so5_#6FR8IFM0R;j2
RRRR8CMRMoCC0sNC6Rz;R

R-RR-VRQRH58MC_sos2RC#oH0RCs7RQhkM#HopRBiR
RRnRzRRR:H5VR8_HMs2CoRMoCC0sNCR
RRRRRRsRbF#OC#BR5pRi,72QhRoLCHRM
RRRRRRRRRHRRVBR5p=iRR''4R8NMRiBp'CCPMR020MEC
RRRRRRRRRRRRRRRR_HMs_Co#=R<Rh7Q;R
RRRRRRRRRRMRC8VRH;R
RRRRRRMRC8sRbF#OC#R;
RCRRMo8RCsMCNR0Cz
n;RRRRzR(R:VRHRF5M0HR8MC_soo2RCsMCN
0CRRRRRRRRRRRRHsM_C#o_RR<=7;Qh
RRRR8CMRMoCC0sNC(Rz;R

R-RR-VRQRF58ks0_CRo2sHCo#s0CRz7ma#RkHRMomiBp
RRRRRzURH:RV8R5F_k0s2CoRMoCC0sNCR
RRRRRRsRbF#OC#mR5B,piR0Fk_osC_R#2LHCoMR
RRRRRRRRRRVRHRB5mp=iRR''4R8NMRpmBiP'CC2M0RC0EMR
RRRRRRRRRRRRRRmR7z<aR=kRF0C_so;_#
RRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMRFbsO#C#;R
RRMRC8CRoMNCs0zCRUR;
RzRRg:RRRRHV50MFRk8F0C_soo2RCsMCN
0CRRRRRRRRRRRR7amzRR<=F_k0s_Co#R;
RCRRMo8RCsMCNR0Cz
g;
RRRRR--Q5VRNs88_osC2CRso0H#CqsR7R7)kM#HopRBiR
RR4Rzj:RRRRHV58sN8ss_CRo2oCCMsCN0
RRRRRRRRFbsO#C#Rp5Bi),Rq)772CRLo
HMRRRRRRRRRRRRH5VRBRpi=4R''MRN8pRBiP'CC2M0RC0EMR
RRRRRRRRRRRRRRNRs8C_soR_#<)=Rq)7758N8s8IH04E-RI8FMR0Fj
2;RRRRRRRRRRRRCRM8H
V;RRRRRRRRCRM8bOsFC;##
RRRR8CMRMoCC0sNC4RzjR;
RzRR4:4RRRHV50MFR8sN8ss_CRo2oCCMsCN0
RRRRRRRRRRRR8sN_osC_<#R=qR)7;7)
RRRR8CMRMoCC0sNC4Rz4
;
RRRR-Q-RVNR58_8ss2CoRosCHC#0s7Rq7k)R#oHMRiBp
RRRR.z4RRR:H5VRI8N8sC_soo2RCsMCN
0CRRRRRRRRbOsFCR##5iBp,qRW727)RoLCHRM
RRRRRRRRRHRRVBR5p=iRR''4R8NMRiBp'CCPMR020MEC
RRRRRRRRRRRRRRRR8IN_osC_<#R=qRW757)Ns88I0H8ER-48MFI0jFR2R;
RRRRRRRRRCRRMH8RVR;
RRRRRCRRMb8RsCFO#
#;RRRRCRM8oCCMsCN0R.z4;R
RR4RzdRR:H5VRMRF0I8N8sC_soo2RCsMCN
0CRRRRRRRRRRRRI_N8s_Co#=R<R7Wq7
);RRRRCRM8oCCMsCN0Rdz4;R
RRRRRRRR
R-RR-CRtMNCs00CRE)CRqOvRC#DDR8NMRD#CCRO0DHFoOR
RR4RzcRR:VRFsHMRHRk5MlC_ODnD_cRR-482RF0IMFRRjoCCMsCN0
RRRRR--Q5VRNs88I0H8ERR>6M2RCRC80OFRs0CNCsRIHR0CCLMNDNCRMF8Rkk0b0MRCNCLDRD#CCRO0DHFoOR
RRRRRR4Rz6RR:H5VRNs88I0H8ERR>no2RCsMCN
0CRRRRRRRRRRRRRRRRF_k0C#M_5RH2<'=R4I'RERCM58sN_osC_N#58I8sHE80-84RF0IMF2RnRH=R2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0C#M_5RH2<W=R ERIC5MRI_N8s_Co#85N8HsI8-0E4FR8IFM0RRn2=2RHR#CDCjR''R;
RRRRRCRRMo8RCsMCNR0Cz;46
RRRRR--Q5VRNs88I0H8E=R<RR62MIFRsCH0RNCMLRDCFFsRkk0b0MRCNCLDRD#CCRO0DHFoOCRMC88C
RRRRRRRRnz4RH:RVNR58I8sHE80RR<=no2RCsMCN
0CRRRRRRRRRRRRRRRRF_k0C#M_5RH2<'=R4
';RRRRRRRRRRRRRRRRI_s0C#M_5RH2<W=R R;
RRRRRCRRMo8RCsMCNR0Cz;4n
RRRRR--tCCMsCN0RC0ERv)qRDOCDN#RM08Rs#H-0CN0#R
RRRRRR4Rz(RR:VRFs[MRHRH5I8R0E-2R4RI8FMR0FjCRoMNCs0RC
RRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)RzqcvnRD:RNDLCRRH#"a17"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloHC5*2ncR"&RW&"RR0HMCsoC'NHlo[C52RR&"R "&MRH0CCosl'HN5oCo_C0C_M880CbEH55+*42nRc,80CbER22&XR""RR&HCM0o'CsHolNC+5[4
2;RRRRRRRRRRRRLHCoMR
RRRRRRRRRR)RzqcvnRX:R)nqvc7X4RR
RRRRRRRRRRRRRRFRbsl0RN5bR7>R=R_HMs_Co#25[,jRqRR=>D_FII8N8s5_#jR2,q=4R>FRDIN_I8_8s#254,.RqRR=>D_FII8N8s5_#.
2,RRRRRRRRRRRRRRRRRRRRRRRRRdRqRR=>D_FII8N8s5_#dR2,q=cR>FRDIN_I8_8s#25c,6RqRR=>D_FII8N8s5_#6R2,
SSSSRSSR)7uq=jR>FRDIN_s8_8s#25j,uR7)Rq4=D>RFsI_Ns88_4#527,Ru.)qRR=>D_FIs8N8s5_#.
2,SSSSSRSR7qu)d>R=RIDF_8sN8#s_5,d2R)7uq=cR>FRDIN_s8_8s#25c,uR7)Rq6=D>RFsI_Ns88_6#52
,RSSSSSRSRW= R>sRI0M_C_H#52W,RBRpi=B>RpRi,7Rum=F>RkL0_kn#_cH#5,2[2;R
RRRRRRRRRRRRRRkRF0C_so5_#[<2R=kRF0k_L#c_n#,5H[I2RERCM50Fk__CM#25HR'=R4R'2CCD#R''Z;R
RRRRRRMRC8CRoMNCs0zCR4
(;RRRRR8CMRMoCC0sNC4RzcR;RRRRRRRRRRRR
RRRRRR
RR-R-RMtCC0sNCRRNdI.RFRs88bCCRv)qRDOCDVRHRbNbssFbHCN0RRRRRRRRRRRRR
RRRRRRzR4U:VRHRk5MlC_ODdD_.RR=4o2RCsMCN
0CRRRR-Q-RVNR58I8sHE80R(>R2CRMC08RFsROCCN0RHIs0CCRMDNLCMRN8kRF00bkRNCMLRDC#CCDOD0RFOoH
RRRRRRRRgz4NRR:H5VRNs88I0H8ERR>no2RCsMCN
0CRRRRRRRRRRRRRRRRF_k0CdM_.=R<R''4RCIEM5R5s_N8s_Co#85N8HsI8-0E4FR8IFM0RRn2=kRMlC_ODnD_cN2RM58Rs_N8s_Co#256R'=Rj2'2R#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_M._dRR<=WI RERCM5N5I8C_so5_#Ns88I0H8ER-48MFI0nFR2RR=M_klODCD_2ncR8NMRN5I8C_so5_#6=2RR''j2C2RDR#C';j'
RRRRRRRR8CMRMoCC0sNC4Rzg
N;RRRRRRRRzL4gRH:RVNR58I8sHE80Rn=RR8NMRlMk_DOCDc_nRj=R2CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_M._dRR<='R4'IMECRs55Ns8_C#o_5R62=jR''R22CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C_Rd.<W=R ERIC5MR58IN_osC_6#52RR='2j'2DRC#'CRj
';RRRRRRRRCRM8oCCMsCN0Rgz4LR;RR-R-RRQV58N8s8IH0<ER=2R6RRMFI0sHCMRCNCLDRRFsFbk0kC0RMDNLCCR#D0CORoDFHMORCCC88R
RRRRRR.RzjRR:H5VRNs88I0H8E=R<RR62oCCMsCN0
RRRRRRRRRRRRRRRR0Fk__CMd<.R=4R''R;
RRRRRRRRRRRRRIRRsC0_M._dRR<=W
 ;RRRRRRRRCRM8oCCMsCN0Rjz.;R
RR-R-RMtCC0sNCER0CqR)vCRODNDRM08Rs#H-0CN0
RRRRRRRR4z.RV:RF[sRRRHM58IH0-ERRR428MFI0jFRRMoCC0sNCR
RRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqz)vRd.:NRDLRCDH"#R1"7aRH&RMo0CCHs'lCNo58IH0RE2&7R""RR&HCM0o'CsHolNCk5MlC_ODnD_cc*n2RR&"RW"&MRH0CCosl'HN5oC[&2RR"" RH&RMo0CCHs'lCNo50oC_8CM_b8C0ME5kOl_C_DDnnc*cRR+dR.,80CbER22&XR""RR&HCM0o'CsHolNC+5[4
2;RRRRRRRRRRRRLHCoMR
RRRRRRRRRR)Rzq.vdRX:R)dqv.7X4RR
RRRRRRRRRRRRRRFRbsl0RN5bR7>R=R_HMs_Co#25[,jRqRR=>D_FII8N8s5_#jR2,q=4R>FRDIN_I8_8s#254,.RqRR=>D_FII8N8s5_#.
2,RRRRRRRRRRRRRRRRRRRRRRRRRdRqRR=>D_FII8N8s5_#dR2,q=cR>FRDIN_I8_8s#25c,SR
SSSSS7RRuj)qRR=>D_FIs8N8s5_#jR2,7qu)4>R=RIDF_8sN8#s_5,42R)7uq=.R>FRDIN_s8_8s#25.,S
SSSSSRuR7)Rqd=D>RFsI_Ns88_d#527,Ruc)qRR=>D_FIs8N8s5_#cR2,
SSSSRSSRRW =I>RsC0_M._d,BRWp=iR>pRBi7,Ru=mR>kRF0k_L#._d#k5MlC_ODdD_.2,[2R;
RRRRRRRRRRRRRFRRks0_C#o_5R[2<F=RkL0_kd#_.M#5kOl_C_DDd[.,2ERIC5MRF_k0CdM_.RR='24'R#CDCZR''R;
RRRRRRRRCRM8oCCMsCN0R4z.;R
RRCRRMo8RCsMCNR0Cz;4URRRRRRRRR
R
RRRR-t-RCsMCNR0CNnR4RsIF8CR8C)bRqOvRCRDDHNVRbFbsbNsH0RCRRRRRRRRRRRRRRR
RR.Rz.RR:H5VRM_klODCD_R4n=2R4RMoCC0sNCR
RR-R-RRQV58N8s8IH0>ERRR62M8CCRR0FONsC0ICRsCH0RNCMLRDCNRM8Fbk0kC0RMDNLCCR#D0CORoDFHRO
RRRRRzRR.RdN:VRHR85N8HsI8R0E>RRnNRM8M_klODCD_Rd.=2R4RMoCC0sNCR
RRRRRRRRRRRRRRkRF0M_C_R4n<'=R4I'RERCM5N5s8C_so5_#Ns88I0H8ER-48MFI0nFR2RR=M_klODCD_2ncR8NMRN5s8C_so5_#6=2RR''42MRN8sR5Ns8_C#o_5Rc2=jR''R22CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C_R4n<W=R ERIC5MR58IN_osC_N#58I8sHE80-84RF0IMF2RnRM=RkOl_C_DDnRc2NRM858IN_osC_6#52RR='24'R8NMRN5I8C_so5_#c=2RR''j2C2RDR#C';j'
RRRRRRRR8CMRMoCC0sNC.Rzd
N;RRRRRRRRzL.dRH:RVNR58I8sHE80Rn>RR8NMRlMk_DOCD._dRR/=4o2RCsMCN
0CRRRRRRRRRRRRRRRRF_k0C4M_n=R<R''4RCIEM5R5s_N8s_Co#85N8HsI8-0E4FR8IFM0RRn2=kRMlC_ODnD_cN2RM58Rs_N8s_Co#256R'=RjR'2NRM858sN_osC_c#52RR='2j'2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0C4M_n=R<RRW IMECRI55Ns8_C#o_58N8s8IH04E-RI8FMR0Fn=2RRlMk_DOCDc_n2MRN8IR5Ns8_C#o_5R62=jR''N2RM58RI_N8s_Co#25cR'=Rj2'2R#CDCjR''R;
RRRRRCRRMo8RCsMCNR0CzL.d;R
RRRRRR.Rzd:ORRRHV58N8s8IH0=ERRNnRMM8RkOl_C_DDd=.RRR42oCCMsCN0
RRRRRRRRRRRRRRRR0Fk__CM4<nR=4R''ERIC5MR58sN_osC_6#52RR='24'R8NMRN5s8C_so5_#c=2RR''j2C2RDR#C';j'
RRRRRRRRRRRRRRRR0Is__CM4<nR= RWRCIEM5R5I_N8s_Co#256R'=R4R'2NRM858IN_osC_c#52RR='2j'2DRC#'CRj
';RRRRRRRRCRM8oCCMsCN0Rdz.OR;
RRRRRzRR.Rd8:VRHR85N8HsI8R0E=RR6NRM8M_klODCD_Rd./4=R2CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_Mn_4RR<='R4'IMECRs55Ns8_C#o_58N8s8IH04E-RI8FMR0Fc=2RRlMk_DOCD._d2C2RDR#C';j'
RRRRRRRRRRRRRRRR0Is__CM4<nR= RWRCIEM5R5I_N8s_Co#85N8HsI8-0E4FR8IFM0RRc2=kRMlC_ODdD_.R22CCD#R''j;R
RRRRRRMRC8CRoMNCs0zCR.;d8RRRR-Q-RVNR58I8sHE80RR<=6M2RFsRIHR0CCLMNDFCRskRF00bkRNCMLRDC#CCDOD0RFOoHRCMC8
C8RRRRRRRRzR.c:VRHR85N8HsI8R0E<c=R2CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_Mn_4RR<=';4'
RRRRRRRRRRRRRRRR0Is__CM4<nR= RW;R
RRRRRRMRC8CRoMNCs0zCR.
c;RRRR-t-RCsMCNR0C0REC)RqvODCDR8NMRH0s-N#00RC
RRRRRzRR.:6RRsVFRH[RMIR5HE80R4-R2FR8IFM0RojRCsMCN
0CRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FzVR)4qvnRR:DCNLD#RHR7"1a&"RR0HMCsoC'NHloIC5HE802RR&"R7"&MRH0CCosl'HN5oCM_klODCD_*ncn+cRRlMk_DOCD._d*2d.R"&RW&"RR0HMCsoC'NHlo[C52RR&"R "&MRH0CCosl'HN5oCo_C0C_M880CbEk5MlC_ODnD_cc*nRM+RkOl_C_DDdd.*.RR+4Rn,80CbER22&XR""RR&HCM0o'CsHolNC+5[4
2;RRRRRRRRRRRRLHCoMR
RRRRRRRRRR)Rzqnv4R):Rqnv4XR47
RRRRRRRRRRRRRRRRsbF0NRlb7R5RR=>HsM_C#o_5,[2RRqj=D>RFII_Ns88_j#52q,R4>R=RIDF_8IN8#s_5,42RRq.=D>RFII_Ns88_.#52R,
RRRRRRRRRRRRRRRRRRRRRRRRRRqd=D>RFII_Ns88_d#527,Ruj)qRR=>D_FIs8N8s5_#jR2,7qu)4>R=RIDF_8sN8#s_5,42R)7uq=.R>FRDIN_s8_8s#25.,S
SSSSSRuR7)Rqd=D>RFsI_Ns88_d#52W,R >R=R0Is__CM4Rn,WiBpRR=>B,piRm7uRR=>F_k0L_k#45n#M_klODCD_,4n[;22
RRRRRRRRRRRRRRRR0Fk_osC_[#52=R<R0Fk_#Lk_#4n5lMk_DOCDn_4,R[2IMECRk5F0M_C_R4n=4R''C2RDR#C';Z'
RRRRRRRR8CMRMoCC0sNC.Rz6R;
RCRRMo8RCsMCNR0Cz;..RRRR
CRRMo8RCsMCNR0Cz;cc
8CMRONsECH0Os0kCDRLF_O	s;Nl
s
NO0EHCkO0sMCRFI_s_COEOF	RVqR)v__)W#RH
lOFbCFMMX0R)dqv.7X4RbRRFRs05R
RRRRRRuR7mRRR:kRF00R#8D_kFOoH;RRRRRRRRR
RRRRRRuR1mRRR:kRF00R#8D_kFOoH;R

RRRRRqRRjRRRRH:RM0R#8D_kFOoH;R
RRRRRR4RqRRRR:MRHR8#0_FkDo;HO
RRRRRRRRRq.R:RRRRHM#_08koDFH
O;RRRRRRRRqRdRRRR:H#MR0k8_DHFoOR;
RRRRRqRRcRRRRH:RM0R#8D_kFOoH;R
RRRRRRRR7RRRR:MRHR8#0_FkDo;HO
RRRRRRRR)7uq:jRRRHM#_08koDFH
O;RRRRRRRR7qu)4RR:H#MR0k8_DHFoOR;
RRRRR7RRu.)qRH:RM0R#8D_kFOoH;R
RRRRRRuR7)Rqd:MRHR8#0_FkDo;HO
RRRRRRRR)7uq:cRRRHM#_08koDFH
O;RRRRRRRRWiBpRRR:H#MR0k8_DHFoOR;RRRRRRRR
RRRRRWRR RRRRH:RM0R#8D_kFOoH
RRRRRRR2R;R
8CMRlOFbCFMM
0;ObFlFMMC0)RXqcvnXR47RFRbs50R
RRRRRRRRm7uR:RRR0FkR8#0_FkDo;HORRRRRRRR
RRRRRRRRm1uR:RRR0FkR8#0_FkDo;HO
R
RRRRRRjRqRRRR:MRHR8#0_FkDo;HO
RRRRRRRRRq4R:RRRRHM#_08koDFH
O;RRRRRRRRqR.RRRR:H#MR0k8_DHFoOR;
RRRRRqRRdRRRRH:RM0R#8D_kFOoH;R
RRRRRRcRqRRRR:MRHR8#0_FkDo;HO
RRRRRRRRRq6R:RRRRHM#_08koDFH
O;RRRRRRRR7RRRRRR:H#MR0k8_DHFoOR;
RRRRR7RRuj)qRH:RM0R#8D_kFOoH;R
RRRRRRuR7)Rq4:MRHR8#0_FkDo;HO
RRRRRRRR)7uq:.RRRHM#_08koDFH
O;RRRRRRRR7qu)dRR:H#MR0k8_DHFoOR;
RRRRR7RRuc)qRH:RM0R#8D_kFOoH;R
RRRRRRuR7)Rq6:MRHR8#0_FkDo;HO
RRRRRRRRpWBi:RRRRHM#_08koDFHRO;RRRRR
RRRRRRRRRRWR RRRR:H#MR0k8_DHFoOR
RRRRRRR2;RM
C8FROlMbFC;M0
MVkOF0HMkRVMHO_M5H0LRR:LDFFC2NMR0sCkRsM#H0sMHoR#C
Lo
HMRVRHR25LRC0EMR
RRCRs0Mks5F"hRNsC8s/IHR0COVFMD0HORCOEOR	31kHlDHN0FlMRHN#l0ROEb#F#HCLDR"!!2R;
R#CDCR
RRCRs0Mks5F"BkRD8MRF0HDlbCMlC0DRAFRO	)3qvRRQ#0RECs8CNR8N8s#C#RosCHC#0sRC8kM#HoER0CNR#lOCRD	FORRN#0REC)?qv"
2;RMRC8VRH;M
C8kRVMHO_M;H0
MVkOF0HMCRo0M_C8C_8b50E#CHxRH:RMo0CC;sRRb8C0:ERR0HMCsoC2CRs0MksR0HMCsoCR
H#PHNsNCLDRMlH_x#HCRR:HCM0oRCs:j=R;C
Lo
HMRHRlMH_#x:CR=CR8b;0E
HRRV#R5HRxC<CR8b20ERC0EMR
RRHRlMH_#x:CR=HR#x
C;RMRC8VRH;R
RskC0slMRH#M_H;xC
8CMR0oC_8CM_b8C0
E;Ns00H0LkCCRoMNCs0_FssFCbs:0RRs#0H;Mo
0N0skHL0oCRCsMCNs0F_bsCFRs0FMVRFI_s_COEO:	RRONsECH0Os0kC#RHRMVkOM_HHs05Ns88_osC2-;
-CRLoRHMLODF	NRsllRHblDCCNM00MHFRo#HM#ND
b0$CMRH0s_NsRN$HN#Rs$sNRR5j06FR2VRFR0HMCsoC;F
OMN#0MI0RHE80_sNsN:$RR0HM_sNsN:$R=4R5,,R.RRc,g4,RUd,Rn
2;O#FM00NMRb8C0NE_s$sNRH:RMN0_s$sNRR:=5d4nURc,U.4g,jRcgRn,.Ujc,jR4.Rc,624.;F
OMN#0M80RH.PdRH:RMo0CC:sR=IR5HE80-/42d
n;O#FM00NMRP8H4:nRR0HMCsoCRR:=58IH04E-2U/4;F
OMN#0M80RHRPU:MRH0CCos=R:RH5I8-0E4g2/;F
OMN#0M80RHRPc:MRH0CCos=R:RH5I8-0E4c2/;F
OMN#0M80RHRP.:MRH0CCos=R:RH5I8-0E4.2/;F
OMN#0M80RHRP4:MRH0CCos=R:RH5I8-0E442/;O

F0M#NRM0LDFF4RR:LDFFCRNM:5=R84HPRj>R2O;
F0M#NRM0LDFF.RR:LDFFCRNM:5=R8.HPRj>R2O;
F0M#NRM0LDFFcRR:LDFFCRNM:5=R8cHPRj>R2O;
F0M#NRM0LDFFURR:LDFFCRNM:5=R8UHPRj>R2O;
F0M#NRM0LDFF4:nRRFLFDMCNRR:=5P8H4>nRR;j2
MOF#M0N0FRLF.DdRL:RFCFDN:MR=8R5H.PdRj>R2
;
O#FM00NMRP8H4UndcRR:HCM0oRCs:5=R80CbE2-4/d4nU
c;O#FM00NMRP8HU.4gRH:RMo0CC:sR=8R5CEb0-/42U.4g;F
OMN#0M80RHjPcg:nRR0HMCsoCRR:=5b8C04E-2j/cg
n;O#FM00NMRP8H.UjcRH:RMo0CC:sR=8R5CEb0-/42.Ujc;F
OMN#0M80RHjP4.:cRR0HMCsoCRR:=5b8C04E-2j/4.
c;O#FM00NMRP8H6R4.:MRH0CCos=R:RC58b-0E462/4
.;
MOF#M0N0FRLF4D6.RR:LDFFCRNM:5=R86HP4>.RR;j2
MOF#M0N0FRLFjD4.:cRRFLFDMCNRR:=5P8H4cj.Rj>R2O;
F0M#NRM0LDFF.UjcRL:RFCFDN:MR=8R5HjP.c>URR;j2
MOF#M0N0FRLFjDcg:nRRFLFDMCNRR:=5P8HcnjgRj>R2O;
F0M#NRM0LDFFU.4gRL:RFCFDN:MR=8R5H4PUg>.RR;j2
MOF#M0N0FRLFnD4dRUc:FRLFNDCM=R:RH58Pd4nU>cRR;j2
F
OMN#0M#0RkIl_HE80RH:RMo0CC:sR=mRAmqp hF'b#F5LF2D4RA+Rm mpqbh'FL#5F.FD2RR+Apmm 'qhb5F#LDFFc+2RRmAmph q'#bF5FLFDRU2+mRAmqp hF'b#F5LFnD42O;
F0M#NRM0#_kl80CbERR:HCM0oRCs:6=RR5-RApmm 'qhb5F#LDFF624.RA+Rm mpqbh'FL#5F4FDj2.cRA+Rm mpqbh'FL#5F.FDj2cURA+Rm mpqbh'FL#5FcFDj2gnRA+Rm mpqbh'FL#5FUFD42g.2
;
O#FM00NMROI_EOFHCH_I8R0E:MRH0CCos=R:R8IH0NE_s$sN5l#k_8IH0;E2
MOF#M0N0_RIOHEFO8C_CEb0RH:RMo0CC:sR=CR8b_0ENNss$k5#lH_I820E;F
OMN#0M80R_FOEH_OCI0H8ERR:HCM0oRCs:I=RHE80_sNsN#$5k8l_CEb02O;
F0M#NRM08E_OFCHO_b8C0:ERR0HMCsoCRR:=80CbEs_Ns5N$#_kl80CbE
2;
MOF#M0N0_RII0H8Ek_MlC_ODRD#:MRH0CCos=R:RH5I8-0E4I2/_FOEH_OCI0H8ERR+4O;
F0M#NRM0IC_8b_0EM_klODCD#RR:HCM0oRCs:5=R80CbE2-4/OI_EOFHCC_8bR0E+;R4
F
OMN#0M80R_8IH0ME_kOl_C#DDRH:RMo0CC:sR=IR5HE80-/428E_OFCHO_8IH0+ERR
4;O#FM00NMR88_CEb0_lMk_DOCD:#RR0HMCsoCRR:=5b8C04E-2_/8OHEFO8C_CEb0R4+R;O

F0M#NRM0IH_#x:CRR0HMCsoCRR:=IH_I8_0EM_klODCD#RR*IC_8b_0EM_klODCD#O;
F0M#NRM08H_#x:CRR0HMCsoCRR:=8H_I8_0EM_klODCD#RR*8C_8b_0EM_klODCD#
;
O#FM00NMRFLFDR_8:FRLFNDCM=R:R_58#CHxRI-R_x#HC=R<R;j2
MOF#M0N0FRLFID_RL:RFCFDN:MR=FRM0F5LF8D_2
;
O#FM00NMRFOEH_OCI0H8ERR:HCM0oRCs:5=RApmm 'qhb5F#LDFF_R82*_R8OHEFOIC_HE802RR+5mAmph q'#bF5FLFD2_IRI*R_FOEH_OCI0H8E
2;O#FM00NMRFOEH_OC80CbERR:HCM0oRCs:5=RApmm 'qhb5F#LDFF_R82*_R8OHEFO8C_CEb02RR+5mAmph q'#bF5FLFD2_IRI*R_FOEH_OC80CbE
2;O#FM00NMR8IH0ME_kOl_C#DDRH:RMo0CC:sR=AR5m mpqbh'FL#5F_FD8*2R58IH04E-2_/8OHEFOIC_HE802RR+5mAmph q'#bF5FLFD2_IR5*RI0H8E2-4/OI_EOFHCH_I820ER4+R;F
OMN#0M80RCEb0_lMk_DOCD:#RR0HMCsoCRR:=5mAmph q'#bF5FLFD2_8R8*5CEb0-/428E_OFCHO_b8C0RE2+AR5m mpqbh'FL#5F_FDI*2RRC58b-0E4I2/_FOEH_OC80CbE+2RR
4;0C$bR0Fk_#Lk4$_0bHCR#sRNsRN$5b8C0ME_kOl_C#DD-84RF0IMF,RjR8IH0ME_kOl_C#DD-84RF0IMF2RjRRFV#_08DHFoO#;
HNoMDkRF0k_L#:4RR0Fk_#Lk4$_0bRC;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RV_Rs80FkRM5HbRk000FRs#H-0CN0#02
$RbCF_k0L.k#_b0$C#RHRsNsN5$R80CbEk_MlC_OD-D#4FR8IFM0RRj,.H*I8_0EM_klODCD#R+48MFI0jFR2VRFR8#0_oDFH
O;#MHoNFDRkL0_kR#.:kRF0k_L#0._$;bCRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$FsVR_k8F0HR5M0bkRR0F0-sH#00NC
#20C$bR0Fk_#Lkc$_0bHCR#sRNsRN$5b8C0ME_kOl_C#DD-84RF0IMF,RjRIc*HE80_lMk_DOCDd#+RI8FMR0FjF2RV0R#8F_Do;HO
o#HMRNDF_k0Lck#RF:RkL0_k_#c0C$b;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFVsF_8k50RHkMb0FR0RH0s-N#002C#
b0$CkRF0k_L#0U_$RbCHN#Rs$sNRC58b_0EM_klODCD#R-48MFI0jFR,*RUI0H8Ek_MlC_OD+D#(FR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNR0Fk_#LkURR:F_k0LUk#_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFR8s_FRk05bHMk00RFsR0H0-#N#0C2$
0bbCRN0sH$k_L#0U_$RbCHN#Rs$sNRC58b_0EM_klODCD#R-48MFI0jFR,HRI8_0EM_klODCD#R-48MFI0jFR2VRFR8#0_oDFH
O;#MHoNbDRN0sH$k_L#:URRsbNH_0$LUk#_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$FsVR_k8F0HR5M0bkRR0F0-sH#00NC
#20C$bR0Fk_#Lk40n_$RbCHN#Rs$sNRC58b_0EM_klODCD#R-48MFI0jFR,nR4*8IH0ME_kOl_C#DD+R468MFI0jFR2VRFR8#0_oDFH
O;#MHoNFDRkL0_kn#4RF:RkL0_kn#4_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFR8s_FRk05bHMk00RFsR0H0-#N#0C2$
0bbCRN0sH$k_L#_4n0C$bRRH#NNss$8R5CEb0_lMk_DOCD4#-RI8FMR0Fj.,R*8IH0ME_kOl_C#DD+84RF0IMF2RjRRFV#_08DHFoO#;
HNoMDNRbs$H0_#Lk4:nRRsbNH_0$L4k#n$_0bRC;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RV_Rs80FkRM5HbRk000FRs#H-0CN0#02
$RbCF_k0Ldk#.$_0bHCR#sRNsRN$5b8C0ME_kOl_C#DD-84RF0IMF,RjR*d.I0H8Ek_MlC_OD+D#d84RF0IMF2RjRRFV#_08DHFoO#;
HNoMDkRF0k_L#Rd.:kRF0k_L#_d.0C$b;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFVsF_8k50RHkMb0FR0RH0s-N#002C#
b0$CNRbs$H0_#Lkd0._$RbCHN#Rs$sNRC58b_0EM_klODCD#R-48MFI0jFR,*RcI0H8Ek_MlC_OD+D#dFR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNRsbNH_0$Ldk#.RR:bHNs0L$_k.#d_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFR8s_FRk05bHMk00RFsR0H0-#N#0C2H
#oDMNR0Fk_RCM:0R#8F_Do_HOP0COF8s5CEb0_lMk_DOCD4#-RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-C-RMDNLCV#RF0sRs#H-0CN0#H
#oDMNR0Is_RCM:0R#8F_Do_HOP0COF8s5CEb0_lMk_DOCD4#-RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-I-RsCH0RNCML#DCRsVFROCNEFRsIVRFRv)qRDOCD##
HNoMDMRH_osCR#:R0D8_FOoH_OPC05FsI0H8E6+dRI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RCk#8FR0RosCHC#0sQR7h#R
HNoMDkRF0C_soRR:#_08DHFoOC_POs0F58IH0dE+6FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RCk#8FR0RosCHC#0smR7z#a
HNoMDkRF0C_so:4RR8#0_oDFHPO_CFO0sH5I8-0E4FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--k8#CRR0FOFEF#LCRCC0IC7MRQNhRMF8Rkk0b0VRFRFADO)	Rq#v
HNoMDNRs8C_soRR:#_08DHFoOC_POs0F58N8s8IH04E-RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RCk#8FR0RosCHC#0sqR)7
7)#MHoNIDRNs8_C:oRR8#0_oDFHPO_CFO0s85N8HsI8-0E4FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-#RkC08RFCRso0H#CWsRq)77
o#HMRNDD_FIs8N8sRR:#_08DHFoOC_POs0F5R4d8MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--s8N8sHRL0H#RM0bkRR0F)RqvODCD#cR5R0LH#CRsJskHC
82#MHoNDDRFII_Ns88R#:R0D8_FOoH_OPC05Fs48dRF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-I-RNs88R0LH#MRHbRk00)FRqOvRC#DDRR5cL#H0RJsCkCHs8#2
HNoMD_RsNs88_osCR#:R0D8_FOoH_OPC05FsNs88I0H8ER-48MFI0jFR2-;
-MRC8DRLFRO	sRNlHDlbCMlC0HN0F#MRHNoMD-#
-CRLoRHM#CCDOs0RNHlRlCbDl0CMNF0HMHR#oDMN#k
VMHO0FoMRCM0_knl_cC58b:0ER0HMCsoC2CRs0MksR0HMCsoCR
H#PHNsNCLDRDPNRH:RMo0CC:sR=;Rj
oLCHRM
RDPNRR:=80CbEc/n;R
RH5VR5b8C0lERFn8Rc>2RR2cURC0EMR
RRNRPD=R:RDPNR4+R;R
RCRM8H
V;RCRs0MksRDPN;M
C8CRo0k_Mlc_n;k
VMHO0FoMRCD0_CFV0P_Csd8.5CEb0RH:RMo0CCRs2skC0sHMRMo0CCHsR#C
Lo
HMRCRs0Mks5b8C0lERFn8Rc
2;CRM8o_C0D0CVFsPC_;d.
MVkOF0HMCRo0C_DVP0FC8s5CEb0RH:RMo0CCRs;lRNG:MRH0CCoss2RCs0kMMRH0CCos#RH
sPNHDNLCNRPDRR:HCM0oRCs:j=R;C
Lo
HMRVRHRC58bR0E-NRlG=R>RRj20MEC
RRRRDPNRR:=80CbERR-l;NG
CRRD
#CRRRRPRND:8=RCEb0;R
RCRM8H
V;RCRs0Mks5DPN2C;
Mo8RCD0_CFV0P;Cs
MVkOF0HMCRo0k_Ml._d5b8C0:ERR0HMCsoC2CRs0MksR0HMCsoCR
H#PHNsNCLDRDPNRH:RMo0CC:sR=;Rj
oLCHRM
RRHV5b8C0<ER=URcR8NMRb8C0>ERR24nRC0EMR
RRPRRN:DR=;R4
CRRMH8RVR;
R0sCkRsMP;ND
8CMR0oC_lMk_;d.
MVkOF0HMCRo0k_Mln_45b8C0:ERR0HMCsoC2CRs0MksR0HMCsoCR
H#PHNsNCLDRDPNRH:RMo0CC:sR=;Rj
oLCHRM
RRHV5b8C0<ER=nR4R8NMRb8C0>ERRRj20MEC
RRRRNRPD=R:R
4;RMRC8VRH;R
RskC0sPMRN
D;CRM8o_C0M_kl4
n;O#FM00NMRlMk_DOCDc_nRH:RMo0CC:sR=CRo0k_Mlc_n5b8C0;E2
MOF#M0N0CRDVP0FCds_.RR:HCM0oRCs:o=RCD0_CFV0P_Csd8.5CEb02O;
F0M#NRM0M_klODCD_Rd.:MRH0CCos=R:R0oC_lMk_5d.D0CVFsPC_2d.;F
OMN#0MD0RCFV0P_Cs4:nRR0HMCsoCRR:=o_C0D0CVFsPC5VDC0CFPs._d,.Rd2O;
F0M#NRM0M_klODCD_R4n:MRH0CCos=R:R0oC_lMk_54nD0CVFsPC_24n;0

$RbCF_k0L_k#0C$b_#ncRRH#NNss$MR5kOl_C_DDn8cRF0IMF,RjR8IH04E-RI8FMR0FjF2RV0R#8F_Do;HO
b0$CkRF0k_L#$_0bdC_.H#R#sRNsRN$5lMk_DOCD._dRI8FMR0FjI,RHE80-84RF0IMF2RjRRFV#_08DHFoO0;
$RbCF_k0L_k#0C$b_#4nRRH#NNss$MR5kOl_C_DD48nRF0IMF,RjR8IH04E-RI8FMR0FjF2RV0R#8F_Do;HO
o#HMRNDF_k0L_k#nRc#:kRF0k_L#$_0bnC_cR#;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RVFR8k50RHkMb0FR0RH0s-N#002C#
o#HMRNDF_k0L_k#dR.#:kRF0k_L#$_0bdC_.R#;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RVFR8k50RHkMb0FR0RH0s-N#002C#
o#HMRNDF_k0L_k#4Rn#:kRF0k_L#$_0b4C_nR#;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RVFR8k50RHkMb0FR0RH0s-N#002C#
o#HMRNDF_k0C#M_R#:R0D8_FOoH_OPC05FsM_klODCD_Rnc8MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-MRCNCLD#FRVssR0H0-#N#0C
o#HMRNDF_k0CdM_.RR:#_08DHFoO#;
HNoMDkRF0M_C_R4n:0R#8F_Do;HO
o#HMRNDI_s0C#M_R#:R0D8_FOoH_OPC05FsM_klODCD_Rnc8MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-sRIHR0CCLMNDRC#VRFsCENORIsFRRFV)RqvODCD#H
#oDMNR0Is__CMd:.RR8#0_oDFH
O;#MHoNIDRsC0_Mn_4R#:R0D8_FOoH;H
#oDMNR_HMs_Co#RR:#_08DHFoOC_POs0F58IH04E-RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RCk#8FR0RosCHC#0sQR7h#R
HNoMDkRF0C_soR_#:0R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-#RkC08RFCRso0H#C7sRm
za#MHoNsDRNs8_C#o_R#:R0D8_FOoH_OPC05FsNs88I0H8ER-48MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--k8#CRR0FsHCo#s0CR7q7)H
#oDMNR8IN_osC_:#RR8#0_oDFHPO_CFO0s85N8HsI8-0E4FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-#RkC08RFCRso0H#CqsR7
7)#MHoNDDRFsI_Ns88_:#RR8#0_oDFHPO_CFO0sR568MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--Ns88R0LH#MRHbRk00)FRqOvRC#DDRR5cL#H0RJsCkCHs8#2
HNoMDFRDIN_I8_8s#RR:#_08DHFoOC_POs0F586RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-N-R8R8sL#H0RbHMk00RFqR)vCRODRD#5LcRHR0#skCJH8sC2-
-R8CMRD#CCRO0sRNlHDlbCMlC0HN0F#MRHNoMDN#
0H0sLCk0Rs\3NFl_VCV#0:\RRs#0H;Mo
C
Lo
HMRcRzdH:RVsR5Ns88_osC2CRoMNCs0-CR-CRoMNCs0LCRD	FORlsN
RRRRR--QNVR8I8sHE80RO<REOFHCH_I8R0ENH##o'MRj0'RFMRkk8#CR0LH#R
RRjRzRRR:H5VRNs88I0H8ERR=4o2RCsMCN
0CSRRRRIDF_8sN8<sR=jR"jjjjjjjjjjjj"RR&s_N8s5Coj
2;SRRRRIDF_8IN8<sR=jR"jjjjjjjjjjjj"RR&I_N8s5Coj
2;S8CMRMoCC0sNCjRz;R
RR4RzRRR:H5VRNs88I0H8ERR=.o2RCsMCN
0CSFSDIN_s8R8s<"=Rjjjjjjjjjjjj"RR&s_N8s5Co4FR8IFM0R;j2
RSRRFRDIN_I8R8s<"=Rjjjjjjjjjjjj"RR&I_N8s5Co4FR8IFM0R;j2
MSC8CRoMNCs0zCR4R;
RzRR.:RRRRHV58N8s8IH0=ERRRd2oCCMsCN0
DSSFsI_Ns88RR<="jjjjjjjjjjj"RR&s_N8s5Co.FR8IFM0R;j2
RSRRFRDIN_I8R8s<"=Rjjjjjjjjj"jjRI&RNs8_C.o5RI8FMR0Fj
2;S8CMRMoCC0sNC.Rz;R
RRdRzRRR:H5VRNs88I0H8ERR=co2RCsMCN
0CSFSDIN_s8R8s<"=RjjjjjjjjjRj"&NRs8C_soR5d8MFI0jFR2S;
RRRRD_FII8N8s=R<Rj"jjjjjjjjj"RR&I_N8s5CodFR8IFM0R;j2
MSC8CRoMNCs0zCRdR;
RzRRc:RRRRHV58N8s8IH0=ERRR62oCCMsCN0
RSRRFRDIN_s8R8s<"=Rjjjjjjjjj&"RR8sN_osC58cRF0IMF2Rj;R
SRDRRFII_Ns88RR<="jjjjjjjjRj"&NRI8C_soR5c8MFI0jFR2S;
CRM8oCCMsCN0R;zc
RRRRRz6RH:RVNR58I8sHE80Rn=R2CRoMNCs0SC
RRRRD_FIs8N8s=R<Rj"jjjjjjRj"&NRs8C_soR568MFI0jFR2S;
SIDF_8IN8<sR=jR"jjjjj"jjRI&RNs8_C6o5RI8FMR0Fj
2;S8CMRMoCC0sNC6Rz;R
RRnRzRRR:H5VRNs88I0H8ERR=(o2RCsMCN
0CSRRRRIDF_8sN8<sR=jR"jjjjjRj"&NRs8C_soR5n8MFI0jFR2S;
SIDF_8IN8<sR=jR"jjjjjRj"&NRI8C_soR5n8MFI0jFR2S;
CRM8oCCMsCN0R;zn
RRRRRz(RH:RVNR58I8sHE80RU=R2CRoMNCs0SC
RRRRD_FIs8N8s=R<Rj"jjjjj"RR&s_N8s5Co(FR8IFM0R;j2
DSSFII_Ns88RR<="jjjj"jjRI&RNs8_C(o5RI8FMR0Fj
2;S8CMRMoCC0sNC(Rz;R
RRURzRRR:H5VRNs88I0H8ERR=go2RCsMCN
0CSRRRRIDF_8sN8<sR=jR"jjjj"RR&s_N8s5CoUFR8IFM0R;j2
DSSFII_Ns88RR<="jjjjRj"&NRI8C_soR5U8MFI0jFR2S;
CRM8oCCMsCN0R;zU
RRRRRzgRH:RVNR58I8sHE80R4=Rjo2RCsMCN
0CSRRRRIDF_8sN8<sR=jR"j"jjRs&RNs8_Cgo5RI8FMR0Fj
2;SFSDIN_I8R8s<"=Rjjjj"RR&I_N8s5CogFR8IFM0R;j2
MSC8CRoMNCs0zCRgR;
RzRR4RjR:VRHR85N8HsI8R0E=4R42CRoMNCs0SC
RRRRD_FIs8N8s=R<Rj"jj&"RR8sN_osC5R4j8MFI0jFR2S;
SIDF_8IN8<sR=jR"jRj"&NRI8C_soj54RI8FMR0Fj
2;S8CMRMoCC0sNC4RzjR;
RzRR4R4R:VRHR85N8HsI8R0E=.R42CRoMNCs0SC
RRRRD_FIs8N8s=R<Rj"j"RR&s_N8s5Co484RF0IMF2Rj;S
SD_FII8N8s=R<Rj"j"RR&I_N8s5Co484RF0IMF2Rj;C
SMo8RCsMCNR0Cz;44
RRRR.z4RRR:H5VRNs88I0H8ERR=4Rd2oCCMsCN0
RSRRFRDIN_s8R8s<'=Rj&'RR8sN_osC5R4.8MFI0jFR2S;
SIDF_8IN8<sR=jR''RR&I_N8s5Co48.RF0IMF2Rj;C
SMo8RCsMCNR0Cz;4.
RRRRdz4RRR:H5VRNs88I0H8ERR>4Rd2oCCMsCN0
RSRRFRDIN_s8R8s<s=RNs8_C4o5dFR8IFM0R;j2
RSRRFRDIN_I8R8s<I=RNs8_C4o5dFR8IFM0R;j2
MSC8CRoMNCs0zCR4
d;
RRRRR--Q5VR8_HMs2CoRosCHC#0sQR7h#RkHRMoB
piRRRRzR4cRH:RV8R5HsM_CRo2oCCMsCN0
RRRRRRRRFbsO#C#Rp5Bi7,RQRh2LHCoMR
RRRRRRRRRRVRHRp5BiRR='R4'NRM8B'piCMPC002RE
CMRRRRRRRRRRRRRRRRHsM_C<oR="R5jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"RR&72Qh;R
RRRRRRRRRRMRC8VRH;R
RRRRRRMRC8sRbF#OC#S;
CRM8oCCMsCN0Rcz4;R
RR4Rz6:RRRRHV50MFRM8H_osC2CRoMNCs0RC
RRRRRRRRRHRRMC_so=R<Rj5"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jjR7&RQ;h2
MSC8CRoMNCs0zCR4
6;
RRRRR--Q5VRsk8F0C_sos2RC#oH0RCs)m_7zkaR#oHMRm)_B
piRRRRzR4nRH:RV8R5F_k0s2CoRMoCC0sNCR
RRRRRRsRbF#OC#mR5B,piR0Fk_osC4L2RCMoH
RRRRRRRRRRRRRHV5pmBiRR='R4'NRM8miBp'CCPMR020MEC
RRRRRRRRRRRRRRRRz7ma=R<R0Fk_osC4R;
RRRRRRRRRCRRMH8RVR;
RRRRRCRRMb8RsCFO#
#;RRRRRRRRCRM8oCCMsCN0Rnz4;R
RR4Rz(:RRRRHV50MFRk8F0C_soo2RCsMCN
0CRRRRRRRRRRRR7amzRR<=F_k0s4Co;C
SMo8RCsMCNR0Cz;4(
R
RR-R-RRQV58sN8ss_CRo2sHCo#s0CR7)q7k)R#oHMRpmBiR
RR4RznRsR:VRHRN5s8_8ss2CoRMoCC0sNC-
-RRRRRRRRbOsFCR##5pmBi),Rq)772CRLo
HM-R-RRRRRRRRRRVRHRB5mp=iRR''4R8NMRpmBiP'CC2M0RC0EM-
-RRRRRRRRRRRRRRRRs_N8sRCo<)=Rq)7758N8s8IH04E-RI8FMR0Fj
2;-R-RRRRRRRRRRMRC8VRH;-
-RRRRRRRRCRM8bOsFC;##
S--CRM8oCCMsCN0Rnz4s-;
-RRRR(z4sRR:H5VRMRF0s8N8sC_soo2RCsMCN
0CRRRRRRRRRRRRs_N8sRCo<)=Rq)77;C
SMo8RCsMCNR0Czs4n;S

-Q-RVIR5Ns88_osC2CRso0H#CWsRq)77RHk#MWoR_pmBiR
RR4RznRIR:VRHRN5I8_8ss2CoRMoCC0sNCR
RRRRRRsRbF#OC#BR5pRi,W7q7)L2RCMoH
RRRRRRRRRRRRRHV5iBpR'=R4N'RMB8RpCi'P0CM2ER0CRM
RRRRRRRRRRRRRIRRNs8_C<oR=qRW757)Ns88I0H8ER-48MFI0jFR2R;
RRRRRRRRRCRRMH8RVR;
RRRRRCRRMb8RsCFO#
#;S8CMRMoCC0sNC4Rzn
I;RRRRzI4(RH:RVMR5FI0RNs88_osC2CRoMNCs0RC
RRRRRRRRRIRRNs8_C<oR=qRW7;7)
MSC8CRoMNCs0zCR4;(I
R
RR-R-R0 GsDNRFOoHRsVFRN7kDFRbsO0RN
#CSR--7MFRFM0RCRC80#EHRsVFRsMF8OIsEO	RN
#C-z-SsRCo:sRbF#OC#p5BiL2RCMoH
S--RVRHRp5Bie'  RhaNRM8BRpi=4R''02RE
CM-R-SRQR7hl_0b=R<Rh7Q;-
-SRRR)7q7)l_0b=R<R7)q7
);-R-SRqRW7_7)0Rlb<W=Rq)77;-
-SRRRW0 _l<bR= RW;-
-SCRRMH8RV-;
-MSC8sRbF#OC#
;
SR--Q)VRCRN8qs88CR##=sRWHR0Cqs88C,##RbL$NR##7RQh0FFRkk0b0VRHRRW HC#RMDNLCS8
zGlkRb:RsCFO#F#5ks0_C
o2SLRRCMoH
S--RRRRH5VRW7q7)l_0bRR=)7q7)l_0bMRN8 RW_b0lR'=R4R'20MEC
S--SFRRks0_CRo4<7=RQ0h_l
b;-S-SCCD#
RSSR0Fk_osC4=R<R0Fk_osC58IH04E-RI8FMR0Fj
2;-S-SCRM8H
V;S8CMRFbsO#C#;R
SR
RRRRRR-t-RCsMCNR0C0REC)RqvODCD#MRN8CR#D0CORoDFHVORF)sRq4vAn4_1_
14SUz4RH:RVOR5EOFHCH_I8R0E=2R4RMoCC0sNC-
S-HRVGFRVsNROD4DRd(UU,CR#D0CORRFV0#sH0CN0R0MFRHLCMsoRC#oH0CCs8R
SRORzER	:H5VRNs88I0H8ERR>4Rc2oCCMsCN0
RRRRRRRRDkO	RR:bOsFC5##B2pi
RRRRRRRRCRLo
HMRRRRRRRRRVRHRp5BiP'CCRM0NRM8BRpi=4R''02RE
CMRRRRRRRRRRRRs8_N8ss_CNo58I8sHE80-84RF0IMFcR42=R<R7)q7N)58I8sHE80-84RF0IMFcR42R;
RRRRRRRRR8CMR;HV
RRRRRRRR8CMRFbsO#C#RDkO	S;
RMRC8CRoMNCs0zCRO;E	
RRRR4SzgRR:VRFsHMRHRC58b_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
-S-RRQV58N8s8IH0>ERR24cRCMC8FR0RCOsNR0CI0sHCMRCNCLDR8NMR0FkbRk0CLMND#CRCODC0FRDo
HORRRRRRRRSjz.RH:RVNR58I8sHE80R4>Rco2RCsMCN
0CSR--VRHGVRFsODNDRU4dUR(,#CCDOF0RVsR0HN#00MCRFL0RCoHMRosCHC#0s
C8SSSSF_k0CHM52=R<R''4RCIEMsR5_8N8sC_so85N8HsI8-0E4FR8IFM0R24cRH=R2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0CHM52=R<RRW IMECRN5I8C_so85N8HsI8-0E4FR8IFM0R24cRH=R2DRC#'CRj
';RRRRRRRRS8CMRMoCC0sNC.RzjS;
-Q-RVNR58I8sHE80RR<=4Rc2MIFRsCH0RNCMLRDCFFsRkk0b0MRCNCLDRD#CCRO0DHFoOCRMC88C
RRSRSRRzR.4:VRHR85N8HsI8R0E<4=Rco2RCsMCN
0CSSSSF_k0CHM52=R<R''4;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R R;
RRRRRSRRCRM8oCCMsCN0R4z.;-
S-CRtMNCs00CRE)CRqOvRC#DDR8NMRH0s-N#00
C#RRRRRRRRS.z.RV:RF[sRRRHM58IH0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CRRRRRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FAVR)_qv4Undc7X4RD:RNDLCRRH#";W"
RRRRRRRRRRRRRRRRoLCHRM
RRRRRRRRRSRRAv)q_d4nU4cX7RR:)Aqv41n_44_1
RSRRRRRRRRRRFRbsl0RN5bR75Qqj=2R>MRH_osC5,[2R7q7)=qR>FRDIN_I858s48dRF0IMF2Rj,QR7A>R=R""j,7Rq7R)A=D>RFsI_Ns885R4d8MFI0jFR2S,
S SSh=qR>4R''1,R1R)q='>RjR',WR q=I>RsC0_M25H,pRBi=qR>pRBi ,Rh=AR>4R''1,R1R)A='>RjR',WR A='>RjR',BApiRR=>B,pi
SSSRRRR7Rmq=F>Rb,CMRA7m5Rj2=F>RkL0_k5#4H2,[2
;
RRRRRRRRRRRRRRRRF_k0s5Co[<2R=kRF0k_L#H45,R[2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRMSC8CRoMNCs0zCR.
.;RRRRRMSC8CRoMNCs0zCR4
g;RRRRCRM8oCCMsCN0RUz4;RRRRR
RRRRR
RRRRR--tCCMsCN0RC0ERv)qRDOCDN#RM#8RCODC0FRDoRHOVRFs)Aqv41n_.._1
.SzdRR:H5VROHEFOIC_HE80R.=R2CRoMNCs0SC
-V-RHVGRFOsRNRDD4UdU(#,RCODC0VRFRH0s#00NCFRM0CRLHRMosHCo#s0CCS8
RORzE:	RRRHV58N8s8IH0>ERR24dRMoCC0sNCR
RRRRRRORkD:	RRFbsO#C#5iBp2R
RRRRRRLRRCMoH
RRRRRRRRHRRVBR5pCi'P0CMR8NMRiBpR'=R4R'20MEC
RRRRRRRRRRRRNs_8_8ss5CoNs88I0H8ER-48MFI04FRd<2R=qR)757)Ns88I0H8ER-48MFI04FRd
2;RRRRRRRRRMRC8VRH;R
RRRRRRMRC8sRbF#OC#ORkD
	;SCRRMo8RCsMCNR0Cz	OE;R
RRzRS.:cRRsVFRHHRM8R5CEb0_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNC-
S-VRQR85N8HsI8R0E>dR42CRMC08RFsROCCN0RHIs0CCRMDNLCMRN8kRF00bkRNCMLRDC#CCDOD0RFOoH
RRRRRRRR.Sz6RR:H5VRNs88I0H8ERR>4Rd2oCCMsCN0
-S-RGVHRsVFRDONDdR4U,U(RD#CCRO0F0VRs0H#NR0CMRF0LMCHoCRso0H#C8sC
RRRRRRRRRRRRRRRR0Fk_5CMH<2R=4R''ERIC5MRs8_N8ss_CNo58I8sHE80-84RF0IMFdR42RR=HC2RDR#C';j'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RWRCIEMIR5Ns8_CNo58I8sHE80-84RF0IMFdR42RR=HC2RDR#C';j'
RRRRRRRRMSC8CRoMNCs0zCR.
6;SR--Q5VRNs88I0H8E=R<R24dRRMFI0sHCMRCNCLDRRFsFbk0kC0RMDNLCCR#D0CORoDFHMORCCC88S
RRRRRSnz.RH:RVNR58I8sHE80RR<=4Rd2oCCMsCN0
RSRRRRRRRRRRkRF0M_C5RH2<'=R4
';RRRRRRRRRRRRRRRRI_s0CHM52=R<R;W 
RRRRRRRRMSC8CRoMNCs0zCR.
n;SR--tCCMsCN0RC0ERv)qRDOCDN#RM08Rs#H-0CN0#R
RRRRRRzRS.:(RRsVFRH[RMIR5HE80_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNCR
RRRRRRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqA)v4_Ug..X7RR:DCNLD#RHR""W;R
RRRRRRRRRRRRRRCRLo
HMRRRRRRRRRRRRSqA)v4_Ug..X7RR:)Aqv41n_.._1
RSRRRRRRRRRRFRbsl0RN5bR7RQq=H>RMC_so*5.[R+48MFI0.FR*,[2R7q7)=qR>FRDIN_I858s48.RF0IMF2Rj,QR7A>R=Rj"j"q,R7A7)RR=>D_FIs8N8s.54RI8FMR0Fj
2,SRSSR RRh=qR>4R''1,R1R)q='>RjR',WR q=I>RsC0_M25H,pRBi=qR>pRBi ,Rh=AR>4R''1,R1R)A='>RjR',WR A='>RjR',BApiRR=>B,pi
SSSRRRR7Rmq=F>Rb,CMRA7m5R42=F>RkL0_k5#.H*,.[2+4,mR7A25jRR=>F_k0L.k#5RH,.2*[2R;
RRRRRRRRRRRRRFRRks0_C.o5*R[2<F=RkL0_k5#.H*,.[I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co.+*[4<2R=kRF0k_L#H.5,[.*+R42IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRMSC8CRoMNCs0zCR.
(;RRRRRMSC8CRoMNCs0zCR.
c;RRRRCRM8oCCMsCN0Rdz.;
RR
RSRR-R-RMtCC0sNCER0CqR)vCRODRD#NRM8#CCDOD0RFOoHRsVFRv)qA_4n11c_cz
S.:URRRHV5FOEH_OCI0H8ERR=co2RCsMCN
0CSR--VRHGVRFsODNDRU4dUR(,#CCDOF0RVsR0HN#00MCRFL0RCoHMRosCHC#0s
C8SzRRO:E	RRHV58N8s8IH0>ERR24.RMoCC0sNCRR
RRRRRkRRORD	:sRbF#OC#p5BiR2
RRRRRRRRLHCoMR
RRRRRRRRRH5VRB'piCMPC0MRN8pRBiRR='24'RC0EMR
RRRRRRRRRR_RsNs88_osC58N8s8IH04E-RI8FMR0F4R.2<)=Rq)7758N8s8IH04E-RI8FMR0F4;.2
RRRRRRRRCRRMH8RVR;
RRRRRCRRMb8RsCFO#k#RO;D	
RSRCRM8oCCMsCN0REzO	R;
RSRRzR.g:FRVsRRHH5MR80CbEk_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0SC
-Q-RVNR58I8sHE80R4>R.M2RCRC80OFRs0CNCsRIHR0CCLMNDNCRMF8Rkk0b0MRCNCLDRD#CCRO0DHFoOR
RRRRRRzRSd:jRRRHV58N8s8IH0>ERR24.RMoCC0sNC-
S-HRVGFRVsNROD4DRd(UU,CR#D0CORRFV0#sH0CN0R0MFRHLCMsoRC#oH0CCs8R
RRRRRRRRRRRRRRkRF0M_C5RH2<'=R4I'RERCM5Ns_8_8ss5CoNs88I0H8ER-48MFI04FR.=2RRRH2CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R ERIC5MRI_N8s5CoNs88I0H8ER-48MFI04FR.=2RRRH2CCD#R''j;R
RRRRRRCRSMo8RCsMCNR0Cz;dj
-S-RRQV58N8s8IH0<ER=.R42FRMRHIs0CCRMDNLCsRFR0FkbRk0CLMND#CRCODC0FRDoRHOM8CCCR8
SRRRRdSz4RR:H5VRNs88I0H8E=R<R24.RMoCC0sNCS
SSkSF0M_C5RH2<'=R4
';RRRRRRRRRRRRRRRRI_s0CHM52=R<R;W 
RRRRRRRRMSC8CRoMNCs0zCRd
4;SR--tCCMsCN0RC0ERv)qRDOCDN#RM08Rs#H-0CN0#R
RRRRRRzRSd:.RRsVFRH[RMIR5HE80_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNCR
RRRRRRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqA)vj_cgcnX7RR:DCNLD#RHR""W;R
RRRRRRRRRRRRRRCRLo
HMRRRRRRRRRRRRSqA)vj_cgcnX7RR:)Aqv41n_cc_1
RSRRRRRRRRRRFRbsl0RN5bR7RQq=H>RMC_so*5c[R+d8MFI0cFR*,[2R7q7)=qR>FRDIN_I858s484RF0IMF2Rj,QR7A>R=Rj"jj,j"R7q7)=AR>FRDIN_s858s484RF0IMF2Rj,S
SShS q>R=R''4,1R1)=qR>jR''W,R =qR>sRI0M_C5,H2RiBpq>R=RiBp,hR A>R=R''4,1R1)=AR>jR''W,R =AR>jR''B,RpRiA=B>Rp
i,SSSS7Rmq=F>Rb,CMRA7m5Rd2=F>RkL0_k5#cHc,R*d[+27,Rm.A52>R=R0Fk_#Lkc,5Hc+*[.R2,
SSSSA7m5R42=F>RkL0_k5#cH*,c[2+4,mR7A25jRR=>F_k0Lck#5RH,c2*[2R;
RRRRRRRRRRRRRFRRks0_Cco5*R[2<F=RkL0_k5#cH*,c[I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Coc+*[4<2R=kRF0k_L#Hc5,[c*+R42IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5[c*+R.2<F=RkL0_k5#cH*,c[2+.RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so*5c[2+dRR<=F_k0Lck#5cH,*d[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''
;
RRRRRRRRS8CMRMoCC0sNCdRz.R;
RRRRS8CMRMoCC0sNC.RzgR;
RCRRMo8RCsMCNR0Cz;.U
R
SR-RR-CRtMNCs00CRE)CRqOvRC#DDR8NMRD#CCRO0DHFoOFRVsqR)vnA4__1g1Sg
zRdd:VRHRE5OFCHO_8IH0=ERRRg2oCCMsCN0
-S-RGVHRsVFRDONDdR4U,U(RD#CCRO0F0VRs0H#NR0CMRF0LMCHoCRso0H#C8sC
RSRz	OERH:RVNR58I8sHE80R4>R4o2RCsMCN
0CRRRRRRRRk	ODRb:RsCFO#B#5p
i2RRRRRRRRRoLCHRM
RRRRRRRRRRHV5iBp'CCPMN0RMB8Rp=iRR''42ER0CRM
RRRRRRRRRsRR_8N8sC_so85N8HsI8-0E4FR8IFM0R244RR<=)7q7)85N8HsI8-0E4FR8IFM0R244;R
RRRRRRRRRCRM8H
V;RRRRRRRRCRM8bOsFCR##k	OD;R
SR8CMRMoCC0sNCORzE
	;RRRRSczdRV:RFHsRRRHM5b8C0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CSR--Q5VRNs88I0H8ERR>4R42M8CCRR0FONsC0ICRsCH0RNCMLRDCNRM8Fbk0kC0RMDNLCCR#D0CORoDFHRO
RRRRRSRRzRd6:VRHR85N8HsI8R0E>4R42CRoMNCs0SC
-V-RHVGRFOsRNRDD4UdU(#,RCODC0VRFRH0s#00NCFRM0CRLHRMosHCo#s0CCR8
RRRRRRRRRRRRRFRRkC0_M25HRR<='R4'IMECR_5sNs88_osC58N8s8IH04E-RI8FMR0F4R42=2RHR#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=WI RERCM58IN_osC58N8s8IH04E-RI8FMR0F4R42=2RHR#CDCjR''R;
RRRRRSRRCRM8oCCMsCN0R6zd;-
S-VRQR85N8HsI8R0E<4=R4M2RFsRIHR0CCLMNDFCRskRF00bkRNCMLRDC#CCDOD0RFOoHRCMC8
C8RRSRRzRSd:nRRRHV58N8s8IH0<ER=4R42CRoMNCs0SC
RRRRRRRRRRRRF_k0CHM52=R<R''4;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R R;
RRRRRSRRCRM8oCCMsCN0Rnzd;-
S-CRtMNCs00CRE)CRqOvRC#DDR8NMRH0s-N#00
C#RRRRRRRRS(zdRV:RF[sRRRHM58IH0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CRRRRRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FAVR)_qv.UjcXRU7:NRDLRCDH"#RW
";RRRRRRRRRRRRRRRRLHCoMR
RRRRRRRRRRARS)_qv.UjcXRU7:qR)vnA4__1g1Rg
RRRRRRRRRRRRRRRRRsbF0NRlb7R5Q=qR>MRH_osC5[g*+8(RF0IMF*Rg[R2,q)77q>R=RIDF_8IN84s5jFR8IFM0R,j2RA7QRR=>"jjjjjjjjR",q)77A>R=RIDF_8sN84s5jFR8IFM0R,j2
SSSSq hRR=>',4'R)11q>R=R''j, RWq>R=R0Is_5CMHR2,BqpiRR=>B,piRA hRR=>',4'R)11A>R=R''j, RWA>R=R''j,pRBi=AR>pRBi
,RSSSS7Rmq=F>Rb,CMRA7m5R(2=F>RkL0_k5#UH*,U[2+(,mR7A25nRR=>F_k0LUk#5UH,*n[+2
,RSSSS75mA6=2R>kRF0k_L#HU5,[U*+,62RA7m5Rc2=F>RkL0_k5#UH*,U[2+c,mR7A25dRR=>F_k0LUk#5UH,*d[+2
,RSSSS75mA.=2R>kRF0k_L#HU5,[U*+,.2RA7m5R42=F>RkL0_k5#UH*,U[2+4,mR7A25jRR=>F_k0LUk#5UH,*,[2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRQR7ujq52>R=R_HMs5Cog+*[UR2,7AQuRR=>",j"Ru7mq>R=RCFbM7,Rm5uAj=2R>NRbs$H0_#LkU,5H[;22
RRRRRRRRRRRRRRRR0Fk_osC5[g*2=R<R0Fk_#LkU,5HU2*[RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so*5g[2+4RR<=F_k0LUk#5UH,*4[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cgo5*.[+2=R<R0Fk_#LkU,5HU+*[.I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cog+*[d<2R=kRF0k_L#HU5,[U*+Rd2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5[g*+Rc2<F=RkL0_k5#UH*,U[2+cRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so*5g[2+6RR<=F_k0LUk#5UH,*6[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cgo5*n[+2=R<R0Fk_#LkU,5HU+*[nI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cog+*[(<2R=kRF0k_L#HU5,[U*+R(2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5[g*+RU2<b=RN0sH$k_L#HU5,R[2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRMSC8CRoMNCs0zCRd
(;RRRRRMSC8CRoMNCs0zCRd
c;RRRRCRM8oCCMsCN0Rdzd;S

RRRR-t-RCsMCNR0C0REC)RqvODCD#MRN8CR#D0CORoDFHVORF)sRq4vAn4_1U4_1Uz
Sd:URRRHV5FOEH_OCI0H8ERR=4RU2oCCMsCN0
-S-RGVHRsVFRDONDdR4U,U(RD#CCRO0F0VRs0H#NR0CMRF0LMCHoCRso0H#C8sC
RSRREzO	RR:H5VRNs88I0H8ERR>4Rj2oCCMsCN0
RRRRRRRRDkO	RR:bOsFC5##B2pi
RRRRRRRRCRLo
HMRRRRRRRRRVRHRp5BiP'CCRM0NRM8BRpi=4R''02RE
CMRRRRRRRRRRRRs8_N8ss_CNo58I8sHE80-84RF0IMFjR42=R<R7)q7N)58I8sHE80-84RF0IMFjR42R;
RRRRRRRRR8CMR;HV
RRRRRRRR8CMRFbsO#C#RDkO	S;
RCRRMo8RCsMCNR0Cz	OE;R
RRzRSd:gRRsVFRHHRM8R5CEb0_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNC-
S-VRQR85N8HsI8R0E>jR42CRMC08RFsROCCN0RHIs0CCRMDNLCMRN8kRF00bkRNCMLRDC#CCDOD0RFOoH
RRRRRRRRcSzjRR:H5VRNs88I0H8ERR>4Rj2oCCMsCN0
-S-RGVHRsVFRDONDdR4U,U(RD#CCRO0F0VRs0H#NR0CMRF0LMCHoCRso0H#C8sC
RRRRRRRRRRRRRRRR0Fk_5CMH<2R=4R''ERIC5MRs8_N8ss_CNo58I8sHE80-84RF0IMFjR42RR=HC2RDR#C';j'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RWRCIEMIR5Ns8_CNo58I8sHE80-84RF0IMFjR42RR=HC2RDR#C';j'
RRRRRRRRMSC8CRoMNCs0zCRc
j;SR--Q5VRNs88I0H8E=R<R24jRRMFI0sHCMRCNCLDRRFsFbk0kC0RMDNLCCR#D0CORoDFHMORCCC88S
RRRRRS4zcRH:RVNR58I8sHE80RR<=4Rj2oCCMsCN0
RSRRRRRRRRRRkRF0M_C5RH2<'=R4
';RRRRRRRRRRRRRRRRI_s0CHM52=R<R;W 
RRRRRRRRMSC8CRoMNCs0zCRc
4;SR--tCCMsCN0RC0ERv)qRDOCDN#RM08Rs#H-0CN0#R
RRRRRRzRSc:.RRsVFRH[RMIR5HE80_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNCR
RRRRRRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqA)vj_4.4cXn:7RRLDNCHDR#WR""R;
RRRRRRRRRRRRRLRRCMoH
RRRRRRRRRRRR)SAq4v_jX.c4Rn7:qR)vnA4_U14_U14
RRRRRRRRRRRRRRRRbRRFRs0lRNb5q7QRR=>HsM_C4o5U+*[486RF0IMFUR4*,[2R7q7)=qR>FRDIN_I858sgFR8IFM0R,j2RA7QRR=>"jjjjjjjjjjjjjjjjR",q)77A>R=RIDF_8sN8gs5RI8FMR0Fj
2,SSSS Rhq='>R4R',1q1)RR=>',j'RqW RR=>I_s0CHM52B,RpRiq=B>RpRi, RhA='>R4R',1A1)RR=>',j'RAW RR=>',j'RiBpA>R=RiBp,SR
S7SSm=qR>bRFCRM,75mA4R62=F>RkL0_kn#454H,n+*[4,62RA7m524cRR=>F_k0L4k#n,5H4[n*+24c,SR
S7SSm4A5d=2R>kRF0k_L#54nHn,4*4[+dR2,75mA4R.2=F>RkL0_kn#454H,n+*[4,.2RA7m5244RR=>F_k0L4k#n,5H4[n*+244,SR
S7SSm4A5j=2R>kRF0k_L#54nHn,4*4[+jR2,75mAg=2R>kRF0k_L#54nHn,4*g[+27,RmUA52>R=R0Fk_#Lk4Hn5,*4n[2+U,SR
S7SSm(A52>R=R0Fk_#Lk4Hn5,*4n[2+(,mR7A25nRR=>F_k0L4k#n,5H4[n*+,n2RA7m5R62=F>RkL0_kn#454H,n+*[6R2,
SSSSA7m5Rc2=F>RkL0_kn#454H,n+*[cR2,75mAd=2R>kRF0k_L#54nHn,4*d[+27,Rm.A52>R=R0Fk_#Lk4Hn5,*4n[2+.,SR
S7SSm4A52>R=R0Fk_#Lk4Hn5,*4n[2+4,mR7A25jRR=>F_k0L4k#n,5H4[n*2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRR7qQuRR=>HsM_C4o5U+*[48(RF0IMFUR4*4[+nR2,7AQuRR=>""jj,mR7u=qR>bRFC
M,RRRRRRRRRRRRRRRRRRRRRRRRRRRR7Amu5R42=b>RN0sH$k_L#54nH*,.[2+4,mR7ujA52>R=RsbNH_0$L4k#n,5H.2*[2R;
RRRRRRRRRRRRRFRRks0_C4o5U2*[RR<=F_k0L4k#n,5H4[n*2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[4<2R=kRF0k_L#54nHn,4*4[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[.<2R=kRF0k_L#54nHn,4*.[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[d<2R=kRF0k_L#54nHn,4*d[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[c<2R=kRF0k_L#54nHn,4*c[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[6<2R=kRF0k_L#54nHn,4*6[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[n<2R=kRF0k_L#54nHn,4*n[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[(<2R=kRF0k_L#54nHn,4*([+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[U<2R=kRF0k_L#54nHn,4*U[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[g<2R=kRF0k_L#54nHn,4*g[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[4Rj2<F=RkL0_kn#454H,n+*[4Rj2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[4+42=R<R0Fk_#Lk4Hn5,*4n[4+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[4R.2<F=RkL0_kn#454H,n+*[4R.2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[d+42=R<R0Fk_#Lk4Hn5,*4n[d+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[4Rc2<F=RkL0_kn#454H,n+*[4Rc2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[6+42=R<R0Fk_#Lk4Hn5,*4n[6+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[4Rn2<b=RN0sH$k_L#54nH*,.[I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+24(RR<=bHNs0L$_kn#45.H,*4[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRSRRCRM8oCCMsCN0R.zc;R
RRSRRCRM8oCCMsCN0Rgzd;R
RRMRC8CRoMNCs0zCRd
U;
RSRR-R-RMtCC0sNCER0CqR)vCRODRD#NRM8#CCDOD0RFOoHRsVFRv)qA_4n1_dn1
dnSUzdNRR:H5VROHEFOIC_HE80Rd=Rno2RCsMCN
0CSR--VRHGVRFsODNDRU4dUR(,#CCDOF0RVsR0HN#00MCRFL0RCoHMRosCHC#0s
C8SRRRz	OERH:RVNR58I8sHE80Rg>R2CRoMNCs0SC
RRRRk	ODRb:RsCFO#B#5p
i2SLSRCMoH
RSSRRHV5iBp'CCPMN0RMB8Rp=iRR''42ER0CSM
SRRRRNs_8_8ss5CoNs88I0H8ER-48MFI0gFR2=R<R7)q7N)58I8sHE80-84RF0IMF2Rg;S
SRMRC8VRH;S
SCRM8bOsFCR##k	OD;R
SRMRC8CRoMNCs0zCRO;E	
RSRRdRzg:NRRsVFRHHRM8R5CEb0_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNC-
S-VRQR85N8HsI8R0E>2RgRCMC8FR0RCOsNR0CI0sHCMRCNCLDR8NMR0FkbRk0CLMND#CRCODC0FRDo
HOSzSScRjN:VRHR85N8HsI8R0E>2RgRMoCC0sNC-
S-HRVGFRVsNROD4DRd(UU,CR#D0CORRFV0#sH0CN0R0MFRHLCMsoRC#oH0CCs8S
SSkSF0M_C5RH2<'=R4I'RERCM5Ns_8_8ss5CoNs88I0H8ER-48MFI0gFR2RR=HC2RDR#C';j'
SSSS0Is_5CMH<2R= RWRCIEMIR5Ns8_CNo58I8sHE80-84RF0IMF2RgRH=R2DRC#'CRj
';SCSSMo8RCsMCNR0CzNcj;-
S-VRQR85N8HsI8R0E<g=R2FRMRHIs0CCRMDNLCsRFR0FkbRk0CLMND#CRCODC0FRDoRHOM8CCCS8
ScSz4:NRRRHV58N8s8IH0<ER=2RgRMoCC0sNCS
SSkSF0M_C5RH2<'=R4
';SSSSI_s0CHM52=R<R;W 
SSSCRM8oCCMsCN0R4zcNS;
-t-RCsMCNR0C0REC)RqvODCD#MRN8sR0H0-#N#0C
SSSzNc.RV:RF[sRRRHM58IH0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CRRRRRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FAVR)_qv6X4.dR.7:NRDLRCDH"#RW
";RRRRRRRRRRRRRRRRLHCoMS
SS)SAq6v_4d.X.:7RRv)qA_4n1_dn1
dnRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRFRbsl0RN5bR7RQq=H>RMC_son5d*d[+4FR8IFM0R*dn[R2,q)77q>R=RIDF_8IN8Us5RI8FMR0FjR2,7RQA=">Rjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"q,R7A7)RR=>D_FIs8N8sR5U8MFI0jFR2S,
S SSh=qR>4R''1,R1R)q='>RjR',WR q=I>RsC0_M25H,pRBi=qR>pRBi ,Rh=AR>4R''1,R1R)A='>RjR',WR A='>RjR',BApiRR=>B,pi
SSSSq7mRR=>FMbC,mR7A45d2>R=R0Fk_#LkdH.5,*d.[4+d27,RmdA5j=2R>kRF0k_L#5d.H.,d*d[+j
2,SSSS75mA.Rg2=F>RkL0_k.#d5dH,.+*[.,g2RA7m52.URR=>F_k0Ldk#.,5Hd[.*+2.U,mR7A(5.2>R=R0Fk_#LkdH.5,*d.[(+.2S,
S7SSm.A5n=2R>kRF0k_L#5d.H.,d*.[+nR2,75mA.R62=F>RkL0_k.#d5dH,.+*[.,62RA7m52.cRR=>F_k0Ldk#.,5Hd[.*+2.c,S
SSmS7Ad5.2>R=R0Fk_#LkdH.5,*d.[d+.27,Rm.A5.=2R>kRF0k_L#5d.H.,d*.[+.R2,75mA.R42=F>RkL0_k.#d5dH,.+*[.,42
SSSSA7m52.jRR=>F_k0Ldk#.,5Hd[.*+2.j,mR7Ag542>R=R0Fk_#LkdH.5,*d.[g+427,Rm4A5U=2R>kRF0k_L#5d.H.,d*4[+U
2,SSSS75mA4R(2=F>RkL0_k.#d5dH,.+*[4,(2RA7m524nRR=>F_k0Ldk#.,5Hd[.*+24n,mR7A6542>R=R0Fk_#LkdH.5,*d.[6+42S,
S7SSm4A5c=2R>kRF0k_L#5d.H.,d*4[+cR2,75mA4Rd2=F>RkL0_k.#d5dH,.+*[4,d2RA7m524.RR=>F_k0Ldk#.,5Hd[.*+24.,S
SSmS7A4542>R=R0Fk_#LkdH.5,*d.[4+427,Rm4A5j=2R>kRF0k_L#5d.H.,d*4[+jR2,75mAg=2R>kRF0k_L#5d.H.,d*g[+2S,
S7SSmUA52>R=R0Fk_#LkdH.5,*d.[2+U,mR7A25(RR=>F_k0Ldk#.,5Hd[.*+,(2RA7m5Rn2=F>RkL0_k.#d5dH,.+*[n
2,SSSS75mA6=2R>kRF0k_L#5d.H.,d*6[+27,RmcA52>R=R0Fk_#LkdH.5,*d.[2+c,mR7A25dRR=>F_k0Ldk#.,5Hd[.*+,d2
SSSSA7m5R.2=F>RkL0_k.#d5dH,.+*[.R2,75mA4=2R>kRF0k_L#5d.H.,d*4[+27,RmjA52>R=R0Fk_#LkdH.5,*d.[
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR7qQuRR=>HsM_Cdo5n+*[d86RF0IMFnRd*d[+.R2,7AQuRR=>"jjjjR",7qmuRR=>FMbC,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7udA52>R=RsbNH_0$Ldk#.,5Hc+*[dR2,7Amu5R.2=b>RN0sH$k_L#5d.H*,c[2+.,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7u4A52>R=RsbNH_0$Ldk#.,5Hc+*[4R2,7Amu5Rj2=b>RN0sH$k_L#5d.H*,c[;22
SSSS0Fk_osC5*dn[<2R=kRF0k_L#5d.H.,d*R[2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
SSSS0Fk_osC5*dn[2+4RR<=F_k0Ldk#.,5Hd[.*+R42IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
SSSS0Fk_osC5*dn[2+.RR<=F_k0Ldk#.,5Hd[.*+R.2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
SSSS0Fk_osC5*dn[2+dRR<=F_k0Ldk#.,5Hd[.*+Rd2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
SSSS0Fk_osC5*dn[2+cRR<=F_k0Ldk#.,5Hd[.*+Rc2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
SSSS0Fk_osC5*dn[2+6RR<=F_k0Ldk#.,5Hd[.*+R62IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
SSSS0Fk_osC5*dn[2+nRR<=F_k0Ldk#.,5Hd[.*+Rn2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
SSSS0Fk_osC5*dn[2+(RR<=F_k0Ldk#.,5Hd[.*+R(2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
SSSS0Fk_osC5*dn[2+URR<=F_k0Ldk#.,5Hd[.*+RU2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
SSSS0Fk_osC5*dn[2+gRR<=F_k0Ldk#.,5Hd[.*+Rg2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
SSSS0Fk_osC5*dn[j+42=R<R0Fk_#LkdH.5,*d.[j+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''S;
SFSSks0_Cdo5n+*[4R42<F=RkL0_k.#d5dH,.+*[4R42IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
SSSS0Fk_osC5*dn[.+42=R<R0Fk_#LkdH.5,*d.[.+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''S;
SFSSks0_Cdo5n+*[4Rd2<F=RkL0_k.#d5dH,.+*[4Rd2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
SSSS0Fk_osC5*dn[c+42=R<R0Fk_#LkdH.5,*d.[c+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''S;
SFSSks0_Cdo5n+*[4R62<F=RkL0_k.#d5dH,.+*[4R62IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
SSSS0Fk_osC5*dn[n+42=R<R0Fk_#LkdH.5,*d.[n+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''S;
SFSSks0_Cdo5n+*[4R(2<F=RkL0_k.#d5dH,.+*[4R(2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
SSSS0Fk_osC5*dn[U+42=R<R0Fk_#LkdH.5,*d.[U+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''S;
SFSSks0_Cdo5n+*[4Rg2<F=RkL0_k.#d5dH,.+*[4Rg2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
SSSS0Fk_osC5*dn[j+.2=R<R0Fk_#LkdH.5,*d.[j+.2ERIC5MRF_k0CHM52RR='24'R#CDCZR''S;
SFSSks0_Cdo5n+*[.R42<F=RkL0_k.#d5dH,.+*[.R42IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
SSSS0Fk_osC5*dn[.+.2=R<R0Fk_#LkdH.5,*d.[.+.2ERIC5MRF_k0CHM52RR='24'R#CDCZR''S;
SFSSks0_Cdo5n+*[.Rd2<F=RkL0_k.#d5dH,.+*[.Rd2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
SSSS0Fk_osC5*dn[c+.2=R<R0Fk_#LkdH.5,*d.[c+.2ERIC5MRF_k0CHM52RR='24'R#CDCZR''S;
SFSSks0_Cdo5n+*[.R62<F=RkL0_k.#d5dH,.+*[.R62IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
SSSS0Fk_osC5*dn[n+.2=R<R0Fk_#LkdH.5,*d.[n+.2ERIC5MRF_k0CHM52RR='24'R#CDCZR''S;
SFSSks0_Cdo5n+*[.R(2<F=RkL0_k.#d5dH,.+*[.R(2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
SSSS0Fk_osC5*dn[U+.2=R<R0Fk_#LkdH.5,*d.[U+.2ERIC5MRF_k0CHM52RR='24'R#CDCZR''S;
SFSSks0_Cdo5n+*[.Rg2<F=RkL0_k.#d5dH,.+*[.Rg2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
SSSS0Fk_osC5*dn[j+d2=R<R0Fk_#LkdH.5,*d.[j+d2ERIC5MRF_k0CHM52RR='24'R#CDCZR''S;
SFSSks0_Cdo5n+*[dR42<F=RkL0_k.#d5dH,.+*[dR42IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
SSSS0Fk_osC5*dn[.+d2=R<RsbNH_0$Ldk#.,5Hc2*[RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;S
SSkSF0C_son5d*d[+d<2R=NRbs$H0_#LkdH.5,[c*+R42IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
SSSS0Fk_osC5*dn[c+d2=R<RsbNH_0$Ldk#.,5Hc+*[.I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';SSSSF_k0s5Cod[n*+2d6RR<=bHNs0L$_k.#d5cH,*d[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''S;
SMSC8CRoMNCs0zCRc;.N
CSSMo8RCsMCNR0CzNdg;C
SMo8RCsMCNR0CzNdU;R
RCRM8oCCMsCN0Rdzc;R

RczcRH:RVMR5Fs0RNs88_osC2CRoMNCs0-CR-CRoMNCs0#CRCODC0NRslR
RR-R-RRQVNs88I0H8ERR<6#RN#MHoR''jRR0Fk#MkCL8RH
0#RRRRzRjR:VRHR85N8HsI8R0E=2R4RMoCC0sNCR
RRRRRRFRDIN_s8_8s#=R<Rj"jj"jjRs&RNs8_C#o_5;j2
RRRRRRRRIDF_8IN8#s_RR<="jjjjRj"&NRI8C_so5_#j
2;RRRRCRM8oCCMsCN0R;zj
RRRRRz4RH:RVNR58I8sHE80R.=R2CRoMNCs0RC
RRRRRDRRFsI_Ns88_<#R=jR"j"jjRs&RNs8_C#o_584RF0IMF2Rj;R
RRRRRRFRDIN_I8_8s#=R<Rj"jjRj"&NRI8C_so5_#4FR8IFM0R;j2
RRRR8CMRMoCC0sNC4Rz;R
RR.RzRRR:H5VRNs88I0H8ERR=do2RCsMCN
0CRRRRRRRRD_FIs8N8sR_#<"=Rj"jjRs&RNs8_C#o_58.RF0IMF2Rj;R
RRRRRRFRDIN_I8_8s#=R<Rj"jj&"RR8IN_osC_.#5RI8FMR0Fj
2;RRRRCRM8oCCMsCN0R;z.
RRRRRzdRH:RVNR58I8sHE80Rc=R2CRoMNCs0RC
RRRRRDRRFsI_Ns88_<#R=jR"j&"RR8sN_osC_d#5RI8FMR0Fj
2;RRRRRRRRD_FII8N8sR_#<"=RjRj"&NRI8C_so5_#dFR8IFM0R;j2
RRRR8CMRMoCC0sNCdRz;z
ScRS:H5VRNs88I0H8ERR=6o2RCsMCN
0CSFSDIN_s8_8s#=R<R''jRs&RNs8_C#o_58cRF0IMF2Rj;S
SD_FII8N8sR_#<'=Rj&'RR8IN_osC_c#5RI8FMR0Fj
2;S8CMRMoCC0sNCcRz;R
RR6RzRRR:H5VRNs88I0H8ERR>6o2RCsMCN
0CRRRRRRRRD_FIs8N8sR_#<s=RNs8_C#o_586RF0IMF2Rj;R
RRRRRRFRDIN_I8_8s#=R<R8IN_osC_6#5RI8FMR0Fj
2;RRRRCRM8oCCMsCN0R;z6
R
RR-R-RRQV5M8H_osC2CRso0H#C7sRQkhR#oHMRiBp
RRRRRznRH:RV8R5HsM_CRo2oCCMsCN0
RRRRRRRRFbsO#C#Rp5Bi7,RQRh2LHCoMR
RRRRRRRRRRVRHRp5BiRR='R4'NRM8B'piCMPC002RE
CMRRRRRRRRRRRRRRRRHsM_C#o_RR<=7;Qh
RRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMRFbsO#C#;R
RRMRC8CRoMNCs0zCRnR;
RzRR(:RRRRHV50MFRM8H_osC2CRoMNCs0RC
RRRRRRRRRHRRMC_soR_#<7=RQ
h;RRRRCRM8oCCMsCN0R;z(
R
RR-R-RRQV5k8F0C_sos2RC#oH0RCs7amzRHk#MmoRB
piRRRRzRUR:VRHRF58ks0_CRo2oCCMsCN0
RRRRRRRRFbsO#C#RB5mpRi,F_k0s_Co#L2RCMoH
RRRRRRRRRRRRRHV5pmBiRR='R4'NRM8miBp'CCPMR020MEC
RRRRRRRRRRRRRRRRz7ma=R<R0Fk_osC_
#;RRRRRRRRRRRRCRM8H
V;RRRRRRRRCRM8bOsFC;##
RRRR8CMRMoCC0sNCURz;R
RRgRzRRR:H5VRMRF080Fk_osC2CRoMNCs0RC
RRRRRRRRR7RRmRza<F=Rks0_C#o_;R
RRMRC8CRoMNCs0zCRg
;
RRRR-Q-RVNR58_8ss2CoRosCHC#0s7Rq7k)R#oHMRiBp
RRRRjz4RRR:H5VRs8N8sC_soo2RCsMCN
0CRRRRRRRRbOsFCR##5iBp,qR)727)RoLCHRM
RRRRRRRRRHRRVBR5p=iRR''4R8NMRiBp'CCPMR020MEC
RRRRRRRRRRRRRRRR8sN_osC_<#R=qR)757)Ns88I0H8ER-48MFI0jFR2R;
RRRRRRRRRCRRMH8RVR;
RRRRRCRRMb8RsCFO#
#;RRRRCRM8oCCMsCN0Rjz4;R
RR4Rz4RR:H5VRMRF0s8N8sC_soo2RCsMCN
0CRRRRRRRRRRRRs_N8s_Co#=R<R7)q7
);RRRRCRM8oCCMsCN0R4z4;R

R-RR-VRQR85N8ss_CRo2sHCo#s0CR7q7)#RkHRMoB
piRRRRzR4.RH:RVIR5Ns88_osC2CRoMNCs0RC
RRRRRbRRsCFO#5#RB,piR7Wq7R)2LHCoMR
RRRRRRRRRRVRHRp5BiRR='R4'NRM8B'piCMPC002RE
CMRRRRRRRRRRRRRRRRI_N8s_Co#=R<R7Wq7N)58I8sHE80-84RF0IMF2Rj;R
RRRRRRRRRRMRC8VRH;R
RRRRRRMRC8sRbF#OC#R;
RCRRMo8RCsMCNR0Cz;4.
RRRRdz4RH:RVMR5FI0RNs88_osC2CRoMNCs0RC
RRRRRRRRRIRRNs8_C#o_RR<=W7q7)R;
RCRRMo8RCsMCNR0Cz;4d
RRRRRRRRR
RR-R-RMtCC0sNCER0CqR)vCRODRD#NRM8#CCDOD0RFOoH
RRRRcz4RV:RFHsRRRHM5lMk_DOCDc_nR4-R2FR8IFM0RojRCsMCN
0CRRRR-Q-RVNR58I8sHE80R6>R2CRMC08RFsROCCN0RHIs0CCRMDNLCMRN8kRF00bkRNCMLRDC#CCDOD0RFOoH
RRRRRRRR6z4RH:RVNR58I8sHE80Rn>R2CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_M5_#H<2R=4R''ERIC5MRs_N8s_Co#85N8HsI8-0E4FR8IFM0RRn2=2RHR#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_M5_#H<2R= RWRCIEMIR5Ns8_C#o_58N8s8IH04E-RI8FMR0Fn=2RRRH2CCD#R''j;R
RRRRRRMRC8CRoMNCs0zCR4
6;RRRR-Q-RVNR58I8sHE80RR<=6M2RFsRIHR0CCLMNDFCRskRF00bkRNCMLRDC#CCDOD0RFOoHRCMC8
C8RRRRRRRRzR4n:VRHR85N8HsI8R0E<n=R2CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_M5_#H<2R=4R''R;
RRRRRRRRRRRRRIRRsC0_M5_#H<2R= RW;R
RRRRRRMRC8CRoMNCs0zCR4
n;RRRR-t-RCsMCNR0C0REC)RqvODCD#MRN8sR0H0-#N#0C
RRRRRRRR(z4RV:RF[sRRRHM58IH0-ERRR428MFI0jFRRMoCC0sNCR
RRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqz)vRnc:NRDLRCDH"#R1"7aRH&RMo0CCHs'lCNo58IH0RE2&7R""RR&HCM0o'CsHolNC*5HnRc2&WR""RR&HCM0o'CsHolNC25[R"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05+5H4n2*c8,RCEb02&2RR""XRH&RMo0CCHs'lCNo54[+2R;
RRRRRRRRRLRRCMoH
RRRRRRRRRRRRqz)vRnc:)RXqcvnXR47
RRRRRRRRRRRRRRRRsbF0NRlb7R5RR=>HsM_C#o_5,[2RRqj=D>RFII_Ns88_j#52q,R4>R=RIDF_8IN8#s_5,42RRq.=D>RFII_Ns88_.#52R,
RRRRRRRRRRRRRRRRRRRRRRRRRRqd=D>RFII_Ns88_d#52q,Rc>R=RIDF_8IN8#s_5,c2RRq6=D>RFII_Ns88_6#52
,RSSSSSRSR7qu)j>R=RIDF_8sN8#s_5,j2R)7uq=4R>FRDIN_s8_8s#254,uR7)Rq.=D>RFsI_Ns88_.#52S,
SSSSS7RRud)qRR=>D_FIs8N8s5_#dR2,7qu)c>R=RIDF_8sN8#s_5,c2R)7uq=6R>FRDIN_s8_8s#256,SR
SSSSSWRR >R=R0Is__CM#25H,BRWp=iR>pRBi7,Ru=mR>kRF0k_L#c_n#,5H[;22
RRRRRRRRRRRRRRRR0Fk_osC_[#52=R<R0Fk_#Lk_#nc5[H,2ERIC5MRF_k0C#M_5RH2=4R''C2RDR#C';Z'
RRRRRRRR8CMRMoCC0sNC4Rz(R;
RRRRCRM8oCCMsCN0Rcz4;RRRRRRRRRRRRR
RRRRR
RRRRR--tCCMsCN0RdNR.FRIs88RCRCb)RqvODCDRRHVNsbbFHbsNR0CRRRRRRRRRRRRRRR
RzRR4:URRRHV5lMk_DOCD._dR4=R2CRoMNCs0RC
R-RR-VRQR85N8HsI8R0E>2R(RCMC8FR0RCOsNR0CI0sHCMRCNCLDR8NMR0FkbRk0CLMND#CRCODC0FRDo
HORRRRRRRRzN4gRH:RVNR58I8sHE80Rn>R2CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_M._dRR<='R4'IMECRs55Ns8_C#o_58N8s8IH04E-RI8FMR0Fn=2RRlMk_DOCDc_n2MRN8sR5Ns8_C#o_5R62=jR''R22CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C_Rd.<W=R ERIC5MR58IN_osC_N#58I8sHE80-84RF0IMF2RnRM=RkOl_C_DDnRc2NRM858IN_osC_6#52RR='2j'2DRC#'CRj
';RRRRRRRRCRM8oCCMsCN0Rgz4NR;
RRRRRzRR4RgL:VRHR85N8HsI8R0E=RRnNRM8M_klODCD_Rnc=2RjRMoCC0sNCR
RRRRRRRRRRRRRRkRF0M_C_Rd.<'=R4I'RERCM5N5s8C_so5_#6=2RR''j2C2RDR#C';j'
RRRRRRRRRRRRRRRR0Is__CMd<.R= RWRCIEM5R5I_N8s_Co#256R'=Rj2'2R#CDCjR''R;
RRRRRCRRMo8RCsMCNR0CzL4g;RRRRR--Q5VRNs88I0H8E=R<RR62MIFRsCH0RNCMLRDCFFsRkk0b0MRCNCLDRD#CCRO0DHFoOCRMC88C
RRRRRRRRjz.RH:RVNR58I8sHE80RR<=6o2RCsMCN
0CRRRRRRRRRRRRRRRRF_k0CdM_.=R<R''4;R
RRRRRRRRRRRRRRsRI0M_C_Rd.<W=R R;
RRRRRCRRMo8RCsMCNR0Cz;.j
RRRRR--tCCMsCN0RC0ERv)qRDOCDMRN8sR0H0-#N
0CRRRRRRRRzR.4:FRVsRR[H5MRI0H8ERR-482RF0IMFRRjoCCMsCN0
RRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVzv)qd:.RRLDNCHDR#1R"7Ra"&MRH0CCosl'HN5oCI0H8E&2RR""7RH&RMo0CCHs'lCNo5lMk_DOCDc_n*2ncR"&RW&"RR0HMCsoC'NHlo[C52RR&"R "&MRH0CCosl'HN5oCo_C0C_M880CbEk5MlC_ODnD_cc*nRd+R.8,RCEb02&2RR""XRH&RMo0CCHs'lCNo54[+2R;
RRRRRRRRRLRRCMoH
RRRRRRRRRRRRqz)vRd.:)RXq.vdXR47
RRRRRRRRRRRRRRRRsbF0NRlb7R5RR=>HsM_C#o_5,[2RRqj=D>RFII_Ns88_j#52q,R4>R=RIDF_8IN8#s_5,42RRq.=D>RFII_Ns88_.#52R,
RRRRRRRRRRRRRRRRRRRRRRRRRRqd=D>RFII_Ns88_d#52q,Rc>R=RIDF_8IN8#s_5,c2RS
SSSSSRuR7)Rqj=D>RFsI_Ns88_j#527,Ru4)qRR=>D_FIs8N8s5_#4R2,7qu).>R=RIDF_8sN8#s_5,.2
SSSSRSSR)7uq=dR>FRDIN_s8_8s#25d,uR7)Rqc=D>RFsI_Ns88_c#52
,RSSSSSRSRW= R>sRI0M_C_,d.RpWBi>R=RiBp,uR7m>R=R0Fk_#Lk_#d.5lMk_DOCD._d,2[2;R
RRRRRRRRRRRRRRkRF0C_so5_#[<2R=kRF0k_L#._d#k5MlC_ODdD_.2,[RCIEMFR5kC0_M._dR'=R4R'2CCD#R''Z;R
RRRRRRCRRMo8RCsMCNR0Cz;.4
RRRRMRC8CRoMNCs0zCR4RU;RRRRRRRRRR

R-RR-CRtMNCs0NCRRR4nI8FsRC8CbqR)vCRODHDRVbRNbbsFs0HNCRRRRRRRRRRRRRRR
RRRR.z.RH:RVMR5kOl_C_DD4=nRRR42oCCMsCN0
RRRRR--Q5VRNs88I0H8ERR>6M2RCRC80OFRs0CNCsRIHR0CCLMNDNCRMF8Rkk0b0MRCNCLDRD#CCRO0DHFoOR
RRRRRR.Rzd:NRRRHV58N8s8IH0>ERRNnRMM8RkOl_C_DDd=.RRR42oCCMsCN0
RRRRRRRRRRRRRRRR0Fk__CM4<nR=4R''ERIC5MR58sN_osC_N#58I8sHE80-84RF0IMF2RnRM=RkOl_C_DDnRc2NRM858sN_osC_6#52RR='24'R8NMRN5s8C_so5_#c=2RR''j2C2RDR#C';j'
RRRRRRRRRRRRRRRR0Is__CM4<nR= RWRCIEM5R5I_N8s_Co#85N8HsI8-0E4FR8IFM0RRn2=kRMlC_ODnD_cN2RM58RI_N8s_Co#256R'=R4R'2NRM858IN_osC_c#52RR='2j'2DRC#'CRj
';RRRRRRRRCRM8oCCMsCN0Rdz.NR;
RRRRRzRR.RdL:VRHR85N8HsI8R0E>RRnNRM8M_klODCD_Rd./4=R2CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_Mn_4RR<='R4'IMECRs55Ns8_C#o_58N8s8IH04E-RI8FMR0Fn=2RRlMk_DOCDc_n2MRN8sR5Ns8_C#o_5R62=jR''N2RM58Rs_N8s_Co#25cR'=Rj2'2R#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_Mn_4RR<=WI RERCM5N5I8C_so5_#Ns88I0H8ER-48MFI0nFR2RR=M_klODCD_2ncR8NMRN5I8C_so5_#6=2RR''j2MRN8IR5Ns8_C#o_5Rc2=jR''R22CCD#R''j;R
RRRRRRMRC8CRoMNCs0zCR.;dL
RRRRRRRRdz.ORR:H5VRNs88I0H8ERR=nMRN8kRMlC_ODdD_.RR=4o2RCsMCN
0CRRRRRRRRRRRRRRRRF_k0C4M_n=R<R''4RCIEM5R5s_N8s_Co#256R'=R4R'2NRM858sN_osC_c#52RR='2j'2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0C4M_n=R<RRW IMECRI55Ns8_C#o_5R62=4R''N2RM58RI_N8s_Co#25cR'=Rj2'2R#CDCjR''R;
RRRRRCRRMo8RCsMCNR0CzO.d;R
RRRRRR.Rzd:8RRRHV58N8s8IH0=ERRN6RMM8RkOl_C_DDd/.R=2R4RMoCC0sNCR
RRRRRRRRRRRRRRkRF0M_C_R4n<'=R4I'RERCM5N5s8C_so5_#Ns88I0H8ER-48MFI0cFR2RR=M_klODCD_2d.2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0C4M_n=R<RRW IMECRI55Ns8_C#o_58N8s8IH04E-RI8FMR0Fc=2RRlMk_DOCD._d2C2RDR#C';j'
RRRRRRRR8CMRMoCC0sNC.RzdR8;R-RR-VRQR85N8HsI8R0E<6=R2FRMRHIs0CCRMDNLCsRFR0FkbRk0CLMND#CRCODC0FRDoRHOM8CCCR8
RRRRRzRR.:cRRRHV58N8s8IH0<ER=2RcRMoCC0sNCR
RRRRRRRRRRRRRRkRF0M_C_R4n<'=R4
';RRRRRRRRRRRRRRRRI_s0C4M_n=R<R;W 
RRRRRRRR8CMRMoCC0sNC.RzcR;
R-RR-CRtMNCs00CRE)CRqOvRCRDDNRM80-sH#00NCR
RRRRRR.Rz6RR:VRFs[MRHRH5I8R0E-2R4RI8FMR0FjCRoMNCs0RC
RRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)Rzqnv4RD:RNDLCRRH#"a17"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloMC5kOl_C_DDnnc*cRR+M_klODCD_*d.dR.2&WR""RR&HCM0o'CsHolNC25[R"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05lMk_DOCDc_n*Rnc+kRMlC_ODdD_..*dR4+Rn8,RCEb02&2RR""XRH&RMo0CCHs'lCNo54[+2R;
RRRRRRRRRLRRCMoH
RRRRRRRRRRRRqz)vR4n:qR)vX4n4
7RRRRRRRRRRRRRRRRRb0FsRblNRR57=H>RMC_so5_#[R2,q=jR>FRDIN_I8_8s#25j,4RqRR=>D_FII8N8s5_#4R2,q=.R>FRDIN_I8_8s#25.,R
RRRRRRRRRRRRRRRRRRRRRRRRRq=dR>FRDIN_I8_8s#25d,uR7)Rqj=D>RFsI_Ns88_j#527,Ru4)qRR=>D_FIs8N8s5_#4R2,7qu).>R=RIDF_8sN8#s_5,.2
SSSSRSSR)7uq=dR>FRDIN_s8_8s#25d, RWRR=>I_s0C4M_nW,RBRpi=B>RpRi,7Rum=F>RkL0_k4#_nM#5kOl_C_DD4[n,2
2;RRRRRRRRRRRRRRRRF_k0s_Co#25[RR<=F_k0L_k#45n#M_klODCD_,4n[I2RERCM50Fk__CM4=nRR''42DRC#'CRZ
';RRRRRRRRCRM8oCCMsCN0R6z.;R
RRMRC8CRoMNCs0zCR.R.;R
RRRMRC8CRoMNCs0zCRc
c;CRM8NEsOHO0C0CksR_MFsOI_E	CO;-

--
-R#pN0lRHblDCCNM00MHFRRH#8NCVk
D0-N-
sHOE00COkRsC#CCDOs0_NFlRVqR)v__)W#RH
MVkOF0HMCRo0M_C8C_8b50E#CHxRH:RMo0CC;sRRb8C0:ERR0HMCsoC2CRs0MksR0HMCsoCR
H#PHNsNCLDRMlH_x#HCRR:HCM0oRCs:j=R;C
Lo
HMRHRlMH_#x:CR=CR8b;0E
HRRV#R5HRxC<CR8b20ERC0EMR
RRHRlMH_#x:CR=HR#x
C;RMRC8VRH;R
RskC0slMRH#M_H;xC
8CMR0oC_8CM_b8C0
E;O#FM00NMRlMk_DOCD:#RR0HMCsoCRR:=5C58bR0E-2R4/24n;RRRRRRRRRRRRR--yVRFRv)q44nX7CRODRD#M8CCC08
$RbCF_k0L_k#0C$bRRH#NNss$MR5kOl_C#DDRI8FMR0FjI,RHE80-84RF0IMF2RjRRFV#_08DHFoO#;
HNoMDkRF0k_L#RR:F_k0L_k#0C$b;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$F8VRFRk05bHMk00RFsR0H0-#N#0C2H
#oDMNR0Fk_RCM:0R#8F_Do_HOP0COFMs5kOl_C#DDRI8FMR0FjR2;RRRRR-RR-MRCNCLD#FRVssR0H0-#N#0C
o#HMRNDI_s0C:MRR8#0_oDFHPO_CFO0sk5MlC_ODRD#8MFI0jFR2R;RRRRRR-R-RHIs0CCRMDNLCV#RFCsRNROEsRFIF)VRqOvRC#DD
o#HMRNDHsM_C:oRR8#0_oDFHPO_CFO0sH5I8-0E4FR8IFM0R;j2RRRRRRRRR-R-RCk#8FR0RosCHC#0sQR7h#R
HNoMDkRF0C_soRR:#_08DHFoOC_POs0F58IH04E-RI8FMR0FjR2;RRRRRRRR-k-R#RC80sFRC#oH0RCs7amz
o#HMRNDs_N8sRCo:0R#8F_Do_HOP0COFNs58I8sHE80-84RF0IMF2Rj;RRRR-R-RCk#8FR0RosCHC#0sqR)7
7)#MHoNIDRNs8_C:oRR8#0_oDFHPO_CFO0s85N8HsI8-0E4FR8IFM0R;j2RRRRRR--k8#CRR0FsHCo#s0CR7Wq7#)
HNoMDFRDIN_s8R8s:0R#8F_Do_HOP0COFds5RI8FMR0FjR2;RRRRRRRRRRRR-s-RNs88R0LH#MRHbRk00)FRqOvRC#DDRR5cL#H0RJsCkCHs8#2
HNoMDFRDIN_I8R8s:0R#8F_Do_HOP0COFds5RI8FMR0FjR2;RRRRRRRRRRRR-I-RNs88R0LH#MRHbRk00)FRqOvRC#DDRR5cL#H0RJsCkCHs8N2
0H0sLCk0Rs\3NFl_VCV#0:\RRs#0H;Mo
C
Lo
HM
RRRRR--QNVR8I8sHE80Rc<RR#N#HRoM'Rj'0kFRMCk#8HRL0R#
RzRR4:RRRRHV58N8s8IH0=ERRR42oCCMsCN0
RRRRRRRRIDF_8sN8<sR=jR"jRj"&NRs8C_so25j;R
RRRRRRFRDIN_I8R8s<"=Rj"jjRI&RNs8_Cjo52R;
RCRRMo8RCsMCNR0Cz
4;RRRRzR.R:VRHR85N8HsI8R0E=2R.RMoCC0sNCR
RRRRRRFRDIN_s8R8s<"=RjRj"&NRs8C_soR548MFI0jFR2R;
RRRRRDRRFII_Ns88RR<=""jjRI&RNs8_C4o5RI8FMR0Fj
2;RRRRCRM8oCCMsCN0R;z.
RRRRRzdRH:RVNR58I8sHE80Rd=R2CRoMNCs0RC
RRRRRDRRFsI_Ns88RR<='Rj'&NRs8C_soR5.8MFI0jFR2R;
RRRRRDRRFII_Ns88RR<='Rj'&NRI8C_soR5.8MFI0jFR2R;
RCRRMo8RCsMCNR0Cz
d;RRRRzRcR:VRHR85N8HsI8R0E>2RdRMoCC0sNCR
RRRRRRFRDIN_s8R8s<s=RNs8_Cdo5RI8FMR0Fj
2;RRRRRRRRD_FII8N8s=R<R8IN_osC58dRF0IMF2Rj;R
RRMRC8CRoMNCs0zCRc
;
RRRR-Q-RV8R5HsM_CRo2sHCo#s0CRh7QRHk#MBoRpRi
RzRR6:RRRRHV5M8H_osC2CRoMNCs0RC
RRRRRbRRsCFO#5#RB,piRh7Q2CRLo
HMRRRRRRRRRRRRH5VRBRpi=4R''MRN8pRBiP'CC2M0RC0EMR
RRRRRRRRRRRRRRMRH_osCRR<=7;Qh
RRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMRFbsO#C#;R
RRMRC8CRoMNCs0zCR6R;
RzRRn:RRRRHV50MFRM8H_osC2CRoMNCs0RC
RRRRRRRRRHRRMC_so=R<Rh7Q;R
RRMRC8CRoMNCs0zCRn
;
RRRR-Q-RV8R5F_k0s2CoRosCHC#0smR7zkaR#oHMRpmBiR
RR(RzRRR:H5VR80Fk_osC2CRoMNCs0RC
RRRRRbRRsCFO#5#RmiBp,kRF0C_soL2RCMoH
RRRRRRRRRRRRRHV5pmBiRR='R4'NRM8miBp'CCPMR020MEC
RRRRRRRRRRRRRRRRz7ma=R<R0Fk_osC;R
RRRRRRRRRRMRC8VRH;R
RRRRRRMRC8sRbF#OC#R;
RCRRMo8RCsMCNR0Cz
(;RRRRzRUR:VRHRF5M0FR8ks0_CRo2oCCMsCN0
RRRRRRRRRRRRz7ma=R<R0Fk_osC;R
RRMRC8CRoMNCs0zCRU
;
RRRR-Q-RVsR5Ns88_osC2CRso0H#C)sRq)77RHk#MmoRB
piRRRRzRgR:VRHRN5s8_8ss2CoRMoCC0sNCR
RRRRRRsRbF#OC#mR5B,piR7)q7R)2LHCoMR
RRRRRRRRRRVRHRB5mp=iRR''4R8NMRpmBiP'CC2M0RC0EMR
RRRRRRRRRRRRRRNRs8C_so=R<R7)q7N)58I8sHE80-84RF0IMF2Rj;R
RRRRRRRRRRMRC8VRH;R
RRRRRRMRC8sRbF#OC#R;
RCRRMo8RCsMCNR0Cz
g;RRRRzR4j:VRHRF5M0NRs8_8ss2CoRMoCC0sNCR
RRRRRRRRRRNRs8C_so=R<R7)q7
);RRRRCRM8oCCMsCN0Rjz4;R
RRRRRRRR
R-RR-VRQRN5I8_8ss2CoRosCHC#0sqRW7R7)kM#HopRBiR
RR4Rz6:RRRRHV58IN8ss_CRo2oCCMsCN0
RRRRRRRRFbsO#C#Rp5BiW,Rq)772CRLo
HMRRRRRRRRRRRRH5VRBRpi=4R''MRN8pRBiP'CC2M0RC0EMR
RRRRRRRRRRRRRRNRI8C_so=R<R7Wq7N)58I8sHE80-84RF0IMF2Rj;R
RRRRRRRRRRMRC8VRH;R
RRRRRRMRC8sRbF#OC#R;
RCRRMo8RCsMCNR0Cz;46
RRRRnz4RH:RVMR5FI0RNs88_osC2CRoMNCs0RC
RRRRRRRRRIRRNs8_C<oR=qRW7;7)
RRRR8CMRMoCC0sNC4Rzn
;
RRRR-t-RCsMCNR0C0REC)RqvODCD#MRN8CR#D0CORoDFHRO
RzRR4:4RRsVFRHHRMkRMlC_ODRD#8MFI0jFRRMoCC0sNCR
RRRRRR-R-RRQV58N8s8IH0>ERRRc2M8CCRR0FONsC0ICRsCH0RNCMLRDCNRM8Fbk0kC0RMDNLCCR#D0CORoDFHRO
RRRRRzRR4:.RRRHV58N8s8IH0>ERRRc2oCCMsCN0
RRRRRRRRRRRRRRRR0Fk_5CMH<2R=4R''ERIC5MRs_N8s5CoNs88I0H8ER-48MFI0cFR2RR=HC2RDR#C';j'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RWRCIEMIR5Ns8_CNo58I8sHE80-84RF0IMF2RcRH=R2DRC#'CRj
';RRRRRRRRCRM8oCCMsCN0R.z4;R
RRRRRR-R-RRQV58N8s8IH0<ER=2RcRRMFI0sHCMRCNCLDRRFsFbk0kC0RMDNLCCR#D0CORoDFHMORCCC88R
RRRRRR4RzdRR:H5VRNs88I0H8E=R<RRc2oCCMsCN0
RRRRRRRRRRRRRRRR0Fk_5CMH<2R=4R''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=W
 ;RRRRRRRRRRRRCRM8oCCMsCN0Rdz4;R
RR-R-RCtMsCN0RC0ERv)qRDOCDN#RM08Rs#H-0CN0#R
RRRRRR4RzcRR:VRFs[MRHRH5I8R0E-2R4RI8FMR0FjCRoMNCs0RC
RRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)Rzq:vRRLDNCHDR#1R"7Ra"&MRH0CCosl'HN5oCI0H8E&2RR""7RH&RMo0CCHs'lCNo54H*n&2RR""WRH&RMo0CCHs'lCNo5R[2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50E54H+2n*4,CR8b20E2RR&"RX"&MRH0CCosl'HN5oC[2+4;R
RRRRRRRRRRCRLo
HMRRRRRRRRRRRRzv)q:qR)vX4n4
7RRRRRRRRRRRRRRRRRb0FsRblNRR57=H>RMC_so25[,jRqRR=>D_FII8N8s25j,4RqRR=>D_FII8N8s254,.RqRR=>D_FII8N8s25.,R
RRRRRRRRRRRRRRRRRRRRRRRRRq=dR>FRDIN_I858sdR2,7qu)j>R=RIDF_8sN8js527,Ru4)qRR=>D_FIs8N8s254,RR
RRRRRRRRRRRRRRRRRRRRRRRRR)7uq=.R>FRDIN_s858s.R2,7qu)d>R=RIDF_8sN8ds52W,R >R=R0Is_5CMHR2,
RRRRRRRRRRRRRRRRRRRRRRRRWRRBRpi=B>RpRi,7Rum=F>RkL0_kH#5,2[2;R
RRRRRRRRRRkRF0C_so25[RR<=F_k0L5k#H2,[RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRMRC8CRoMNCs0zCR4
c;RRRRRRRRCRM8oCCMsCN0R4z4;R
RRRRRRRRRRRRRRRRRRRRRRRRRR
RRCRM8NEsOHO0C0CksRD#CC_O0s;Nl
