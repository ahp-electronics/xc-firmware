--
@ER--RbBF$osHE50RO42RgRgg1b$MDHHO0R$,Q3MO
R--RDqDRosHER0#sCC#s8PC3-
-
R--fN]C8:CsR#//$DMbH0OH$N/lb0DN.Uj4J4.b/blNb#Cs/DOb8H/DLC/oMN_D0O0HC8/N8E3P8Ry4f-
-
-
-
R--oCCMsCN0RFbsbNNo0OCRC3DDRDONONkD0RC#OsNsHRC#LCN#8MRFRMoC/FbsbMRHb#k0

--DsHLNRs$HCCC;#
kCCRHC#C30D8_FOoH_n44cD3NDC;
M00H$bRo_NDCV#RHRo
SCsMCH5OR
#SSHRxC:MRH0CCos=R:RS4
2S;
b0FsRS5
SMoCFRk0:kRF00R#8F_Do;HO
bSSsFFbk:0RR0FkR8#0_oDFH
O;SFSOk:0RR0FkR8#0_oDFHPO_CFO0sH5#x4C-RI8FMR0Fj
2;SCSoMRHM:MRHR8#0_oDFHPO_CFO0sH5#x4C-RI8FMR0Fj
2;SsSbFMbHRH:RM0R#8F_Do_HOP0COF#s5H-xC4FR8IFM0R;j2
OSSH:MRRRHM#_08DHFoO
2;CRM8oDb_C;NV
s
NO0EHCkO0sLCRFCFDNFMRVbRo_NDCV#RHR#
SHNoMDoR0:0R#8F_Do_HOP0COF#s5H-xC4FR8IFM0R;j2
HS#oDMNR:0bR8#0_oDFHPO_CFO0sH5#x4C-RI8FMR0Fj
2;LHCoM0
Sb25jRR<=bbsFHjM52S;
0jo52=R<RMoCHjM52S;
O0Fk5Rj2<0=Ro25jRRFs550bjN2RMO8RH;M2Sb
SsCFO#5#RO,HMRFbsb,HMRMoCHRM,0Ro,0Rb2
PSSNNsHLRDCHRR:HCM0o;Cs
CSLo
HMSFSVsRRHH4MRRR0F#CHx-D4RF
FbS0SSb25HRR<=bbsFHHM52MRN8bR054H-2S;
SoS05RH2<o=RCMMH5RH2F5sRbbsFHHM52MRN8oR054H-2
2;SOSSF5k0H<2R=oR05RH2F5sR0Hb52MRN8HROM
2;SMSC8FRDF
b;S8CMRFbsO#C#;o
SCkMF0=R<R50o#CHx-;42
sSbFkbF0=R<R50b#CHx-;42
M
C8FRLFNDCM
;
---
-NROsRs$D	FFNNEC88RN8RCsIEH0RF0IRPDCCRD#FDVRFRF	NNEC8-
-R0HMCCsl80HNC8RN8#CsRCNsRbsHbRDCNC88s-#
-H
DLssN$CRHC
C;kR#CHCCC38#0_oDFH4O_43ncN;DD
0CMHR0$Ns88oHbR#o
SCsMCH5OR
#SSHRxC:MRH0CCos=R:R;.g
DSSC#NVHRxC:MRH0CCos=R:RSn
2S;
b0FsRS5
SkOF0RR:FRk0#_08DHFoOS;
S:8RR0FkR8#0_oDFHPO_CFO0sH5#x4C-RI8FMR0Fj
2;SRSN:MRHR8#0_oDFHPO_CFO0sH5#x4C-RI8FMR0Fj
2;SRSL:MRHR8#0_oDFHPO_CFO0sH5#x4C-RI8FMR0Fj
2;SHSOMRR:H#MR0D8_FOoH2C;
MN8R8o8sb
;
NEsOHO0C0CksRFLFDMCNRRFVNs88oHbR#S

VOkM0MHFRDONO0OMRF5OMN#0M#0RxD,RC#NVxRR:HCM0o2CsR0sCkRsMHCM0oRCsHS#
PHNsNCLDRNDCVb0l,MsO0RR:HCM0o;Cs
CSLo
HMSCSDNlV0b=R:RR#x/CRDNxV#;S
SH5VR5R#xlRF8DVCN#Rx2=2RjRC0EMS
SSMsO0=R:RNDCVb0lRS;
S#CDCSR
SOSsM:0R=DR5C0NVl+bRR;42
CSSMH8RVS;
S0sCkRsMs0OM;C
SMO8RNODOM
0;
FSOMN#0MD0RCONVM:0RR0HMCsoCRR:=OONDO5M0#CHx,CRDNHV#x;C2
V
Sk0MOHRFM0#EHDVCN#CHxRF5OMN#0MM0RRH:RMo0CCRs2skC0sHMRMo0CCHsR#P
SNNsHLRDC#:xRR0HMCsoC;L
SCMoH
HSSVMR5R5=RDVCNO-M04R220MECRS
SSR#x:#=RHRxClRF8DVCN#CHx;S
SSRHV5R#x=2RjRC0EMSR
S#SSx=R:RNDCVx#HC
;RSCSSMH8RVS;
S#CDCS
SSR#x:D=RC#NVH;xC
CSSMH8RVS;
S0sCkRsM#
x;S8CMRH0E#NDCVx#HC
;
SMVkOF0HMNRlG0LHRF5OMN#0MM0RRH:RMo0CCRs2skC0sHMRMo0CCHsR#P
SNNsHLRDClRNG:MRH0CCosS;
LHCoMS
SlRNG:5=RM2+4*NDCVx#HCRR-4S;
SRHV5GlNRR>=#CHx2ER0CSM
SNSlG=R:Rx#HC;-4
CSSMH8RVS;
S0sCkRsMl;NG
MSC8NRlG0LH;S

#MHoNoDRCLMN:0R#8F_Do_HOP0COF#s5H-xC4FR8IFM0R;j2
HS#oDMNRFbsb:NLR8#0_oDFHPO_CFO0sH5#x4C-RI8FMR0Fj
2;So#HMRNDO0HM:0R#8F_Do_HOP0COFDs5CONVM80RF0IMF2Rj;#
SHNoMDHROM:0LR8#0_oDFHPO_CFO0sC5DNMVO0FR8IFM0R;j2
HS#oDMNRHOsMR0:#_08DHFoOC_POs0F5x#HCFR8IFM0R;j2
HS#oDMNRMoCFRk0:0R#8F_Do;HO
HS#oDMNRFbsb0FkR#:R0D8_FOoH;S

ObFlFMMC0bRo_NDCV#RHRS
SoCCMsRHO5S
SSx#HCRR:HCM0o
CsS;S2
bSSFRs05S
SSMoCFRk0:kRF00R#8F_Do;HO
SSSbbsFFRk0:kRF00R#8F_Do;HO
SSSO0FkRF:Rk#0R0D8_FOoH_OPC05Fs#CHx-84RF0IMF2Rj;S
SSMoCH:MRRRHM#_08DHFoOC_POs0F5x#HCR-48MFI0jFR2S;
SsSbFMbHRH:RM0R#8F_Do_HOP0COF#s5H-xC4FR8IFM0R;j2
SSSORHM:MRHR8#0_oDFH;O2
MSC8FROlMbFC;M0
O
SFFlbM0CMR8N8sbHbDHCR#S
SoCCMsRHO5S
SSx#HCRR:HCM0o
CsS;S2
bSSFRs05S
SSkOF0RR:FRk0#_08DHFoOS;
SRS8:kRF00R#8F_Do_HOP0COF#s5H-xC4FR8IFM0R;j2
SSSNRR:H#MR0D8_FOoH_OPC05Fs#CHx-84RF0IMF2Rj;S
SS:LRRRHM#_08DHFoOC_POs0F5x#HCR-48MFI0jFR2S;
SHSOMRR:H#MR0D8_FOoH
2SS;C
SMO8RFFlbM0CM;S

ObFlFMMC0YRBuwAzRRH#
bSSFRs05S
SNRR:H#MR0D8_FOoH;S
SLRR:FRk0#_08DHFoOS
S2S;
CRM8ObFlFMMC0
;
So#HMRNDLLo,bRR:#_08DHFoOC_POs0F5x#HCR-48MFI0jFR2S;
#MHoNLDRoL0,b:0RR8#0_oDFHPO_CFO0sH5#x4C-RI8FMR0Fj
2;So#HMRNDoR,b:0R#8F_Do_HOP0COFDs5CONVM40-RI8FMR0Fj
2;So#HMRNDobL,LRR:#_08DHFoOC_POs0F5NDCV0OM-84RF0IMF2Rj;#
SHNoMDFRVFRR:#_08DHFoOL;
CMoH
o
SCLMNRR<=NMRN8;RL
sSbFLbNRR<=NsRFR
L;SMOH025jRR<=O;HM
HSOM50Lj<2R=HROM
;
SR--	bCCRC0ERLDNCRD##sEF0sRFRC0ERlMNCo#RC00RFDFRF
MoSRq:VRFsMMRHR0jRFCRDNMVO0R-4oCCMsCN0
OSSF0M#NRM0l0GLRH:RMo0CC:sR=NRlG0LH5;M2
OSSF0M#NRM0DxV#RH:RMo0CC:sR=ER0HC#DNHV#xMC52S;
SMOF#M0N0MRlL:0RR0HMCsoCRR:=DVCN#CHx*
M;SFSOMN#0MN0RDMDFC:#RR8#0_oDFHPO_CFO0sG5lL80RF0IMFMRlLR02:5=RFC0Es>#=R''42S;
LHCoMSR
S5Lol0ML2=R<RMoCNlL5M2L0;S
SLlb5M2L0RR<=bbsFNlL5M2L0;S
SL5o0l0ML2=R<R5Lol0ML2S;
S0Lb5LlM0<2R=bRL5LlM0
2;
-SS-NRODDOkNR0C0RECL-H0ICH#R#o'R8NMR#b'R8NMRVLkVRCs0lEC
ASS:FRVsRRlHlMRM+L04FR0RLlG0CRoMNCs0
CRSLSSol052=R<RMoCNlL52sRFRs5bFLbN5Rl2NRM8L5o0l2-42S;
StSAXB:RYzuAwFRbsl0RN5bRL5o0lR2,Llo52
2;SLSSbl052=R<RFbsb5NLlN2RML8Rbl05-;42
SSSA:uXRuBYARzwb0FsRblNRb5L025l,bRL52l2;S
SCRM8oCCMsCN0;S

SR--O$FbRC0ERNDCVR'#oMRN8RRbVlsFRC0ERRLoNRM8LSb
S5oLM<2R=oRL5LlG0
2;SLSb5RM2<L=RbG5lL;02
S
S-L-RkCVVsER0CNROsRs$H5MRVlsFRC0ERsONso$RCsMCNs0F2SR
SRB:H5VRM=R/RRj2oCCMsCN0RS
SSXBA:YRBuwAzRsbF0NRlbH5OMM052O,RHLM052M2;S
SCRM8oCCMsCN0;S

SR--OONDk0DNCER0CHRL0H-I#OCRNHssCV#RsRFl0RECL-H0ICH#R'ob#MRN8HROMS
S8H:RVlR5GRL0>MRlLR02oCCMsCN0RS
SSRC:VRFslMRHRLlG0FR8IFM0RLlM0R+4oCCMsCN0
SSSSHOsMl052=R<R5Lol2-4RRFs5MOH0ML52MRN8bRL54l-2
2;SCSSMo8RCsMCN;0C
CSSMo8RCsMCN;0C
OSSs0HM5LlM0<2R=HROM50LM
2;
-SS-NRODDOkNR0C0REC#
klS5S8l0GLRI8FMR0Fl0ML2=R<RlN5GRL08MFI0lFRM2L0
SSSGRFsLG5lL80RF0IMFMRlLR02GRFsOMsH0G5lL80RF0IMFMRlL;02
MSC8CRoMNCs0
C;
-S-RMoCC0sNCER0CNROsCsH#O
Soo:RbC_DNSV
SMoCCOsHRblNRS5
SHS#x=CR>CRDNMVO0S
S2S
Sb0FsRblNRS5
SCSoM0FkRR=>oFCMk
0,SbSSsFFbk=0R>sRbFkbF0S,
SFSOk=0R>HROMD05CONVM80RF0IMF2R4,S
SSMoCH=MR>LRo5NDCV0OM-84RF0IMF2Rj,S
SSFbsbRHM=b>RLC5DNMVO0R-48MFI0jFR2S,
SHSOM>R=RMOH
2SS;S

O0FkRR<=O0HM5NDCV0OM2
;
CRM8LDFFC;NM
-
-
R--VDkDRbsHbRDCNC88s-
-
LDHs$NsRCHCCk;
#HCRC3CC#_08DHFoO4_4nNc3D
D;CHM00N$R8H8sbCbDR
H#SMoCCOsHRS5
Sx#HCRR:HCM0oRCs:g=R
;S2
FSbs50R
OSSFRk0:kRF00R#8F_Do;HO
8SSRF:Rk#0R0D8_FOoH_OPC05Fs#CHx-84RF0IMF2Rj;S
SNRR:H#MR0D8_FOoH_OPC05Fs#CHx-84RF0IMF2Rj;S
SLRR:H#MR0D8_FOoH_OPC05Fs#CHx-84RF0IMF2Rj;S
SORHM:MRHR8#0_oDFH;O2
8CMR8N8sbHbD
C;
ONsECH0Os0kCFRLFNDCMVRFR8N8sbHbDHCR##
SHNoMDCRoM0FkR#:R0D8_FOoH;#
SHNoMDsRbFkbF0RR:#_08DHFoOS;
#MHoNODRH:M0R8#0_oDFHPO_CFO0sH5#x8CRF0IMF2Rj;#
SHNoMDCRoM:NLR8#0_oDFHPO_CFO0sH5#x4C-RI8FMR0Fj
2;So#HMRNDbbsFNRL:#_08DHFoOC_POs0F5x#HCR-48MFI0jFR2L;
CMoH
CSoMRNL<N=RR8NMR
L;SFbsbRNL<N=RRRFsLS;
O0HM5x#HCFR8IFM0RR42<5=RbbsFNNLRMO8RH5M0#CHx-84RF0IMF2Rj2sRFRMoCN
L;SMOH025jRR<=O;HM
RS8<N=RRsGFRGLRFOsRH5M0#CHx-84RF0IMF2Rj;O
SFRk0<O=RH5M0#CHx2C;
ML8RFCFDN
M;

---0-RFDbRCDPCR0CMHR0$VRFsNC88sCRoMNCs0
Fs-k-R#RC#sbHbDHCRVCRD#0#RERNMv)qXQpuu C,RDR#Ck##CRsONsD$RFNF	E8CN

--DsHLNRs$HCCC;kR
#HCRC3CC#_08DHFoO4_4nNc3D
D;CHM00q$R7H7R#R
RRCRoMHCsOH5I8R0E:MRH0CCos=R:R24n;-R-Ro[N
RRRRsbF0:5qRRHM#_08DHFoOC_POs0F58IH0-ER4FR8IFM0R;j2
RRRRRRRR:RARRHM#_08DHFoOC_POs0F58IH0-ER4FR8IFM0R;j2
RRRRRRRRQRBhRR:H#MR0D8_FOoH;R
RRRRRRmRRRF:Rk#0R0D8_FOoH_OPC05FsI0H8E4R-RI8FMR0Fj
2;RRRRRRRRRzBmaF:Rk#0R0D8_FOoH2C;
Mq8R7
7;
ONsECH0Os0kCCRODDD_CDPCRRFVqR77HS#
O#FM00NMRXvq)uQup: RR0HMCsoCRR:=U
;
SMVkOF0HMNRODCODNHV#x5CRO#FM00NMRRI:HCM0o2CsR0sCkRsMHCM0oRCsHS#
SsPNHDNLCPRsNHD:Mo0CC:sR=;R4
CSLo
HMSESIHRDC5NsPDRR*sDPNRI<R2FRDFSb
SPSsN:DR=PRsN+DRR
4;SMSC8FRDF
b;SVSHRP5sN<DRRRc20MECRS
SSNsPD=R:RRc;
CSSMH8RVS;
S0sCkRsMsDPN;C
SMO8RNDDOC#NVH;xC
O
SFFlbM0CMR8N8sRobHS#
SMoCCOsHRS5
SHS#x:CRR0HMCsoC;S
SSNDCVx#HCRR:HCM0oRCs
2SS;S
Sb0FsRS5
SFSOk:0RR0FkR8#0_oDFH
O;S8SSRF:Rk#0R0D8_FOoH_OPC05Fs#CHx-84RF0IMF2Rj;S
SS:NRRRHM#_08DHFoOC_POs0F5x#HCR-48MFI0jFR2S;
SRSL:MRHR8#0_oDFHPO_CFO0sH5#x4C-RI8FMR0Fj
2;SOSSH:MRRRHM#_08DHFoOS
S2S;
CRM8ObFlFMMC0
;
SlOFbCFMMN0R8H8sbCbDR
H#SCSoMHCsO
R5S#SSHRxC:MRH0CCosS
S2S;
SsbF0
R5SOSSFRk0:kRF00R#8F_Do;HO
SSS8RR:FRk0#_08DHFoOC_POs0F5x#HCR-48MFI0jFR2S;
SRSN:MRHR8#0_oDFHPO_CFO0sH5#x4C-RI8FMR0Fj
2;SLSSRH:RM0R#8F_Do_HOP0COF#s5H-xC4FR8IFM0R;j2
SSSORHM:MRHR8#0_oDFHSO
S
2;S8CMRlOFbCFMM
0;
oLCHSM
LRN:H5VRI0H8ERR>v)qXQpuu o2RCsMCN
0CS4SN:8RN8bsoRS
SSMoCCOsHRblNRS5
S#SSHRxC=I>RHE80,S
SS-S-RNDCVx#HC>R=RDONONDCVx#HCH5I820E
SSSSNDCVx#HC>R=RSc
S
S2SbSSFRs0lRNb5S
SSFSOk=0R>FROk
0,SSSS8>R=R
F,SSSSN>R=R
N,SSSSL>R=R
L,SSSSORHM=O>RHSM
S;S2
MSC8CRoMNCs0
C;
NS#:VRHRH5I8R0E<v=RqQX)u up2CRoMNCs0SC
S:N4R8N8sbHbD
CRSoSSCsMCHlORN5bR
SSSSx#HC>R=R8IH0SE
S
S2SbSSFRs0lRNb5S
SSFSOk=0R>FROk
0,SSSS8>R=R
F,SSSSN>R=R
N,SSSSL>R=R
L,SSSSORHM=O>RHSM
S;S2
MSC8CRoMNCs0
C;
8CMRDOCDC_DP;CD




