--
@ER--B$FbsEHo0OR52gR4g-cRRj.jd$R1MHbDO$H0ROQM
R--fN]C8:CsR#//$DMbH0OH$N/lb0DN.Uj4J4.b/blNb#Cs/0N0/LDH/MoC_OFsN/cCs_Nls3_IPyE84
Rf-
-


-----
-kR7NbD-FRs0)RqvIEH0Rb#CC0sNC7Rq71) 1FRVsCRsNN8RMI8RsCH0
R--aoNsC:0RROpkCRM0-)RmBdqRB-
-
LDHs$NsRCHCCk;
#HCRC3CC#_08DHFoO4_4nNc3D
D;kR#CHCCC38#0_oDFH#O_HCoM8D3NDk;
#HCRC3CC#_08DHFoOs_NH30EN;DD
LDHs$NsROFsN
d;kR#CFNsOds3FOFNOlNb3D
D;CHM00)$Rq)v__HWR#R
RRCRoMHCsO
R5RRRRRRRRVHNlDR$:#H0sM:oR=MR"F"MC;R
RRRRRRHRI8R0E:MRH0CCos=R:RR(;
RRRRRRRR8N8s8IH0:ERR0HMCsoCRR:=(R;RRRRRR-R-RoLHRFCMkRoEVRFs80CbER
RRRRRRCR8bR0E:MRH0CCos=R:R.R4UR;
RRRRR8RRF_k0sRCo:FRLFNDCM=R:RDVN#RC;RRRR-E-RNF#Rkk0b0CRsoR
RRRRRRHR8MC_soRR:LDFFCRNM:V=RNCD#;RRRR-RR-NRE#NR80HNRM0bkRosC
RRRRRRRR8sN8ss_C:oRRFLFDMCNRR:=V#NDCR;RR-R-R8ENRNsC88RN8#sC#CRsoR
RRRRRRNRI8_8ssRCo:FRLFNDCM=R:RDVN#RCRR-RR-NRE8sRIHR0CNs88CR##s
CoRRRRRRRR2R;
RbRRFRs05R
RRRRRRmR7zRaR:kRF00R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj;R
RRRRRRqR)7R7):MRHR0R#8F_Do_HOP0COFNs58I8sHE80-84RF0IMF2Rj;R
RRRRRRQR7hRRR:MRHR0R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj;R
RRRRRRqRW7R7):MRHR0R#8F_Do_HOP0COFNs58I8sHE80-84RF0IMF2Rj;R
RRRRRR RWRRRR:MRHR0R#8F_Do;HORRRRR-RR-sRIHR0CCLMNDVCRFssRNRl
RRRRRBRRpRiRRH:RM#RR0D8_FOoH;RRRRRRR-O-RD	FORsVFRlsN,8RN8Rs,8
HMRRRRRRRRmiBpRRR:HRMR#_08DHFoORRRRRRRRR--FRb0OODF	FRVsFR8kR0
RRRRR2RR;M
C8MRC0$H0Rv)q_W)_;-

--
-RswH#H0RlCbDl0CMNF0HMkRl#L0RCNROD8DCRONsE-j
-s
NO0EHCkO0sNCRsjOERRFV)_qv)R_WHO#
F0M#NRM0M_klODCD#C_8C:bRR0HMCsoCRR:=5C58bR0E-2R4/2d.;RRRRRRRR-R-RFyRVFRsIF#RVBR7 Xd.cCRODRD#M8CCCO8
F0M#NRM0M_klODCD#H_I8:CRR0HMCsoCRR:=5H5I8R0E-2R4/;c2RRRRRRRRR-R-RFyRVFRODMkl#VRFR 7Bdc.XRDOCDM#RCCC88$
0bFCRkL0_k0#_$RbCHN#Rs$sNRk5MlC_OD_D#8bCCRI8FMR0Fj5,RM_klODCD#H_I8cC*2R+d8MFI0jFR2VRFR8#0_oDFH
O;#MHoNFDRkL0_k:#RR0Fk_#Lk_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RVFR8k50RHkMb0FR0RH0s-N#002C#
o#HMRNDF_k0CRMRRRR:#_08DHFoOC_POs0F5lMk_DOCD8#_CRCb8MFI0jFR2R;R-C-RMDNLCV#RF0sRs#H-0CN0#H
#oDMNRCIbjM_CR:RRR8#0_oDFHPO_CFO0sk5MlC_OD_D#8bCCRI8FMR0FjR2;RR--I0sHCMRCNCLD#FRVsNRCOsERFFIRVqR)vCROD
D##MHoNIDRb_C4CRMRR#:R0D8_FOoH_OPC05FsM_klODCD#C_8C8bRF0IMF2Rj;-RR-sRIHR0CCLMNDRC#VRFsCENORIsFRRFV)RqvODCD#H
#oDMNR_HMsRCoR:RRR8#0_oDFHPO_CFO0sH5I8+0EdFR8IFM0R;j2RRRRRRRRRR--k8#CRR0FsHCo#s0CRh7QRH
#oDMNR_W )4 tR:RRR8#0_oDFH
O;#MHoNHDRMC_soR4RR#:R0D8_FOoH_OPC05FsI0H8ER+d8MFI0jFR2R;RR#R
HNoMDkRF0C_soRRR:0R#8F_Do_HOP0COFIs5HE80+8dRF0IMF2Rj;RRRRRRRR-R-RCk#8FR0RosCHC#0smR7z#a
HNoMDNRs8C_soRRR:0R#8F_Do_HOP0COFNs58I8sHE80-84RF0IMF2Rj;RRRR-R-RCk#8FR0RosCHC#0sqR)7
7)#MHoNIDRNs8_CRoRR#:R0D8_FOoH_OPC05FsNs88I0H8ER-48MFI0jFR2R;RR-RR-#RkC08RFCRso0H#CWsRq)77
o#HMRNDD_FIs8N8sRR:#_08DHFoOC_POs0F58cRF0IMF2Rj;RRRRRRRRRRRRRRR-s-RNs88R0LH#MRHbRk00)FRqOvRC#DDRR56L#H0RJsCkCHs8#2
HNoMDFRDIN_I8R8s:0R#8F_Do_HOP0COFcs5RI8FMR0FjR2;RRRRRRRRRRRRR-R-R8IN8LsRHR0#HkMb0FR0Rv)qRDOCD5#R6HRL0s#RCHJks2C8
b0$ClR0b8_N80s_$RbCHN#Rs$sNRk5MlC_OD_D#8bCCRI8FMR0FjF2RV0R#8F_Do_HOP0COF5sRgFR8IFM0R;j2
o#HMRND0_lbNs88RRR:0_lbNs88_b0$C
;
LHCoMR

R-RR-VRQR8N8s8IH0<ERRN6R#o#HMjR''FR0RkkM#RC8L#H0
RRRRRz4RH:RVNR58I8sHE80R4=R2CRoMNCs0RC
RRRRRDRRFsI_Ns88RR<="jjjj&"RR8sN_osC5;j2
RRRRRRRRIDF_8IN8<sR=jR"j"jjRI&RNs8_Cjo52R;
RCRRMo8RCsMCNR0Cz
4;RRRRzR.R:VRHR85N8HsI8R0E=2R.RMoCC0sNCR
RRRRRRFRDIN_s8R8s<"=Rj"jjRs&RNs8_C4o5RI8FMR0Fj
2;RRRRRRRRD_FII8N8s=R<Rj"jj&"RR8IN_osC584RF0IMF2Rj;R
RRMRC8CRoMNCs0zCR.R;
RzRRd:RRRRHV58N8s8IH0=ERRRd2oCCMsCN0
RRRRRRRRIDF_8sN8<sR=jR"j&"RR8sN_osC58.RF0IMF2Rj;R
RRRRRRFRDIN_I8R8s<"=RjRj"&NRI8C_soR5.8MFI0jFR2R;
RCRRMo8RCsMCNR0Cz
d;RRRRzRcR:VRHR85N8HsI8R0E=2RcRMoCC0sNCR
RRRRRRFRDIN_s8R8s<'=Rj&'RR8sN_osC58dRF0IMF2Rj;R
RRRRRRFRDIN_I8R8s<'=Rj&'RR8IN_osC58dRF0IMF2Rj;R
RRMRC8CRoMNCs0zCRcR;
RzRR6:RRRRHV58N8s8IH0>ERRRc2oCCMsCN0
RRRRRRRRIDF_8sN8<sR=NRs8C_soR5c8MFI0jFR2R;
RRRRRDRRFII_Ns88RR<=I_N8s5CocFR8IFM0R;j2
RRRR8CMRMoCC0sNC6Rz;R

R-RR-VRQRH58MC_sos2RC#oH0RCs7RQhkM#HopRBiR
RRnRzRRR:H5VR8_HMs2CoRMoCC0sNCR
RRRRRRsRbF#OC#BR5pRi,72QhRoLCHRM
RRRRRRRRRHRRVBR5p=iRR''4R8NMRiBp'CCPMR020MEC
RRRRRRRRRRRRRRRR_HMsRCo<5=R"jjjj&"RRh7Q2R;
RRRRRRRRRCRRMH8RVR;
RRRRRCRRMb8RsCFO#
#;RRRRCRM8oCCMsCN0R;zn
RRRRRz(RH:RVMR5F80RHsM_CRo2oCCMsCN0
RRRRRRRRRRRR_HMsRCo<5=R"jjjj&"RRh7Q2R;
RCRRMo8RCsMCNR0Cz
(;
RRRRR--Q5VRs8N8sC_sos2RC#oH0RCs)7q7)#RkHRMoB
piRRRRzR4jRH:RVsR5Ns88_osC2CRoMNCs0RC
RRRRRbRRsCFO#5#RmiBp,qR)727)RoLCHRM
RRRRRRRRRHRRVmR5BRpi=4R''MRN8BRmpCi'P0CM2ER0CRM
RRRRRRRRRRRRRsRRNs8_C<oR=qR)757)Ns88I0H8ER-48MFI0jFR2R;
RRRRRRRRRCRRMH8RVR;
RRRRRCRRMb8RsCFO#
#;RRRRCRM8oCCMsCN0Rjz4;R
RR4Rz4RR:H5VRMRF0s8N8sC_soo2RCsMCN
0CRRRRRRRRRRRRs_N8sRCo<)=Rq)7758N8s8IH04E-RI8FMR0Fj
2;RRRRCRM8oCCMsCN0R4z4;R
RRRRRRRR
R-RR-VRQRN5I8_8ss2CoRosCHC#0sqRW7R7)kM#HopRBiR
RR4Rz.:RRRRHV58IN8ss_CRo2oCCMsCN0
RRRRRRRRFbsO#C#Rp5BiW,Rq)772CRLo
HMRRRRRRRRRRRRH5VRBRpi=4R''MRN8pRBiP'CC2M0RC0EMR
RRRRRRRRRRRRRRNRI8C_so=R<R7Wq7N)58I8sHE80-84RF0IMF2Rj;R
RRRRRRRRRRMRC8VRH;R
RRRRRRMRC8sRbF#OC#R;
RCRRMo8RCsMCNR0Cz;4.
RRRRdz4RH:RVMR5FI0RNs88_osC2CRoMNCs0RC
RRRRRRRRRIRRNs8_C<oR=qRW7;7)
RRRR8CMRMoCC0sNC4Rzd
;
RRRR-t-RCsMCNR0C0REC)RqvODCD#MRN8CR#D0CORoDFHRO
RzRR4:cRRsVFRHHRMkRMlC_OD_D#8bCCRI8FMR0FjCRoMNCs0RC
R-RR-kRAHRD8Fbk0kC0RMDNLCCR#D0CORoDFHRO
RRRRR-RR-VRQR85N8HsI8R0E>6R42NROMR'0kR#CNpR1QOBRC
DDRRRRRRRRmn 4RH:RVNR58I8sHE80R4>R6o2RCsMCN
0CRRRRRRRRRRRRRRRRF_k0CHM52=R<R''4RCIEMsR5Ns8_CNo58I8sHE80-84RF0IMF2R6RH=R2DRC#'CRj
';RRRRRRRRCRM8oCCMsCN0R4m nR;
RRRRR-RR-VRQR85N8HsI8R0E>2R6R7qhR85N8HsI8R0E<4=R6k2R#NNRRQ1pBCRODRD
RRRRRmRR R46:VRHR85N8HsI8R0E=6R42CRoMNCs0RC
RRRRRRRRRRRRR0RRlNb_858sHg25RI8FMR0Fj<2R=mRhaF5OM#P_0D8_FOoH_OPC05FsH4,RjR22XRm)s_N8s5CoNs88I0H8ER-48MFI06FR2R;
RRRRRRRRRRRRR1RRq_h74:6RRh1q7R4jb0FsRblNRR5q=0>RlNb_858sHj252A,RRR=>0_lbNs8855H24R2,B>R=Rb0l_8N8s25H5,.2R=7R>lR0b8_N8Hs5225d,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR= R>lR0b8_N8Hs5225c,RRw=0>RlNb_858sH6252t,RRR=>0_lbNs8855H2nR2,]>R=Rb0l_8N8s25H5,(2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR=QR>lR0b8_N8Hs5225U,RRK=0>RlNb_858sHg252Z,RRR=>F_k0CHM52
2;RRRRRRRRCRM8oCCMsCN0R4m 6R;
RRRRRmRR R4c:VRHR85N8HsI8R0E=cR42CRoMNCs0RC
RRRRRRRRRRRRR0RRlNb_858sHU25RI8FMR0Fj<2R=mRhaF5OM#P_0D8_FOoH_OPC05FsHg,R2X2Rms)RNs8_CNo58I8sHE80-84RF0IMF2R6;R
RRRRRRRRRRRRRRqR1h47_cRR:17qh4bjRFRs0lRNb5=qR>lR0b8_N8Hs5225j,RRA=0>RlNb_858sH4252B,RRR=>0_lbNs8855H2.R2,7>R=Rb0l_8N8s25H5,d2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR >R=Rb0l_8N8s25H5,c2R=wR>lR0b8_N8Hs52256,RRt=0>RlNb_858sHn252],RRR=>0_lbNs8855H2(R2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRQ>R=Rb0l_8N8s25H5,U2R=KR>4R''Z,RRR=>F_k0CHM52
2;RRRRRRRRCRM8oCCMsCN0R4m cR;
RRRRRmRR R4d:VRHR85N8HsI8R0E=dR42CRoMNCs0RC
RRRRRRRRRRRRR0RRlNb_858sH(25RI8FMR0Fj<2R=mRhaF5OM#P_0D8_FOoH_OPC05FsHU,R2X2Rms)RNs8_CNo58I8sHE80-84RF0IMF2R6;R
RRRRRRRRRRRRRRqR1h47_dRR:17qhUbRRFRs0lRNb5=qR>lR0b8_N8Hs5225j,RRA=0>RlNb_858sH4252B,RRR=>0_lbNs8855H2.R2,7>R=Rb0l_8N8s25H5,d2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR >R=Rb0l_8N8s25H5,c2R=wR>lR0b8_N8Hs52256,RRt=0>RlNb_858sHn252],RRR=>0_lbNs8855H2(R2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRZ>R=R0Fk_5CMH;22
RRRRRRRR8CMRMoCC0sNC Rm4
d;RRRRRRRRm. 4RH:RVNR58I8sHE80R4=R.o2RCsMCN
0CRRRRRRRRRRRRRRRR0_lbNs8855H2nFR8IFM0RRj2<h=RmOa5F_MP#_08DHFoOC_POs0F5RH,(R22XRm)s_N8s5CoNs88I0H8ER-48MFI06FR2R;
RRRRRRRRRRRRR1RRq_h74:.RRh1q7RURb0FsRblNRR5q=0>RlNb_858sHj252A,RRR=>0_lbNs8855H24R2,B>R=Rb0l_8N8s25H5,.2R=7R>lR0b8_N8Hs5225d,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR= R>lR0b8_N8Hs5225c,RRw=0>RlNb_858sH6252t,RRR=>0_lbNs8855H2nR2,]>R=R''4,RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRZ=F>RkC0_M25H2R;
RRRRRCRRMo8RCsMCNR0Cm. 4;R
RRRRRR Rm4:4RRRHV58N8s8IH0=ERR244RMoCC0sNCR
RRRRRRRRRRRRRRlR0b8_N8Hs52R568MFI0jFR2=R<Rahm5MOFP0_#8F_Do_HOP0COFHs5,2Rn2mRX)NRs8C_so85N8HsI8-0E4FR8IFM0R;62
RRRRRRRRRRRRRRRRh1q74_4R1:Rqnh7RFRbsl0RN5bRq>R=Rb0l_8N8s25H5,j2R=AR>lR0b8_N8Hs52254,RRB=0>RlNb_858sH.2527,RRR=>0_lbNs8855H2d
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR RRRR=>0_lbNs8855H2cR2,w>R=Rb0l_8N8s25H5,62R=ZR>kRF0M_C52H2;R
RRRRRRMRC8CRoMNCs0mCR ;44
RRRRRRRR4m jRR:H5VRNs88I0H8ERR=4Rj2oCCMsCN0
RRRRRRRRRRRRRRRRb0l_8N8s25H58cRF0IMF2RjRR<=h5maOPFM_8#0_oDFHPO_CFO0s,5HR262R)XmR8sN_osC58N8s8IH04E-RI8FMR0F6
2;RRRRRRRRRRRRRRRR17qh_R4j:qR1hR7nRsbF0NRlbqR5RR=>0_lbNs8855H2jR2,A>R=Rb0l_8N8s25H5,42R=BR>lR0b8_N8Hs5225.,RR7=0>RlNb_858sHd252R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR =0>RlNb_858sHc252w,RRR=>',4'R=ZR>kRF0M_C52H2;R
RRRRRRMRC8CRoMNCs0mCR ;4j
RRRRRRRRgm RRR:H5VRNs88I0H8ERR=go2RCsMCN
0CRRRRRRRRRRRRRRRR0_lbNs8855H2dFR8IFM0RRj2<h=RmOa5F_MP#_08DHFoOC_POs0F5RH,cR22XRm)s_N8s5CoNs88I0H8ER-48MFI06FR2R;
RRRRRRRRRRRRR1RRq_h7gRR:17qhcRRRb0FsRblNRR5q=0>RlNb_858sHj252A,RRR=>0_lbNs8855H24R2,B>R=Rb0l_8N8s25H5,.2R=7R>lR0b8_N8Hs5225d,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR=ZR>kRF0M_C52H2;R
RRRRRRMRC8CRoMNCs0mCR 
g;RRRRRRRRmR URH:RVNR58I8sHE80RU=R2CRoMNCs0RC
RRRRRRRRRRRRR0RRlNb_858sH.25RI8FMR0Fj<2R=mRhaF5OM#P_0D8_FOoH_OPC05FsHd,R2X2Rms)RNs8_CNo58I8sHE80-84RF0IMF2R6;R
RRRRRRRRRRRRRRqR1hU7_R1:Rqch7RbRRFRs0lRNb5=qR>lR0b8_N8Hs5225j,RRA=0>RlNb_858sH4252B,RRR=>0_lbNs8855H2.R2,7>R=R''4,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR=ZR>kRF0M_C52H2;R
RRRRRRMRC8CRoMNCs0mCR 
U;RRRRRRRRmR (RH:RVNR58I8sHE80R(=R2CRoMNCs0RC
RRRRRRRRRRRRR0RRlNb_858sH425RI8FMR0Fj<2R=mRhaF5OM#P_0D8_FOoH_OPC05FsH.,R2X2Rms)RNs8_CNo58I8sHE80-84RF0IMF2R6;R
RRRRRRRRRRRRRRqR1h(7_R1:Rq.h7RbRRFRs0lRNb5=qR>lR0b8_N8Hs5225j,RRA=0>RlNb_858sH4252Z,RRR=>F_k0CHM52
2;RRRRRRRRCRM8oCCMsCN0R(m ;R
RRRRRR Rmn:RRRRHV58N8s8IH0=ERRRn2oCCMsCN0
RRRRRRRRRRRRRRRR0Fk_5CMH<2R=4R''ERIC5MRs_N8s5Co6=2RRMOFP0_#8F_Do_HOP0COFHs5,542jR22CCD#R''j;R
RRRRRRMRC8CRoMNCs0mCR 
n;RRRR-Q-RVNR58I8sHE80RR<=6M2RFkRF00bkRNCMLRDC#CCDOD0RFOoHRCMC8
C8RRRRRRRRmR 6:VRHR85N8HsI8R0E<6=R2CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_M25HRR<=';4'
RRRRRRRR8CMRMoCC0sNC Rm6
;
RRRR-Q-RVNR58I8sHE80Rg>R2#RkCuRW 0jRFCR8OCF8R8N8s#C#R0LH#RRn0FEskRoEgMRN8uRW 04RFCR8OCF8R0LH#jR4RR+
RRRRRWRR R4j:VRHR85N8HsI8R0E>2RgRMoCC0sNCR
RRRRRRRRRRRRRRbRICCj_M25HRR<='R4'IMECRN5I8C_soR5U8MFI06FR2RR=OPFM_8#0_oDFHPO_CFO0s,5H.5j2dFR8IFM0R2j2R#CDCjR''R;
RRRRRRRRRRRRRIRRb_C4CHM52=R<R''4RCIEMIR5Ns8_CNo58I8sHE80-84RF0IMF2RgRO=RF_MP#_08DHFoOC_POs0F5.H,jN258I8sHE80-8nRF0IMF2Rc2DRC#'CRj
';RRRRRRRRRRRRCRM8oCCMsCN0R4W jR;
R-RR-VRQR85N8HsI8R0E=RRUFgsR2#RkCuRW 0jRFCR8OCF8R8N8s#C#R0LH#RRn0FEskRoEgR
RRRRRR RWg:RRRRHV585N8HsI8R0E=2RURRm)58N8s8IH0=ERR2g2RMoCC0sNCR
RRRRRRRRRRRRRRbRICCj_M25HRR<='R4'IMECRN5I8C_so85N8HsI8-0E4FR8IFM0RR62=2RHR#CDCjR''R;
RRRRRRRRRRRRRIRRb_C4CHM52=R<R''4;R
RRRRRRRRRRMRC8CRoMNCs0WCR 
g;RRRR-Q-RVNR58I8sHE80R(=R2#RkCuRW 0jRFCR8OCF8RC0EREn0R8N8s#C#R0LHRW&RuR 408FRC8OFCER0C0R(E8RN8#sC#HRL0R
RRRRRR RW(:RRRRHV58N8s8IH0=ERRR(2oCCMsCN0
RRRRRRRRRRRRRRRRCIbjM_C5RH2<'=R4I'RERCM58IN_osC5R62=FROM#P_0D8_FOoH_OPC05FsH2,.52j2R#CDCjR''R;
RRRRRRRRRRRRRIRRb_C4CHM52=R<R''4RCIEMIR5Ns8_Cno52RR=OPFM_8#0_oDFHPO_CFO0s,5H.4252C2RDR#C';j'
RRRRRRRR8CMRMoCC0sNC RW(R;
R-RR-VRQR85N8HsI8R0E=2RnRCk#R WujFR0RO8CFR8C0RECnR0ENs88CR##L
H0RRRRRRRRWR nRH:RVNR58I8sHE80Rn=R2CRoMNCs0RC
RRRRRRRRRRRRRIRRb_CjCHM52=R<R''4RCIEMIR5Ns8_C6o52RR=OPFM_8#0_oDFHPO_CFO0s,5H4j252C2RDR#C';j'
RRRRRRRRRRRRRRRRCIb4M_C5RH2<'=R4
';RRRRRRRRCRM8oCCMsCN0RnW ;R
RR-R-RRQV58N8s8IH0<ER=2R6RRMFI0sHCMRCNCLDRD#CCRO0DHFoOCRMC88C
RRRRRRRR6W RRR:H5VRNs88I0H8E=R<RR62oCCMsCN0
RRRRRRRRRRRRRRRRCIbjM_C5RH2<'=R4
';RRRRRRRRRRRRRRRRI4bC_5CMH<2R=4R''R;
RRRRRCRRMo8RCsMCNR0CW; 6
R
RRMRC8CRoMNCs0zCR4
c;
RRRRFbsO#C#Rp5Bi7,RQRh2LHCoMR
RRRRRRRHV5iBpR'=R4N'RMB8RpCi'P0CM2ER0CRM
RRRRRRRRRMRH_osC4=R<R_HMs;Co
RRRRRRRRRRRW) _ Rt4<W=R R;
RRRRRMRC8VRH;R
RRMRC8sRbF#OC#
;
RRRRzR.6:VRHRF5M0FR8ks0_CRo2oCCMsCN0
RRRRRRRR(z44b:RsCFO#5#RW) _ ,t4R7)q7R),W7q7)H,RMC_soR4,F_k0s2Co
RRRRRRRRoLCHRM
RRRRRRRRRHRRV5R5W) _ Rt4=4R''N2RM58R)7q7)RR=W7q7)R220MEC
RRRRRRRRRRRRRRRRz7ma=R<R_HMs4Co58IH04E-RI8FMR0Fj
2;RRRRRRRRRRRRCCD#
RRRRRRRRRRRRRRRRz7ma=R<R0Fk_osC58IH04E-RI8FMR0Fj
2;RRRRRRRRRRRRCRM8H
V;RRRRRRRRCRM8bOsFCR##z44(;R
RRMRC8CRoMNCs0zCR.
6;
RRRRjzdRRR:H5VR80Fk_osC2CRoMNCs0RC
RRRRRbRRsCFO#5#RmiBp,kRF0C_soL2RCMoH
RRRRRRRRRRRRRHV5pmBiRR='R4'NRM8miBp'CCPMR020MEC
RRRRRRRRRRRRRRRRz7ma=R<R0Fk_osC58IH04E-RI8FMR0Fj
2;RRRRRRRRRRRRCRM8H
V;RRRRRRRRCRM8bOsFC;##
RRRR8CMRMoCC0sNCdRzj
;
RRRR-t-RMNCs00CRE)CRqOvRC#DDR0IHEsR0H0-#N#0C
RRRR6z4RV:RFHsRRRHMM_klODCD#C_8C8bRF0IMFRRjoCCMsCN0
RRRRRRRR(z4RV:RF[sRRRHMM_klODCD#H_I88CRF0IMFRRjoCCMsCN0
RRRRRRRRRRRRqz)v7:RB. dX
cRRRRRRRRRRRRRRRRRb0FsRblNRQ57j>R=R_HMs5Co5c[*2R2,7RQ4=H>RMC_so[55*+c24R2,7RQ.=H>RMC_so[55*+c2.R2,7RQd=H>RMC_so[55*+c2d
2,RRRRRRRRRRRRRRRRRRRRRRRRRqRW7=jR>FRDIN_I858sjR2,W4q7RR=>D_FII8N8s254,qRW7=.R>FRDIN_I858s.R2,Wdq7RR=>D_FII8N8s25d,qRW7=cR>FRDIN_I858sc
2,RRRRRRRRRRRRRRRRRRRRRRRRRqR)7=jR>FRDIN_s858sjR2,)4q7RR=>D_FIs8N8s254,qR)7=.R>FRDIN_s858s.R2,)dq7RR=>D_FIs8N8s25d,qR)7=cR>FRDIN_s858sc
2,-R-RRRRRRRRRRRRRRRRRRRRRRRRRWh) RR=>WR ,Wju RR=>IjbC_5CMHR2,W4u RR=>I4bC_5CMHR2,B=iR>mRhap5BiR2,
RRRRRRRRRRRRRRRRRRRRRRRRWRR)R h=W>R W,RuR j=I>Rb_CjCHM52W,RuR 4=I>Rb_C4CHM52B,Ri>R=RiBp,RR
RRRRRRRRRRRRRRRRRRRRRRRRRj7mRR=>F_k0L5k#H[,5*2c2,mR74>R=R0Fk_#Lk55H,[2*c+,42R.7mRR=>F_k0L5k#H[,5*+c2.R2,7Rmd=F>RkL0_kH#5,*5[cd2+2
2;RRRRRRRRRRRRRRRRF_k0s5Co5c[*2<2R=kRF0k_L#,5H5c[*2I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co5c[*22+4RR<=F_k0L5k#H[,5*+c24I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co5c[*22+.RR<=F_k0L5k#H[,5*+c2.I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co5c[*22+dRR<=F_k0L5k#H[,5*+c2dI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRCRM8oCCMsCN0R(z4;R
RRMRC8CRoMNCs0zCR4
6;
R--RUz.RH:RV8R5F_k0s2CoRMoCC0sNC-
-RRRRRRRRzR4n:FRVsRRHHMMRkOl_C#DD_C8CbFR8IFM0RojRCsMCN
0C-R-RRRRRR4RzURR:VRFs[MRHRlMk_DOCDI#_HR8C8MFI0jFRRMoCC0sNC-
-RRRRRRRRRRRRzv)q:BR7 Xd.c-R
-RRRRRRRRRRRRRRRRsbF0NRlb7R5Q=jR>MRH_osC5*5[c,22R47QRR=>HsM_C5o5[2*c+,42R.7QRR=>HsM_C5o5[2*c+,.2Rd7QRR=>HsM_C5o5[2*c+,d2
R--RRRRRRRRRRRRRRRRRRRRRRRRR7Wqj>R=RIDF_8IN8js52W,RqR74=D>RFII_Ns885,42R7Wq.>R=RIDF_8IN8.s52W,RqR7d=D>RFII_Ns885,d2R7Wqc>R=RIDF_8IN8cs52-,
-RRRRRRRRRRRRRRRRRRRRRRRR)RRqR7j=D>RFsI_Ns885,j2R7)q4>R=RIDF_8sN84s52),RqR7.=D>RFsI_Ns885,.2R7)qd>R=RIDF_8sN8ds52),RqR7c=D>RFsI_Ns885,c2
R--RRRRRRRRRRRRRRRRRRRRRRRRR W)h>R=R,W R Wuj>R=RCIbjM_C5,H2R Wu4>R=RCIb4M_C5,H2RRBi=h>RmBa5p,i2R-
-RRRRRRRRRRRRRRRRRRRRRRRRR7RTm=jR>kRF0k_L#,5H5c[*2R2,T47mRR=>F_k0L5k#H[,5*+c24R2,T.7mRR=>F_k0L5k#H[,5*+c2.R2,Td7mRR=>F_k0L5k#H[,5*+c2d;22

---R-RRRRRRRRRRRRRF_k0s5Co5c[*2<2R=kRF0k_L#,5H5c[*2I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';-R-RRRRRRRRRRRRRRkRF0C_so[55*+c24<2R=kRF0k_L#,5H5c[*22+4RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;-
-RRRRRRRRRRRRRRRRF_k0s5Co5c[*22+.RR<=F_k0L5k#H[,5*+c2.I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';-R-RRRRRRRRRRRRRRkRF0C_so[55*+c2d<2R=kRF0k_L#,5H5c[*22+dRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;-
-RRRRRRRRRRRRCRM8oCCMsCN0RUz4;-
-RRRRRCRRMo8RCsMCNR0Cz;4n
R--RCRRMo8RCsMCNR0Cz;.U
-
-RRRRRURkRH:RV8R5F_k0s2CoRMoCC0sNC-
-RRRRRmR7z<aR=kRF0C_soH5I8-0E4FR8IFM0R;j2
R--R8CMRMoCC0sNCURk;R
RRRRRRCR
MN8RsHOE00COkRsCNEsOj
;

