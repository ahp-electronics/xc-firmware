--------------------------------------------------
@ES--a1m_am7ptRQBVOkM0MHFRObN	CNo
------------------------------------------------
--
LDHs$NsSCHCCk;
#HCRC3CC#_08DHFoO4_4nNc3D
D;
ObN	CNoS8#0_oDFH1O_AHaR#R

RwRRzahBQRmha1F_0F8poRHORRRRRRR5LRR:ARQaRRRRRRRRRRRRRRR2)z a)#hR0D8_FOoH;R
RRCR
M#8R0D8_FOoH_a1A;b

NNO	oLCRFR8$#_08DHFoOA_1a#RH
-
------------------------------------------------------------------R-
RwRRzahBQRmha1F_0F8poRHORRRRRRR5LRR:ARQaRRRRRRRRRRRRRRR2)z a)#hR0D8_FOoHR
Q1RRRRAQ thR
RRRRRRqRB1L RR
Q1RRRRRRRRRRRRWh] R''jRR=>)z a)'hRj
';RRRRRRRRRRRRWh] R''4RR=>)z a)'hR4
';RRRRRRRR Rh7B q1;R
RRhR 7
;
CRM8#_08DHFoOA_1a
;

=--=========================================================================
==-1-RAq_B)R)Y
=--=========================================================================
==
R
RRHRDLssN$CRHC
C;RRRRkR#CHCCC38#0_oDFH4O_43ncN;DD
RRRRCk#RCHCC03#8F_Do_HOkHM#o8MC3DND;R
RRRR
R
RRCHM001$RAq_B)R)YHu#
FRs05QRRjRR:HRMR#_08DHFoOR;
RRRRRQRR4RR:HRMR#_08DHFoOR;
RRRRRBRRQRR:HRMR#_08DHFoOR;
RRRRRBRRmRR:FRk0R8#0_oDFHROR2C;
M18RAq_B);)Y
0N0skHL0#CR$LM_D	NO_GLFRRFV1BA_qY))RO:RFFlbM0CMRRH#0Csk;N

sHOE00COkRsCVOkMRRFV1BA_qY))R
H##MHoNBDRQM_H0#R:0D8_FOoH:j=''L;
CMoH
FbsO#C#52BQ
CSLoRHM
RSRRRHV5RBQ=4R'')RmRRBQ=jR''02RERCMBHQ_M=0<B
Q;SRRRCCD#R_BQH<M0=jR''S;
RCRRMH8RVR;
R8CMRFbsO#C#;B

m=R<RQ5B_0HMR8NMR2QjRRFs5_BQHRM0NRM8QR42F5sRQNjRMQ8R4
2;RM
C8kRVMRO;
-

-============================================================================-
-R_1AB)q)Yh_Q_XvzR-
-============================================================================
R
RRHRDLssN$CRHC
C;RRRRkR#CHCCC38#0_oDFH4O_43ncN;DD
RRRRCk#RCHCC03#8F_Do_HOkHM#o8MC3DND;C

M00H$AR1_)Bq)QY_hz_vX#RH
MoCCOsH5QB_h:QaL_H0P0COF4s5RI8FMR0Fj:2R=jR"j;"2
RRRRsbF0RR5
RSROsNs$M_HHF0_kR0R:kRF0#RR0D8_FOoH;R
SRsONsH$_M_H0HRMR:MRHR0R#8F_DoRHOR;R2
M
C8AR1_)Bq)QY_hz_vX
;RNs00H0LkC$R#MD_LN_O	LRFGF1VRAq_B)_)YQvh_z:XRRlOFbCFMMH0R#sR0k
C;Rs
NO0EHCkO0sVCRkRMOF1VRAq_B)_)YQvh_zHXR#H
#oDMNRD#CC_O0L#H0R0:#8F_Do_HOP0COF4s5RI8FMR0Fj
2;
oLCHbM
sCFO###5CODC0H_L0O#,N$ss_HHM0M_H2L
SCMoHRR
SR#ONCCR#D0CO_0LH##RH
RSRRIRRERCM""jj=N>Os_s$H0MH_0Fk<j=''S;
RRRRRCIEMjR"4>"=OsNs$M_HHF0_k=0<';4'
RSRRIRRERCM""4j=N>Os_s$H0MH_0Fk<N=Os_s$H0MH_;HM
RSRRIRRERCM""44=N>Os_s$H0MH_0Fk<N=Os_s$H0MH_;HM
RSRRIRRERCMFC0Es=#R>sONsH$_M_H0F<k0=''j;R
SR8CMR#ONCS;
RRRR
RRRCRM8bOsFC;##
RRR#CCDOL0_HR0#<a=Rma_17tpmQ BeB)am5QB_h2Qa;

RCRM8VOkM;
R
-=-==========================================================================-=
-AR1_apzc-R
-============================================================================R

RDRRHNLssH$RC;CC
RRRRCk#RCHCC03#8F_Do_HO4c4n3DND;R
RR#RkCCRHC#C30D8_FOoH_#kMHCoM8D3NDR;
R
RRCHM001$RAz_paHcR#R
RRMoCCOsH5apz_QQhaH:L0C_POs0F5R468MFI0jFR2=R:Rj"jjjjjjjjjjjjjj2j";R
RRsbF0RR5
RSRm:RRR0FkR0R#8F_Do;HO
RSRQRjR:MRHR0R#8F_Do;HO
RSRQR4R:MRHR0R#8F_Do;HO
RSRQR.R:MRHR0R#8F_Do;HO
RSRQRdR:MRHR0R#8F_DoRHOR;R2
M
C8AR1_apzc
;RNs00H0LkC$R#MD_LN_O	LRFGF1VRAz_pa:cRRlOFbCFMMH0R#sR0k
C;Rs
NO0EHCkO0sVCRkRMOF1VRAz_paHcR#H
#oDMNR#lN	#R:0D8_FOoH_OPC05Fs486RF0IMF2Rj;H
#oDMNR0Dk#0:#8F_Do:HO=''j;H
#oDMNR_QdH#M:0D8_FOoH:j=''#;
HNoMD.RQ_:HM#_08DHFoO':=j
';#MHoNQDR4M_H:8#0_oDFH=O:';j'
o#HMRNDQHj_M0:#8F_Do:HO=''j;H
#oDMNRuQhz:a1#_08DHFoOC_POs0F58dRF0IMF2Rj;C
Lo
HM
s
bF#OC#d5Q_,HMQH._M4,Q_,HMQHj_MS2
LHCoMRR
RRRRRRRRR_QdH<MR=dRQ;R
RRRRRRRRRQH._M=R<R;Q.
RRRRRRRRQRR4M_HRR<=Q
4;RRRRRRRRRjRQ_RHM<Q=RjS;
RRRRRNRl#<	R=mRa_71apQmtBBe a5m)p_zaQahQ2R;
RRRRRRRRmD<=k;0#
RSRRRRRRuQhz<a1=_QdH&MRR_Q.H&MRR_Q4H&MRR_QjH
M;SR
SRNRO#QCRhauz1#RH
RSRRIRRERCM"jjjj>"=D#k0<l=RN5#	jV2N0RCsj43jR;M#
RSRRIRRERCM"jjj4>"=D#k0<l=RN5#	4V2N0RCsj43jR;M#
RSRRIRRERCM"4jjj>"=D#k0<l=RN5#	.V2N0RCsj43jR;M#
RSRRIRRERCM"4jj4>"=D#k0<l=RN5#	dV2N0RCsj43jR;M#
RSRRIRRERCM"jj4j>"=D#k0<l=RN5#	cV2N0RCsj43jR;M#
RSRRIRRERCM"jj44>"=D#k0<l=RN5#	6V2N0RCsj43jR;M#
RSRRIRRERCM"4j4j>"=D#k0<l=RN5#	nV2N0RCsj43jR;M#
RSRRIRRERCM"4j44>"=D#k0<l=RN5#	(V2N0RCsj43jR;M#
RSSRERIC"MR4jjj"D=>k<0#=NRl#U	520NVCjsR3Rj4M
#;SRRRRERIC"MR44jj"D=>k<0#=NRl#g	520NVCjsR3Rj4M
#;SRRRRERIC"MR4jj4"D=>k<0#=NRl#4	5jV2N0RCsj43jR;M#
RSRRIRRERCM"44j4>"=D#k0<l=RN5#	4N42Vs0CRjj34#RM;R
SRRRRIMECR4"4j=j">0Dk#R<=l	N#524.NCV0s3RjjM4R#S;
RRRRRCIEM4R"4"j4=k>D0=#<R#lN	d5420NVCjsR3Rj4M
#;SRRRRERIC"MR4j44"D=>k<0#=NRl#4	5cV2N0RCsj43jR;M#
RSRRIRRERCM"4444>"=D#k0<l=RN5#	4N62Vs0CRjj34#RM;R
SRRRRIMECREF0C=s#>0Dk#R<=l	N#5Nj2Vs0CRjj34#RM;R
SRMRC8NRO#
C;RMRC8sRbF#OC#
;RCRM8VOkM;


-=-==========================================================================-=
-AR1_w7wR-
-============================================================================
R
RRHRDLssN$CRHC
C;RRRRkR#CHCCC38#0_oDFH4O_43ncN;DD
RRRRCk#RCHCC03#8F_Do_HOkHM#o8MC3DND;C

M00H$AR1_w7wR
H#RbRRFRs05SR
RRRTRF:RkR0R#_08DHFoOS;
RRR7RH:RM#RR0D8_FOoH;R
SRRBR:MRHR0R#8F_DoRHOR
2;S
RRCRM817A_wRw;
0N0skHL0#CR$LM_D	NO_GLFRRFV17A_w:wRRlOFbCFMMH0R#sR0k
C;Rs
NO0EHCkO0sVCRkRMOF1VRAw_7w#RH
oLCHRM
bOsFC5##BR2
RCRLo
HMSHRRV'RBCMPC0MRN8RRB=4R''ER0CSM
SRRT<7=R;R
RRRRRCRM8H
V;RCRRMb8RsCFO#
#;CRM8RMVkO
;

=--=========================================================================
==-1-RAw_7wR1)
=--=========================================================================
==
RRRRLDHs$NsRCHCCR;
RkRR#HCRC3CC#_08DHFoO4_4nNc3D
D;RRRRkR#CHCCC38#0_oDFHkO_Mo#HM3C8N;DD
M
C0$H0R_1A71ww)#RH
RRRb0FsR
5RRRRR):RRRRHMR8#0_oDFH
O;STRRRRR:FRk0R8#0_oDFH
O;S7RRRRR:HRMR#_08DHFoOS;
RRRBRH:RM#RR0D8_FOoHR;R2
RSR
8CMR_1A71ww)
;RNs00H0LkC$R#MD_LN_O	LRFGF1VRAw_7wR1):FROlMbFCRM0H0#Rs;kC
NR
sHOE00COkRsCVOkMRRFV17A_w)w1R
H#LHCoMb
RsCFO#B#52R
RRoLCHSM
RVRHRCB'P0CMR8NMR=BRR''4RC0EMR
SRRRRH)VRR'=R4E'0CSM
SRRRRRRRR<TR=jR''S;
SRRRCCD#
RSSRRRRRTRRRR<=7R;
RRRRRMRC8VRH;R
RRMRC8VRH;R
RR8CMRFbsO#C#;M
C8VRRk;MO
-

-============================================================================-
-R_1A71ww1-R
-============================================================================R

RDRRHNLssH$RC;CC
RRRRCk#RCHCC03#8F_Do_HO4c4n3DND;R
RR#RkCCRHC#C30D8_FOoH_#kMHCoM8D3ND
;
CHM001$RAw_7wR11HR#
RFRbs50RRR
RRRR1RH:RM#RR0D8_FOoH;R
SRRTR:kRF0#RR0D8_FOoH;R
SRR7R:MRHR0R#8F_Do;HO
RSRB:RRRRHMR8#0_oDFHROR2S;
RCR
M18RAw_7w;11R0
N0LsHkR0C#_$MLODN	F_LGVRFR_1A71ww1RR:ObFlFMMC0#RHRk0sCR;

ONsECH0Os0kCkRVMFORVAR1_w7w1H1R#C
Lo
HMRFbsO#C#5
B2RLRRCMoH
RSRHBVR'CCPMN0RMB8RR'=R40'RE
CMSRRRRVRHR=1RR''40MEC
RSSRRRRRTRRRR<=';4'
RSSRDRC#SC
SRRRRRRRR<TR=;R7
RRRRRRRCRM8H
V;RRRRCRM8H
V;RCRRMb8RsCFO#
#;CRM8RMVkO
;

-
-============================================================================
R--17A_wRw)
=--=========================================================================
==
RRRRLDHs$NsRCHCCR;
RkRR#HCRC3CC#_08DHFoO4_4nNc3D
D;RRRRkR#CHCCC38#0_oDFHkO_Mo#HM3C8N;DD
C

M00H$AR1_w7w)#RH
RRRb0FsR
5RRRRR):RRRRHMR8#0_oDFH
O;STRRRRR:FRk0R8#0_oDFH
O;S7RRRRR:HRMR#_08DHFoOS;
RRRBRH:RM#RR0D8_FOoHR;R2
RSR
8CMR_1A7)ww;NR
0H0sLCk0RM#$_NLDOL	_FFGRVAR1_w7w)RR:ObFlFMMC0#RHRk0sCR;

ONsECH0Os0kCkRVMFORVAR1_w7w)#RH
oLCHRM
bOsFC5##BRR,)
R2RLRRCMoH
RSRH5VRBP'CCRM0NRM8BRR='24'RRm)5C)'P0CMR8NMR=)RR''420RRE
CMSRRRRVRHR=)RR''40MEC
RSSRRRRRTRRRR<=';j'
RSSRDRC#SC
SRRRRRRRR<TR=;R7
RRRRRRRCRM8H
V;RRRRCRM8H
V;RCRRMb8RsCFO#
#;CRM8RMVkO
;

=--=========================================================================
==-1-RAw_7w
1R-=-==========================================================================
=
RRRRDsHLNRs$HCCC;R
RR#RkCCRHC#C30D8_FOoH_n44cD3NDR;
RkRR#HCRC3CC#_08DHFoOM_k#MHoCN83D
D;
0CMHR0$17A_wRw1HR#
RFRbs50RRR
RRRR1RH:RM#RR0D8_FOoH;R
SRRTR:kRF0#RR0D8_FOoH;R
SRR7R:MRHR0R#8F_Do;HO
RSRB:RRRRHMR8#0_oDFHROR2S;
RCR
M18RAw_7wR1;
0N0skHL0#CR$LM_D	NO_GLFRRFV17A_wRw1:FROlMbFCRM0H0#Rs;kC
NR
sHOE00COkRsCVOkMRRFV17A_wRw1HL#
CMoH
sRbF#OC#R5B,RR12R
RRoLCHSM
RVRHR'5BCMPC0MRN8RRB=4R''m2R)1R5'CCPMN0RM18RR'=R4R'2RC0EMR
SRRRRH1VRR'=R4E'0CSM
SRRRRRRRR<TR=4R''S;
SRRRCCD#
RSSRRRRRTRRRR<=7R;
RRRRRMRC8VRH;R
RRMRC8VRH;R
RR8CMRFbsO#C#;M
C8VRRk;MO
-

-============================================================================-
-R_1A7 wwR-
-============================================================================
R
RRHRDLssN$CRHC
C;RRRRkR#CHCCC38#0_oDFH4O_43ncN;DD
RRRRCk#RCHCC03#8F_Do_HOkHM#o8MC3DND;


CHM001$RAw_7wH R#R
RRsbF0RR5
RRRRR R:MRHR0R#8F_DoRHO:'=R]
';STRRRRR:FRk0R8#0_oDFH
O;S7RRRRR:HRMR#_08DHFoOS;
RRRBRH:RM#RR0D8_FOoHR;R2
RSR
8CMR_1A7 ww;NR
0H0sLCk0RM#$_NLDOL	_FFGRVAR1_w7w RR:ObFlFMMC0#RHRk0sCR;

ONsECH0Os0kCkRVMFORVAR1_w7w #RH
oLCHRM
bOsFC5##BR2
RCRLo
HMSHRRV'RBCMPC0MRN8RRB=4R''0RRE
CMSRRRRVRHR= RR''40MEC
RSSRRRRRTRRRR<=7S;
SRRRCRM8H
V;RRRRCRM8H
V;RCRRMb8RsCFO#
#;CRM8RMVkO
;

=--=========================================================================
==-1-RAw_7w) 1R-
-============================================================================
R
RRHRDLssN$CRHC
C;RRRRkR#CHCCC38#0_oDFH4O_43ncN;DD
RRRRCk#RCHCC03#8F_Do_HOkHM#o8MC3DND;


CHM001$RAw_7w) 1R
H#RbRRFRs05RR
R RRRRR:HRMR#_08DHFoO=R:R''];R
RRRR)RH:RM#RR0D8_FOoH;R
SRRTR:kRF0#RR0D8_FOoH;R
SRR7R:MRHR0R#8F_Do;HO
RSRB:RRRRHMR8#0_oDFHROR2S;
RCR
M18RAw_7w) 1;NR
0H0sLCk0RM#$_NLDOL	_FFGRVAR1_w7w R1):FROlMbFCRM0H0#Rs;kC
NR
sHOE00COkRsCVOkMRRFV17A_w1w )#RH
oLCHRM
bOsFC5##BR2
RCRLo
HMSHRRV'RBCMPC0MRN8RRB=4R''ER0CSM
RRRRH VRR'=R40'RERCMRR
SRRRRRVRHR=)RR''40MEC
RSSRRRRRRRRR<TR=jR''S;
SRRRRDRC#SC
SRRRRRRRRTRRRR<=7R;
RRRRRMRC8VRH;R
RRRRRCRM8H
V;RRRRCRM8H
V;RCRRMb8RsCFO#
#;CRM8RMVkO
;

=--=========================================================================
==-1-RAw_7w1 1R-
-============================================================================
R
RRHRDLssN$CRHC
C;RRRRkR#CHCCC38#0_oDFH4O_43ncN;DD
RRRRCk#RCHCC03#8F_Do_HOkHM#o8MC3DND;


CHM001$RAw_7w1 1R
H#RbRRFRs05RR
R RRRRR:HRMR#_08DHFoO=R:R''];R
RRRR1RH:RM#RR0D8_FOoH;R
SRRTR:kRF0#RR0D8_FOoH;R
SRR7R:MRHR0R#8F_Do;HO
RSRB:RRRRHMR8#0_oDFHROR2S;
RCR
M18RAw_7w1 1;NR
0H0sLCk0RM#$_NLDOL	_FFGRVAR1_w7w R11:FROlMbFCRM0H0#Rs;kC
NR
sHOE00COkRsCVOkMRRFV17A_w1w 1#RH
oLCHRM
bOsFC5##BR2
RCRLo
HMSHRRV'RBCMPC0MRN8RRB=4R''ER0CSM
RRRRH VRR'=R40'RERCMRR
SRRRRRVRHR=1RR''40MEC
RSSRRRRRRRRR<TR=4R''S;
SRRRRDRC#SC
SRRRRRRRRTRRRR<=7R;
RRRRRMRC8VRH;R
RRRRRCRM8H
V;RRRRCRM8H
V;RCRRMb8RsCFO#
#;CRM8RMVkO
;

=--=========================================================================
==-1-RAw_7wR )
=--=========================================================================
==
RRRRLDHs$NsRCHCCR;
RkRR#HCRC3CC#_08DHFoO4_4nNc3D
D;RRRRkR#CHCCC38#0_oDFHkO_Mo#HM3C8N;DD
C

M00H$AR1_w7w H)R#R
RRsbF0RR5
RRRRR R:MRHR0R#8F_DoRHO:'=R]
';RRRR):RRRRHMR8#0_oDFH
O;STRRRRR:FRk0R8#0_oDFH
O;S7RRRRR:HRMR#_08DHFoOS;
RRRBRH:RM#RR0D8_FOoHR;R2
RSR
8CMR_1A7 ww)
;RNs00H0LkC$R#MD_LN_O	LRFGF1VRAw_7wR ):FROlMbFCRM0H0#Rs;kC
NR
sHOE00COkRsCVOkMRRFV17A_w)w R
H#LHCoMb
RsCFO#B#5R),RRR2
RCRLo
HMSHRRVBR5'CCPMN0RMB8RR'=R4R'2m5)R)P'CCRM0NRM8)RR='24'RER0CSM
RRRRH VRR'=R40'RERCMRR
SRRRRRVRHR=)RR''40MEC
RSSRRRRRRRRR<TR=jR''S;
SRRRRDRC#SC
SRRRRRRRRTRRRR<=7R;
RRRRRRRRCRM8H
V;RRRRRMRC8VRH;R
RRMRC8VRH;R
RR8CMRFbsO#C#;M
C8VRRk;MO
-

-============================================================================-
-R_1A7 ww1-R
-============================================================================R

RDRRHNLssH$RC;CC
RRRRCk#RCHCC03#8F_Do_HO4c4n3DND;R
RR#RkCCRHC#C30D8_FOoH_#kMHCoM8D3ND
;
CHM001$RAw_7wR 1HR#
RFRbs50RRR
RRRR RH:RM#RR0D8_FOoHRR:=';]'
RRRRR1R:MRHR0R#8F_Do;HO
RSRT:RRR0FkR0R#8F_Do;HO
RSR7:RRRRHMR8#0_oDFH
O;SBRRRRR:HRMR#_08DHFoO2RR;R
SRM
C8AR1_w7w R1;
0N0skHL0#CR$LM_D	NO_GLFRRFV17A_w1w RO:RFFlbM0CMRRH#0Csk;

RNEsOHO0C0CksRMVkOVRFR_1A7 ww1#RH
oLCHRM
bOsFC5##BRR,1R2
RCRLo
HMSHRRVBR5'CCPMN0RMB8RR'=R4R'2m5)R1P'CCRM0NRM81RR='24'RER0CSM
RRRRH VRR'=R40'RERCMRR
SRRRRRVRHR=1RR''40MEC
RSSRRRRRRRRR<TR=4R''S;
SRRRRDRC#SC
SRRRRRRRRTRRRR<=7R;
RRRRRRRRCRM8H
V;RRRRRMRC8VRH;R
RRMRC8VRH;R
RR8CMRFbsO#C#;M
C8VRRk;MO
-

-============================================================================-
-R_1A7hwwR-
-============================================================================
R
RRHRDLssN$CRHC
C;RRRRkR#CHCCC38#0_oDFH4O_43ncN;DD
RRRRCk#RCHCC03#8F_Do_HOkHM#o8MC3DND;C

M00H$AR1_w7wh#RH
RRRb0FsR
5RSTRRRRR:FRk0R8#0_oDFH
O;S7RRRRR:HRMR#_08DHFoOS;
RRRBRH:RM#RR0D8_FOoHR;R2
RSR
8CMR_1A7hww;NR
0H0sLCk0RM#$_NLDOL	_FFGRVAR1_w7whRR:ObFlFMMC0#RHRk0sCR;

ONsECH0Os0kCkRVMFORVAR1_w7wh#RH
oLCHRM
bOsFC5##BR2
RCRLo
HMSHRRV'RBCMPC0MRN8RRB=jR''ER0CSM
SRRT<7=R;R
RRRRRCRM8H
V;RCRRMb8RsCFO#
#;CRM8RMVkO
;

=--=========================================================================
==-1-RAw_7w)h1R-
-============================================================================
R
RRHRDLssN$CRHC
C;RRRRkR#CHCCC38#0_oDFH4O_43ncN;DD
RRRRCk#RCHCC03#8F_Do_HOkHM#o8MC3DND;C

M00H$AR1_w7whR1)HR#
RFRbs50RRR
RRRR)RH:RM#RR0D8_FOoH;R
SRRTR:kRF0#RR0D8_FOoH;R
SRR7R:MRHR0R#8F_Do;HO
RSRB:RRRRHMR8#0_oDFHROR2S;
RCR
M18RAw_7w)h1;NR
0H0sLCk0RM#$_NLDOL	_FFGRVAR1_w7whR1):FROlMbFCRM0H0#Rs;kC
NR
sHOE00COkRsCVOkMRRFV17A_w1wh)#RH
oLCHRM
bOsFC5##BR2
RCRLo
HMSHRRV'RBCMPC0MRN8RRB=jR''ER0CSM
RRRRRRHV)RR='04'E
CMSRSRRRRRRRRT<'=Rj
';SRSRR#CDCS
SRRRRRRRRT=R<R
7;RRRRRCRRMH8RVR;
RCRRMH8RVR;
RMRC8sRbF#OC#C;
MR8RVOkM;



=--=========================================================================
==-1-RAw_7w1h1R-
-============================================================================
R
RRHRDLssN$CRHC
C;RRRRkR#CHCCC38#0_oDFH4O_43ncN;DD
RRRRCk#RCHCC03#8F_Do_HOkHM#o8MC3DND;S

CHM001$RAw_7w1h1R
H#SRRRb0FsR
5RSRRRRR1R:MRHR0R#8F_Do;HO
RSSRRTR:kRF0#RR0D8_FOoH;S
SRRR7RH:RM#RR0D8_FOoH;S
SRRRBRH:RM#RR0D8_FOoHR;R2
RSSRC
SM18RAw_7w1h1;SR
Ns00H0LkC$R#MD_LN_O	LRFGF1VRAw_7w1h1RO:RFFlbM0CMRRH#0Csk;R
S
sSNO0EHCkO0sVCRkRMOF1VRAw_7w1h1R
H#SoLCHSM
RFbsO#C#5
B2SRRRLHCoMS
SRVRHRCB'P0CMR8NMR=BRR''jRC0EMS
SRRRRRRHV1RR='04'E
CMSRSSRRRRRTRRRR<=';4'
SSSRCRRD
#CSRSSRRRRRTRRRR<=7S;
RRRRRCRRMH8RVS;
RRRRCRM8H
V;SRRRCRM8bOsFC;##
MSC8VRRk;MO

S
-=-==========================================================================-=
-AR1_w7wh
)R-=-==========================================================================
=
RRRRDsHLNRs$HCCC;R
RR#RkCCRHC#C30D8_FOoH_n44cD3NDR;
RkRR#HCRC3CC#_08DHFoOM_k#MHoCN83D
D;
0CMHR0$17A_w)whR
H#RbRRFRs05RR
R)RRRRR:HRMR#_08DHFoOS;
RRRTRF:RkR0R#_08DHFoOS;
RRR7RH:RM#RR0D8_FOoH;R
SRRBR:MRHR0R#8F_DoRHOR
2;S
RRCRM817A_w)wh;NR
0H0sLCk0RM#$_NLDOL	_FFGRVAR1_w7wh:)RRlOFbCFMMH0R#sR0k
C;Rs
NO0EHCkO0sVCRkRMOF1VRAw_7wRh)HL#
CMoH
sRbF#OC#R5B,RR)2R
RRoLCHSM
RVRHR'5BCMPC0MRN8RRB=jR''m2R))R5'CCPMN0RM)8RR'=R4R'2RC0EMR
SRRRRH)VRR'=R4E'0CSM
SRRRRRRRR<TR=jR''S;
SRRRCCD#
RSSRRRRRTRRRR<=7R;
RRRRRMRC8VRH;R
RRMRC8VRH;R
RR8CMRFbsO#C#;M
C8VRRk;MO
-

-============================================================================-
-R_1A7hww1-R
-============================================================================R

RDRRHNLssH$RC;CC
RRRRCk#RCHCC03#8F_Do_HO4c4n3DND;R
RR#RkCCRHC#C30D8_FOoH_#kMHCoM8D3ND
;

0CMHR0$17A_w1whR
H#RbRRFRs05RR
R1RRRRR:HRMR#_08DHFoOS;
RRRTRF:RkR0R#_08DHFoOS;
RRR7RH:RM#RR0D8_FOoH;R
SRRBR:MRHR0R#8F_DoRHOR
2;S
RRCRM817A_w1wh;NR
0H0sLCk0RM#$_NLDOL	_FFGRVAR1_w7wh:1RRlOFbCFMMH0R#sR0k
C;Rs
NO0EHCkO0sVCRkRMOF1VRAw_7wRh1HL#
CMoH
sRbF#OC#R5B,RR12R
RRoLCHSM
RVRHR'5BCMPC0MRN8RRB=jR''m2R)1R5'CCPMN0RM18RR'=R4R'2RC0EMR
SRRRRH1VRR'=R4E'0CSM
SRRRRRRRR<TR=4R''S;
SRRRCCD#
RSSRRRRRTRRRR<=7R;
RRRRRMRC8VRH;R
RRMRC8VRH;R
RR8CMRFbsO#C#;M
C8VRRk;MO
-

-============================================================================-
-R_1A7hww -R
-============================================================================R

RDRRHNLssH$RC;CC
RRRRCk#RCHCC03#8F_Do_HO4c4n3DND;R
RR#RkCCRHC#C30D8_FOoH_#kMHCoM8D3ND
;

0CMHR0$17A_w whR
H#RbRRFRs05RR
R RRRRR:HRMR#_08DHFoO=R:R''];R
SRRTR:kRF0#RR0D8_FOoH;R
SRR7R:MRHR0R#8F_Do;HO
RSRB:RRRRHMR8#0_oDFHROR2S;
RCR
M18RAw_7w;h R0
N0LsHkR0C#_$MLODN	F_LGVRFR_1A7hww RR:ObFlFMMC0#RHRk0sCR;

ONsECH0Os0kCkRVMFORVAR1_w7whH R#C
Lo
HMRFbsO#C#5
B2RLRRCMoH
RSRHBVR'CCPMN0RMB8RR'=RjR'R0MEC
RSRRHRRVRR =4R''C0EMS
SRRRRRRRRT=R<R
7;SRSRR8CMR;HV
RRRR8CMR;HV
RRRCRM8bOsFC;##
8CMRkRVM
O;
-
-============================================================================
R--17A_w wh1
)R-=-==========================================================================
=
RRRRDsHLNRs$HCCC;R
RR#RkCCRHC#C30D8_FOoH_n44cD3NDR;
RkRR#HCRC3CC#_08DHFoOM_k#MHoCN83D
D;
M
C0$H0R_1A7hww R1)HR#
RFRbs50RRR
RRRR RH:RM#RR0D8_FOoHRR:=';]'
RRRRR)R:MRHR0R#8F_Do;HO
RSRT:RRR0FkR0R#8F_Do;HO
RSR7:RRRRHMR8#0_oDFH
O;SBRRRRR:HRMR#_08DHFoO2RR;R
SRM
C8AR1_w7wh) 1;NR
0H0sLCk0RM#$_NLDOL	_FFGRVAR1_w7wh) 1RO:RFFlbM0CMRRH#0Csk;

RNEsOHO0C0CksRMVkOVRFR_1A7hww R1)HL#
CMoH
sRbF#OC#25B
RRRLHCoMR
SRRHVBP'CCRM0NRM8BRR='Rj'0MEC
RSRRVRHR= RR''4RC0EM
RRSRRRRRRRH)VRR'=R4E'0CSM
SRRRRRRRRTRRRR<=';j'
RSSRRRRCCD#
RSSRRRRRRRRR<TR=;R7
RRRRRRRCRM8H
V;RRRRRMRC8VRH;R
RRMRC8VRH;R
RR8CMRFbsO#C#;M
C8VRRk;MO
-

-============================================================================-
-R_1A7hww R11
=--=========================================================================
==
RRRRLDHs$NsRCHCCR;
RkRR#HCRC3CC#_08DHFoO4_4nNc3D
D;RRRRkR#CHCCC38#0_oDFHkO_Mo#HM3C8N;DD



CHM001$RAw_7w1h 1#RH
RRRb0FsR
5RRRRR :RRRRHMR8#0_oDFH:OR=]R''R;
R1RRRRR:HRMR#_08DHFoOS;
RRRTRF:RkR0R#_08DHFoOS;
RRR7RH:RM#RR0D8_FOoH;R
SRRBR:MRHR0R#8F_DoRHOR
2;S
RRCRM817A_w wh1R1;
0N0skHL0#CR$LM_D	NO_GLFRRFV17A_w wh1:1RRlOFbCFMMH0R#sR0k
C;Rs
NO0EHCkO0sVCRkRMOF1VRAw_7w1h 1#RH
oLCHRM
bOsFC5##BR2
RCRLo
HMSHRRV'RBCMPC0MRN8RRB=jR''ER0CSM
RRRRH VRR'=R40'RERCMRR
SRRRRRVRHR=1RR''40MEC
RSSRRRRRRRRR<TR=4R''S;
SRRRRDRC#SC
SRRRRRRRRTRRRR<=7R;
RRRRRMRC8VRH;R
RRRRRCRM8H
V;RRRRCRM8H
V;RCRRMb8RsCFO#
#;CRM8RMVkO
;

=--=========================================================================
==-1-RAw_7w)h R-
-============================================================================
R
RRHRDLssN$CRHC
C;RRRRkR#CHCCC38#0_oDFH4O_43ncN;DD
RRRRCk#RCHCC03#8F_Do_HOkHM#o8MC3DND;


CHM001$RAw_7w)h R
H#RbRRFRs05RR
R RRRRR:HRMR#_08DHFoO=R:R''];R
RRRR)RH:RM#RR0D8_FOoH;R
SRRTR:kRF0#RR0D8_FOoH;R
SRR7R:MRHR0R#8F_Do;HO
RSRB:RRRRHMR8#0_oDFHROR2S;
RCR
M18RAw_7w)h ;NR
0H0sLCk0RM#$_NLDOL	_FFGRVAR1_w7whR ):FROlMbFCRM0H0#Rs;kC
NR
sHOE00COkRsCVOkMRRFV17A_w wh)#RH
oLCHRM
bOsFC5##BRR,)
R2RLRRCMoH
RSRH5VRBP'CCRM0NRM8BRR='2j'RRm)5C)'P0CMR8NMR=)RR''420RRE
CMSRRRRRHV RR='R4'0MECRSR
RRRRRHRRVRR)=4R''C0EMS
SRRRRRRRRRRRT<'=Rj
';SRSRRCRRD
#CSRSRRRRRRRRRT=R<R
7;RRRRRRRRR8CMR;HV
RRRRCRRMH8RVR;
RCRRMH8RVR;
RMRC8sRbF#OC#C;
MR8RVOkM;


-=-==========================================================================-=
-AR1_w7whR 1
=--=========================================================================
==
RRRRLDHs$NsRCHCCR;
RkRR#HCRC3CC#_08DHFoO4_4nNc3D
D;RRRRkR#CHCCC38#0_oDFHkO_Mo#HM3C8N;DD
M
C0$H0R_1A7hww H1R#R
RRsbF0RR5
RRRRR R:MRHR0R#8F_DoRHO:'=R]
';RRRR1:RRRRHMR8#0_oDFH
O;STRRRRR:FRk0R8#0_oDFH
O;S7RRRRR:HRMR#_08DHFoOS;
RRRBRH:RM#RR0D8_FOoHR;R2
RSR
8CMR_1A7hww R1;
0N0skHL0#CR$LM_D	NO_GLFRRFV17A_w wh1RR:ObFlFMMC0#RHRk0sCR;

ONsECH0Os0kCkRVMFORVAR1_w7whR 1HL#
CMoH
sRbF#OC#R5B,2R1
RRRLHCoMR
SRRHV5CB'P0CMR8NMR=BRR''j2)RmR'51CMPC0MRN8RR1=4R''R2R0MEC
RSRRVRHR= RR''4RC0EM
RRSRRRRRRRH1VRR'=R4E'0CSM
SRRRRRRRRTRRRR<=';4'
RSSRRRRCCD#
RSSRRRRRRRRR<TR=;R7
RRRRRRRRMRC8VRH;R
RRRRRCRM8H
V;RRRRCRM8H
V;RCRRMb8RsCFO#
#;CRM8RMVkO
;

-
--R--Bp pR_1A)cqvihh)W-R--
--DsHLNRs$Q   ;#
kC RQ 1 3ap7_mBtQ_n44cD3NDk;
#QCR 3  1_a7pQmtBh_z1hQt N73D
D;kR#CQ   38#0_oDFHNO_sEH03DND;1
z  RQ M 3kslCH#O_0q83p
p;
0CMHR0$1)A_qivchW)hR
H#
oRRCsMCH5ORRR
RRRRRRRRRRQQhaR_j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QanRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ(a_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QaqRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQAa_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQwa_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jjRR
RRRRRRRRRRRR2;R
RRRRRRRRRb0Fs5RR
RRRRRRRRRRRRR)RR7qqaRF:Rk#0R0D8_FOoH_OPC05FsRR46RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRp)BiRhR:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRBR)pRi :MRHR0R#8F_DoRHO:'=R]
';RRRRRRRRRRRRRRRR)R RRRR:HRMR#_08DHFoO=R:R''];R
RRRRRRRRRRRRRRqR)7R7):MRHR0R#8F_Do_HOP0COFRs5(8RRF0IMF2RjRR;
RRRRRRRRRRRRRWRRBhpiRRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRRWiBp RR:HRMR#_08DHFoO=R:R''];R
RRRRRRRRRRRRRR RWRRRR:MRHR0R#8F_DoRHO:'=R]
';RRRRRRRRRRRRRRRRW7q7)RR:HRMR#_08DHFoOC_POs0F5RR(RI8FMR0Fj;2R
RRRRRRRRRRRRRRRR1vqi:RRRRHMR8#0_oDFHPO_CFO0s45R68RRF0IMF2RjRR;
RRRRRRRRRRRRRWRR7qqaRH:RM#RR0D8_FOoH_OPC05FsRR46RI8FMR0FjR2
RRRRRRRRRRRRR;R2

RRRCR
M18RAq_)vhci);hW
0N0skHL0#CR$LM_D	NO_GLFRRFV1)A_qivchW)hRO:RFFlbM0CMRRH#0Csk;



ONsECH0Os0kCAR1_v)qc)ihheW_RRFV1)A_qivchW)hR
H#RRRR
R
R#MHoNvDR :vRR8#0_oDFHPO_CFO0sj5cg86RF0IMF2RjR
;

#RRHNoMDqR)7_7)H:MRR0HMCsoCRMsNojCRRR0F.R66;R
R#MHoNWDRq)77_RHM:MRH0CCosNRsMRoCjFR0R6.6RR;
Ro#HMRNDqs88C_##BDFDHF#HMC_700COC:8RR8#0_oDFH;OR
C
LoRHM
R
RbOsFC5##)W , q,W7,7))7q7)R2
RRRRRoLCHRM
RRRRRRRRRRHV5WR5 RR='24'RMRN8)R5 RR='24'R8NMRW5Rq)77R)=Rq)772RR20MEC
RRRRRRRRRRRR8Rq8#sC#F_BD#DHH_FM7CC0O80CRR<=';4'
RRRRRRRRCRRD
#CRRRRRRRRRRRRR8q8s#C#_DBFDHH#F7M_CO0C0RC8<'=Rj;'R
RRRRRRRRCRRMH8RV
R;
RRRRRRRRNRR#s#C0qR58C8s#B#_FHDD#MHF_07CCCO08RR='2j'
RRRRRRRRRRRRbsCFRs0"8q8s#C#_DBFDHH#F
M"RRRRRRRRRRRR#CCPs$H0RsINMoHMR
;RRMRC8sRbF#OC#
;R
WRRsCH0ANCEPsHFRb:RsCFO#W#5Bhpi2R

RPRRNNsHLRDCv_ v0bClR#:R0D8_FOoH_OPC05Fsc6jgRI8FMR0Fj:2R=FRa_810pHFoOOeC05FsQahQ_Rw2&R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRa1F_0F8poeHOCFO0sh5QQ a_2
R&RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRFRa_810pHFoOOeC05FsQahQ_R72&R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRa1F_0F8poeHOCFO0sh5QQBa_2
R&RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRFRa_810pHFoOOeC05FsQahQ_RA2&R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRa1F_0F8poeHOCFO0sh5QQqa_2
R&RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRFRa_810pHFoOOeC05FsQahQ_Rg2&R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRa1F_0F8poeHOCFO0sh5QQUa_2
R&RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRFRa_810pHFoOOeC05FsQahQ_R(2&R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRa1F_0F8poeHOCFO0sh5QQna_2
R&RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRFRa_810pHFoOOeC05FsQahQ_R62&R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRa1F_0F8poeHOCFO0sh5QQca_2
R&RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRFRa_810pHFoOOeC05FsQahQ_Rd2&R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRa1F_0F8poeHOCFO0sh5QQ.a_2
R&RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRFRa_810pHFoOOeC05FsQahQ_R42&R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRa1F_0F8poeHOCFO0sh5QQja_2
;
RCRLo
HM
RRRR7Wq7H)_M=R<RMOFPM_H0CCosq5W727)RR;
RR
RRVRHRW5RBhpi'CCPMN0RM58RWiBphRR='2j'R8NMRB5WpRi =4R''N2RM58RW= RR''42RR20MEC
RRRRRRRVRFsHMRHR0jRF6R4RFDFbR
RRRRRRHRRVvR5q51iH=2RR''j2ER0CRM
RRRRRRRRRvRR 0v_C5lb4Wn*q)77_RHM+RRH2:RR=7RWq5aqH;2R
RRRRRRRRMRC8VRHRR;
RRRRRMRC8FRDF;bR
RRRR8CMRRHV;
R
RRRRvR v<v=R 0v_CRlb;


RMRC8sRbF#OC#
R;
R
R)8CNANCEPsHFRb:RsCFO#)#5Bhpi2R
R
RRRRsPNHDNLC7R)q_aq0bClR#:R0D8_FOoH_OPC05FsRR46RI8FMR0Fj;2RRR
RRRR
RoLCH
MR
RRRR7)q7H)_M=R<RMOFPM_H0CCosq5)727)R
;
RRRRH5VRR8q8s#C#_DBFDHH#F7M_CO0C0RC8=4R''02RE
CMRRRRRRRR)a7qqC_0l:bR=FR50sEC#>R=R''X2
R;RRRRCHD#VRR5)iBphP'CCRM0NRM85p)Bi=hRR''j2MRN8)R5B piR'=R4R'2NRM85R) =4R''22RRC0EMR
RRRRRRsVFRHHRMRRj04FR6FRDFRb
RRRRRRRRR)RR7qqa_l0CbR5H2=R:Rvv 5*4n)7q7)M_HRH+RRR2R;R
RRRRRR8CMRFDFb
R;RRRRCRM8H;VRRR

R)RR7qqaRR<=)a7qqC_0l;bR
R

R8CMRFbsO#C#R
;

8CMR_1A)cqvihh)W;_e



----- RBp1pRAq_)vhciW-R--
--DsHLNRs$Q   ;#
kC RQ 1 3ap7_mBtQ_n44cD3NDk;
#QCR 3  1_a7pQmtBh_z1hQt N73D
D;kR#CQ   38#0_oDFHNO_sEH03DND;1
z  RQ M 3kslCH#O_0q83p
p;
0CMHR0$1)A_qivchHWR#R

RMoCCOsHR
5RRRRRRRRRRQRRh_QajRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ4a_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QacRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ6a_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QaURR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQga_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QaBRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ7a_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_ :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
"RRRRRRRRRRRRR2
R;RRRRRRRRRFRbsR05
RRRRRRRRRRRRRRRRq)7a:qRR0FkR8#0_oDFHPO_CFO0s45R68RRF0IMF2RjRR;
RRRRRRRRRRRRR)RRBRpiRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRR)RRB piRH:RM#RR0D8_FOoHRR:=';]'
RRRRRRRRRRRRRRRRR) R:RRRRHMR8#0_oDFH:OR=]R''R;
RRRRRRRRRRRRR)RRq)77RH:RM#RR0D8_FOoH_OPC05FsRR(R8MFI0jFR2
R;RRRRRRRRRRRRRRRRWiBph:RRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRpWBi: RRRHMR8#0_oDFH:OR=]R''R;
RRRRRRRRRRRRRWRR RRRRH:RM#RR0D8_FOoHRR:=';]'
RRRRRRRRRRRRRRRR7Wq7:)RRRHMR8#0_oDFHPO_CFO0s(5RRFR8IFM0RRj2;R
RRRRRRRRRRRRRRqRv1RiR:MRHR0R#8F_Do_HOP0COFRs54R6R8MFI0jFR2
R;RRRRRRRRRRRRRRRRWa7qqRR:HRMR#_08DHFoOC_POs0F56R4RFR8IFM0R
j2RRRRRRRRRRRRR2RR;R
R

RRCRM81)A_qivch
W;Ns00H0LkC$R#MD_LN_O	LRFGF1VRAq_)vhciWRR:ObFlFMMC0#RHRk0sC
;

s
NO0EHCkO0s1CRAq_)vhciWR_eF1VRAq_)vhciW#RH
RRRRR

Ro#HMRNDvR v:0R#8F_Do_HOP0COFcs5jRg68MFI0jFR2
R;
R
R#MHoN)DRq)77_RHM:MRH0CCosNRsMRoCjFR0R6.6RR;
Ro#HMRNDW7q7)M_HRH:RMo0CCssRNCMoR0jRF6R.6
R;RHR#oDMNR8q8s#C#_DBFDHH#F7M_CO0C0RC8:0R#8F_DoRHO;L

CMoHRR

RFbsO#C#5,) WW ,q)77,7)q7
)2RRRRRCRLo
HMRRRRRRRRRVRHR55RW= RR''42NRRM58R)= RR''42MRN8RR5W7q7)RR=)7q7)22RRC0EMR
RRRRRRRRRRqRR8C8s#B#_FHDD#MHF_07CCCO08=R<R''4;R
RRRRRRRRRCCD#
RRRRRRRRRRRR8Rq8#sC#F_BD#DHH_FM7CC0O80CRR<='Rj';R
RRRRRRRRRCRM8H;VR
R
RRRRRRRRRNC##s50Rqs88C_##BDFDHF#HMC_700COC=8RR''j2R
RRRRRRRRRRCRsb0FsR8"q8#sC#F_BD#DHH"FM
RRRRRRRRRRRRP#CC0sH$NRIsMMHoRR;
CRRMb8RsCFO#R#;
R
RW0sHCEACNFPHsRR:bOsFC5##WiBph
2
RRRRPHNsNCLDRvv _l0CbRR:#_08DHFoOC_POs0F5gcj6FR8IFM0RRj2:a=RF0_18opFHCOeOs0F5QQha2_wRR&
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR_aF1p08FOoHe0COFQs5h_Qa &2R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRaRRF0_18opFHCOeOs0F5QQha2_7RR&
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR_aF1p08FOoHe0COFQs5h_QaB&2R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRaRRF0_18opFHCOeOs0F5QQha2_ARR&
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR_aF1p08FOoHe0COFQs5h_Qaq&2R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRaRRF0_18opFHCOeOs0F5QQha2_gRR&
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR_aF1p08FOoHe0COFQs5h_QaU&2R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRaRRF0_18opFHCOeOs0F5QQha2_(RR&
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR_aF1p08FOoHe0COFQs5h_Qan&2R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRaRRF0_18opFHCOeOs0F5QQha2_6RR&
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR_aF1p08FOoHe0COFQs5h_Qac&2R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRaRRF0_18opFHCOeOs0F5QQha2_dRR&
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR_aF1p08FOoHe0COFQs5h_Qa.&2R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRaRRF0_18opFHCOeOs0F5QQha2_4RR&
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR_aF1p08FOoHe0COFQs5h_Qaj
2;
LRRCMoH
R
RRqRW7_7)H<MR=FROMHP_Mo0CCWs5q)772
R;RRR
RHRRVRR5WiBphP'CCRM0NRM85pWBi=hRR''j2MRN8WR5B piR'=R4R'2NRM85RW =4R''22RRC0EMR
RRRRRRsVFRHHRMRRj04FR6FRDFRb
RRRRRRRRH5VRviq15RH2=jR''02RE
CMRRRRRRRRRRRRv_ v0bCl5*4nW7q7)M_HRH+RRR2R:W=R7qqa5RH2;R
RRRRRRCRRMH8RV
R;RRRRRCRRMD8RFRFb;R
RRMRC8VRHR
;R
RRRRvv RR<=v_ v0bClR
;

CRRMb8RsCFO#;#R
R

RN)C8EACNFPHsRR:bOsFC5##)iBp2R
R
RRRRsPNHDNLC7R)q_aq0bClR#:R0D8_FOoH_OPC05FsRR46RI8FMR0Fj;2RRR
RRRR
RoLCH
MR
RRRR7)q7H)_M=R<RMOFPM_H0CCosq5)727)RR;
RR
RRVRHRq5R8C8s#B#_FHDD#MHF_07CCCO08RR='24'RC0EMR
RRRRRR7R)q_aq0bClRR:=5EF0CRs#='>RXR'2;R
RRDRC#RHV5BR)pCi'P0CMR8NMRB5)p=iRR''42MRN8)R5B piR'=R4R'2NRM85R) =4R''22RRC0EMR
RRRRRRsVFRHHRMRRj04FR6FRDFRb
RRRRRRRRR)RR7qqa_l0CbR5H2=R:Rvv 5*4n)7q7)M_HRH+RRR2R;R
RRRRRR8CMRFDFb
R;RRRRCRM8H;VRRR

R)RR7qqaRR<=)a7qqC_0l;bR
R

R8CMRFbsO#C#R
;

8CMR_1A)cqvi_hWe
;

-
--R--Bp pR_1A)cqviRh)-----H
DLssN$ RQ 
 ;kR#CQ   371a_tpmQ4B_43ncN;DD
Ck#R Q  a317m_pt_QBzQh1t7h 3DND;#
kC RQ # 30D8_FOoH_HNs0NE3D
D;zR1 Q   3lMkCOsH_8#03pqp;C

M00H$AR1_v)qc)ihR
H#
oRRCsMCH5ORRR
RRRRRRRRRRQQhaR_j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQda_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QanRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ(a_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QaqRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQAa_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQwa_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jjRR
RRRRRRRRRRRR2;R
RRRRRRRRRb0Fs5RR
RRRRRRRRRRRRR)RR7qqaRF:Rk#0R0D8_FOoH_OPC05FsRR46RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRp)BiRhR:MRHR0R#8F_DoRHO;R
RRRRRRRRRRRRRRBR)pRi :MRHR0R#8F_DoRHO:'=R]
';RRRRRRRRRRRRRRRR)R RRRR:HRMR#_08DHFoO=R:R''];R
RRRRRRRRRRRRRRqR)7R7):MRHR0R#8F_Do_HOP0COFRs5(8RRF0IMF2RjRR;
RRRRRRRRRRRRRWRRBRpiRH:RM#RR0D8_FOoHRR;
RRRRRRRRRRRRRWRRB piRH:RM#RR0D8_FOoHRR:=';]'
RRRRRRRRRRRRRRRRRW R:RRRRHMR8#0_oDFH:OR=]R''R;
RRRRRRRRRRRRRWRRq)77RH:RM#RR0D8_FOoH_OPC05FsRR(R8MFI0jFR2
R;RRRRRRRRRRRRRRRRviq1RRR:HRMR#_08DHFoOC_POs0F56R4RFR8IFM0RRj2;R
RRRRRRRRRRRRRR7RWqRaq:MRHR0R#8F_Do_HOP0COFRs54R6R8MFI0jFR2R
RRRRRRRRRRRRRR
2;RRR
RM
C8AR1_v)qc)ih;0
N0LsHkR0C#_$MLODN	F_LGVRFR_1A)cqviRh):FROlMbFCRM0H0#Rs;kC



NEsOHO0C0CksR_1A)cqvi_h)eVRFR_1A)cqviRh)HR#
R
RR
#RRHNoMD RvvRR:#_08DHFoOC_POs0F5gcj6FR8IFM0RRj2;


RHR#oDMNR7)q7H)_MRR:HCM0oRCssoNMCRRj0.FR6;6R
#RRHNoMDqRW7_7)H:MRR0HMCsoCRMsNojCRRR0F.R66;R
R#MHoNqDR8C8s#B#_FHDD#MHF_07CCCO08RR:#_08DHFoO
R;RLR
CMoHRR

RFbsO#C#5,) WW ,q)77,7)q7
)2RRRRRCRLo
HMRRRRRRRRRVRHR55RW= RR''42NRRM58R)= RR''42MRN8RR5W7q7)RR=)7q7)22RRC0EMR
RRRRRRRRRRqRR8C8s#B#_FHDD#MHF_07CCCO08=R<R''4;R
RRRRRRRRRCCD#
RRRRRRRRRRRR8Rq8#sC#F_BD#DHH_FM7CC0O80CRR<='Rj';R
RRRRRRRRRCRM8H;VR
R
RRRRRRRRRNC##s50Rqs88C_##BDFDHF#HMC_700COC=8RR''j2R
RRRRRRRRRRCRsb0FsR8"q8#sC#F_BD#DHH"FM
RRRRRRRRRRRRP#CC0sH$NRIsMMHoRR;
CRRMb8RsCFO#R#;
R
RW0sHCEACNFPHsRR:bOsFC5##WiBp2R

RPRRNNsHLRDCv_ v0bClR#:R0D8_FOoH_OPC05Fsc6jgRI8FMR0Fj:2R=FRa_810pHFoOOeC05FsQahQ_Rw2&R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRa1F_0F8poeHOCFO0sh5QQ a_2
R&RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRFRa_810pHFoOOeC05FsQahQ_R72&R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRa1F_0F8poeHOCFO0sh5QQBa_2
R&RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRFRa_810pHFoOOeC05FsQahQ_RA2&R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRa1F_0F8poeHOCFO0sh5QQqa_2
R&RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRFRa_810pHFoOOeC05FsQahQ_Rg2&R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRa1F_0F8poeHOCFO0sh5QQUa_2
R&RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRFRa_810pHFoOOeC05FsQahQ_R(2&R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRa1F_0F8poeHOCFO0sh5QQna_2
R&RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRFRa_810pHFoOOeC05FsQahQ_R62&R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRa1F_0F8poeHOCFO0sh5QQca_2
R&RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRFRa_810pHFoOOeC05FsQahQ_Rd2&R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRa1F_0F8poeHOCFO0sh5QQ.a_2
R&RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRFRa_810pHFoOOeC05FsQahQ_R42&R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRa1F_0F8poeHOCFO0sh5QQja_2
;
RCRLo
HM
RRRR7Wq7H)_M=R<RMOFPM_H0CCosq5W727)RR;
RR
RRVRHRW5RB'piCMPC0MRN8WR5BRpi=4R''N2RM58RWiBp RR='24'R8NMR 5WR'=R4R'22ER0CRM
RRRRRFRVsRRHHjMRRR0F4D6RF
FbRRRRRRRRRRHV51vqi25HR'=RjR'20MEC
RRRRRRRRRRRRvv _l0Cbn54*7Wq7H)_MRR+HRR2RR:=Wa7qq25HRR;
RRRRRRRRCRM8H;VR
RRRRRRRCRM8DbFFRR;
RCRRMH8RVRR;
R
RR Rvv=R<Rvv _l0Cb
R;
R
RCRM8bOsFCR##;


RCR)NC8AEHNPF:sRRFbsO#C#5p)Bi
h2RRR
RPRRNNsHLRDC)a7qqC_0l:bRR8#0_oDFHPO_CFO0s45R68RRF0IMF2RjR
;RRRRR
LRRCMoHRR

R)RRq)77_RHM<O=RF_MPHCM0o5Cs)7q7);2R

RRRRRRH5VRR8q8s#C#_DBFDHH#F7M_CO0C0RC8=4R''02RE
CMRRRRRRRR)a7qqC_0l:bR=FR50sEC#>R=R''X2
R;RRRRCHD#VRR5)iBphP'CCRM0NRM85p)Bi=hRR''j2MRN8)R5B piR'=R4R'2NRM85R) =4R''22RRC0EMR
RRRRRRsVFRHHRMRRj04FR6FRDFRb
RRRRRRRRR)RR7qqa_l0CbR5H2=R:Rvv 5*4n)7q7)M_HRH+RRR2R;R
RRRRRR8CMRFDFb
R;RRRRCRM8H;VRRR

R)RR7qqaRR<=)a7qqC_0l;bR
R

R8CMRFbsO#C#R
;
CRM81)A_qivche)_;



----B-R Rpp1)A_qivcR----D-
HNLssQ$R ;  
Ck#R Q  a317m_pt_QB4c4n3DND;#
kC RQ 1 3ap7_mBtQ_1zhQ th7D3NDk;
#QCR 3  #_08DHFoOs_NH30EN;DD
 z1R Q  k3MlHCsO0_#8p3qp
;
CHM001$RAq_)vRciH
#
RCRoMHCsORR5
RRRRRRRRRRRQahQ_:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ.a_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQna_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_QagRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQqa_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RRRRRRRRRRRQahQ_:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";RRRRRRRRRQRRh_Qa7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R;
RRRRRRRRRhRQQ a_RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
RRRRRRRRRRQQhaR_w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjRj"
RRRRRRRRRRRR;2R
RRRRRRRRbRRF5s0RR
RRRRRRRRRRRRRR7R)qRaq:kRF00R#8F_Do_HOP0COFRs54R6R8MFI0jFR2
R;RRRRRRRRRRRRRRRR)iBpRRR:HRMR#_08DHFoO
R;RRRRRRRRRRRRRRRR)iBp RR:HRMR#_08DHFoO=R:R''];R
RRRRRRRRRRRRRR R)RRRR:MRHR0R#8F_DoRHO:'=R]
';RRRRRRRRRRRRRRRR)7q7)RR:HRMR#_08DHFoOC_POs0F5RR(RI8FMR0Fj;2R
RRRRRRRRRRRRRRRRpWBi:RRRRHMR8#0_oDFH;OR
RRRRRRRRRRRRRRRRpWBi: RRRHMR8#0_oDFH:OR=]R''R;
RRRRRRRRRRRRRWRR RRRRH:RM#RR0D8_FOoHRR:=';]'
RRRRRRRRRRRRRRRR7Wq7:)RRRHMR8#0_oDFHPO_CFO0s(5RRFR8IFM0RRj2;R
RRRRRRRRRRRRRRqRv1RiR:MRHR0R#8F_Do_HOP0COFRs54R6R8MFI0jFR2
R;RRRRRRRRRRRRRRRRWa7qqRR:HRMR#_08DHFoOC_POs0F56R4RFR8IFM0R
j2RRRRRRRRRRRRR2RR;R
R

RRCRM81)A_qivc;0
N0LsHkR0C#_$MLODN	F_LGVRFR_1A)cqviRR:ObFlFMMC0#RHRk0sC
;

s
NO0EHCkO0s1CRAq_)v_cieVRFR_1A)cqvi#RH
RRRRR

Ro#HMRNDvR v:0R#8F_Do_HOP0COFcs5jRg68MFI0jFR2
R;
R
R#MHoN)DRq)77_RHM:MRH0CCosNRsMRoCjFR0R6.6RR;
Ro#HMRNDW7q7)M_HRH:RMo0CCssRNCMoR0jRF6R.6
R;RHR#oDMNR8q8s#C#_DBFDHH#F7M_CO0C0RC8:0R#8F_DoRHO;L

CMoHRR

RFbsO#C#5,) WW ,q)77,7)q7
)2RRRRRCRLo
HMRRRRRRRRRVRHR55RW= RR''42NRRM58R)= RR''42MRN8RR5W7q7)RR=)7q7)22RRC0EMR
RRRRRRRRRRqRR8C8s#B#_FHDD#MHF_07CCCO08=R<R''4;R
RRRRRRRRRCCD#
RRRRRRRRRRRR8Rq8#sC#F_BD#DHH_FM7CC0O80CRR<='Rj';R
RRRRRRRRRCRM8H;VR
R
RRRRRRRRRNC##s50Rqs88C_##BDFDHF#HMC_700COC=8RR''j2R
RRRRRRRRRRCRsb0FsR8"q8#sC#F_BD#DHH"FM
RRRRRRRRRRRRP#CC0sH$NRIsMMHoRR;
CRRMb8RsCFO#R#;
R
RW0sHCEACNFPHsRR:bOsFC5##WiBp2R

RPRRNNsHLRDCv_ v0bClR#:R0D8_FOoH_OPC05Fsc6jgRI8FMR0Fj:2R=FRa_810pHFoOOeC05FsQahQ_Rw2&R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRa1F_0F8poeHOCFO0sh5QQ a_2
R&RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRFRa_810pHFoOOeC05FsQahQ_R72&R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRa1F_0F8poeHOCFO0sh5QQBa_2
R&RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRFRa_810pHFoOOeC05FsQahQ_RA2&R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRa1F_0F8poeHOCFO0sh5QQqa_2
R&RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRFRa_810pHFoOOeC05FsQahQ_Rg2&R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRa1F_0F8poeHOCFO0sh5QQUa_2
R&RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRFRa_810pHFoOOeC05FsQahQ_R(2&R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRa1F_0F8poeHOCFO0sh5QQna_2
R&RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRFRa_810pHFoOOeC05FsQahQ_R62&R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRa1F_0F8poeHOCFO0sh5QQca_2
R&RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRFRa_810pHFoOOeC05FsQahQ_Rd2&R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRa1F_0F8poeHOCFO0sh5QQ.a_2
R&RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRFRa_810pHFoOOeC05FsQahQ_R42&R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRa1F_0F8poeHOCFO0sh5QQja_2
;
RCRLo
HM
RRRR7Wq7H)_M=R<RMOFPM_H0CCosq5W727)R
;
RRRRH5VRRpWBiP'CCRM0NRM85pWBiRR='24'R8NMRB5WpRi =4R''N2RM58RW= RR''42RR20MEC
RRRRRRRVRFsHMRHR0jRF6R4RFDFbR
RRRRRRHRRVvR5q51iH=2RR''j2ER0CRM
RRRRRRRRRvRR 0v_C5lb4Wn*q)77_RHM+RRH2:RR=7RWq5aqH;2R
RRRRRRRRMRC8VRHRR;
RRRRRMRC8FRDF;bR
RRRR8CMRRHV;
R
RRRRvR v<v=R 0v_CRlb;


RMRC8sRbF#OC#
R;
R
R)8CNANCEPsHFRb:RsCFO#)#5B2pi

RRRRRRPHNsNCLDRq)7a0q_CRlb:0R#8F_Do_HOP0COFRs54R6R8MFI0jFR2RR;
RRRRR
RLHCoM
R
RRRR)7q7)M_HRR<=OPFM_0HMCsoC57)q7R)2;R
R
RRRRRHV58Rq8#sC#F_BD#DHH_FM7CC0O80CR'=R4R'20MEC
RRRRRRRRq)7a0q_CRlb:5=RFC0Es=#R>XR'';2R
RRRR#CDH5VRRp)BiP'CCRM0NRM85p)BiRR='24'R8NMRB5)pRi =4R''N2RM58R)= RR''42RR20MEC
RRRRRRRVRFsHMRHR0jRF6R4RFDFbR
RRRRRRRRRR7R)q_aq0bCl52HRRR:=v5 v4)n*q)77_RHM+RRH2;RR
RRRRRRRCRM8DbFFRR;
RCRRMH8RVRR;
R
RR7R)qRaq<)=R7qqa_l0Cb
R;
R
RCRM8bOsFCR##;


CRM81)A_qivc_
e;
-----------------------------------------------------------------------------
-SSSSSCbs_
HF----------------------------------------------------------------------------
LDHs$NsRCHCCk;
#HCRC3CC#_08DHFoO4_4nNc3D
D;kR#CHCCC38#0_oDFHNO_sEH03DND;#
kCCRHC#C30D8_FOoH_#kMHCoM8D3ND
;
CHM00b$SsHC_F#SH
b
SFSs05S
SS_L#CSMS:MSHS8#0_oDFHSO;SK--aRqtCLMNDRCRRRRRRRRRRS
SSH#EVS0S:MSHS8#0_oDFHSO;SK--aRqt#VEH0RRRRRRRRRRRRS
SSD0O	:SSSSHM#_08DHFoOS;S-a-KqOtRD	FORRRRRRRRRRRR
SSSkNb80SCS:MSHS8#0_oDFHSO;SK--aRqtkNb80RCRRRRRRRRRRS
SSH#8S:SSSSHM#_08DHFoOS;S-a-Kq#tRCNsHDNR80HNRMRRR
SSSlCF8SSS:H#MS0D8_FOoH;-SS-qKatFRl8RCRRRRRRRRRR
RRSESSHLx_SSS:H#MS0D8_FOoH;-SS-qKatHREoXERRMOF0DsFR
RRS#SS8SFSSF:Sk#0S0D8_FOoH;-SS-qKatCR#sDHNR08NNkRF0
RRS8SSF4k0SSS:FSk0#_08DHFoOS;S-F-hsDlNRbQMkO0RCRDDFbk0k40R
SSS80Fkj:SSS0FkS8#0_oDFHSO;Sh--FNslDMRQbRk0ODCDR0FkbRk0jS
SSs884:SSSSHM#_08DHFoOS;S-F-hsDlNR0mkbRk0ODCDRbHMk40R
SSS8j8sSSS:H#MS0D8_FOoH;-SS-shFlRNDmbk0kO0RCRDDHkMb0
RjSFSSCMbHSSS:H#MS0D8_FOoH;-SS-shFlRNDmkkb0M- NCLDRRRRR
RRSESSFSD8SH:SM0S#8F_Do;HOS-S-hlFsNQDRM0bkRDOCDFROMF0sDSR
S#Ss0SHFSH:SM0S#8F_Do;HOS-S-hlFsNQDRM0bkRDOCDCRs#RC0RSR
SMSHOSD	SH:SM0S#8F_Do;HOS-S-hlFsNQDRM0bkRDOCDDROFRO	RSR
SkSF0	ODSSS:H#MS0D8_FOoH;-SS-shFlRNDmbk0kO0RCRDDOODF	
RRSOSSLSH0SH:SM0S#8F_Do_HOP0COF5sR6FR8IFM0R;j2SB--FHMVoHksFLMRHR0#RSR
SNSb8SHMSH:SM0S#8F_Do;HOS-S-uRq7HkMb0RRRRRRRR
RRSbSSNk8F0:SSS0FkS8#0_oDFHSO;Su--qF7Rkk0b0RRRRRRRRSR
SNSb8MFCSSS:FSk0#_08DHFoOSRS-q-u7kRF00bkRNCMLRDCRS
SS
2;
8CMRCbs_;HF
s
NO0EHCkO0sbCRsHC_FR_PFbVRsHC_F#RH
HS#oDMNS8bNHMM_4M,HO_D	Mb.,NM8H_SMd:0S#8F_Do;HO
HS#oDMNS_HMv_zXM:cSS8#0_oDFH
O;So#HMSNDE8FD_7qh.SS:#_08DHFoOS;
#MHoN8DS8_sjMS44:0S#8F_Do;HO
HS#oDMNS0FkO_D	MS4.:0S#8F_Do;HO
HS#oDMNSs8844_MdSS:#_08DHFoOS;
#MHoNMDS4ScSS#:S0D8_FOoH;#
SHNoMDFS8ks0_Cjo__:MSS8#0_oDFH
O;So#HMSND)_CoFWs_H_sChS4(:0S#8F_Do;HO
HS#oDMNSUM4S:SSS8#0_oDFH
O;So#HMSNDMS4gSSS:#_08DHFoOS;
#MHoN0DSs0H#NS0C:0S#8F_Do;HO
HS#oDMNS0FkO_D	MS..:0S#8F_Do;HO
HS#oDMNSnM.S:SSS8#0_oDFH
O;So#HMSNDF_CMM._McSS:#_08DHFoOS;
#MHoN[DS0_NokNb80MC_d:jSS8#0_oDFH
O;So#HMSND8_HMs_CojSS:#_08DHFoOS;
#MHoNRDR8_HMs_Co4SS:#_08DHFoOS;
#MHoN8DSF_k0s_CojSS:#_08DHFoOS;
#MHoN8DSF_k0s_Co4SS:#_08DHFoOS;
#MHoN0DSs0H#N_0CJSS:#_08DHFoOS;
#MHoN[DS0_NoFsC_C:oSS8#0_oDFH
O;So#HMSND0bCl4C,0lSb.S#:S0D8_FOoH_OPC0RFs584RF0IMF2Rj;#
SHNoMDFS8kj0_SSS:#_08DHFoOS;S-I-SHRsCVRFsb0FsRo#HMRNDko#NCC
Lo
HMSN[0ob_k8CN0_jMdSS<=MSF05_L#CNMRM58RMRF0kNb802C2;

SSF#8S=S<SM8H_osC_
j;Sk8F0S4R<S=R8_HMs_Co4-;
-------------------------------------------------------------SS
bHN8M4_M_:HSSFbsO#C#SF58ks0_Cjo_,NRb8,HMRH#EV
02SSSSLHCoMS
SSHSSV#S5E0HV=''42ES0CSM
SSSSS8bNHMM_4=S<Sk8F0C_so;_j
SSSSDSC#SC
SSSSS8bNHMM_4=S<S8bNH
M;SSSSS8CMR;HV
SSSS8CMSFbsO#C#;

SSOHMDM	_.S_H:sSbF#OC#LS5#M_C,OR0DR	,HDMO	S2
SLSSCMoH
SSSSVSHS#5L_=CM'24'SC0EMS
SSSSSHDMO	._MSS<=0	OD;S
SSCSSD
#CSSSSSMSHO_D	M<.S=MSHO;D	
SSSSMSC8VRH;S
SSMSC8sRbF#OC#
;
SM8H_osC_Hj_Sb:SsCFO#5#SHDMO	._M,#Rs02HF
SSSSoLCHSM
SSSSH5VSsH#0F4=''02SE
CMSSSSSHS8MC_soS_j<'=Sj
';SSSSS#CDH5VSHDMO	._MRP'CCRM0NRM8HDMO	._M=''42ER0CSM
SSSSSM8H_osC_<jS=NSb8_HMM
4;SSSSS8CMR;HV
SSSS8CMRFbsO#C#;-
----------------------------------------------------------S--S
SSS8bNHMM_dS_H:sSbF#OC#LS5#M_C,HR8MC_so,_jR8bNH
M2SSSSLHCoMS
SSHSSVLS5#M_C=''42ES0CSM
SSSSS8bNHMM_d=S<SM8H_osC_
j;SSSSS#CDCS
SSSSSbHN8Md_MSS<=bHN8MS;
SSSSCRM8H
V;SSSSCSM8bOsFC;##
SS
8_HMs_Co4S_H:sSbF#OC#HS5M	OD_,M.R0s#H
F2SSSSLHCoMS
SSHSSVsS5#F0H=''42ES0CSM
SSSSSM8H_osC_<4S=jS''S;
SSSSCHD#VHS5M	OD_RM.'CCPMN0RMH8RM	OD_=M.'2j'RC0EMS
SSSSSH5VS[o0N_8kbN_0CM=dj'24'SC0EMS
SSSSSSM8H_osC_<4S=NSb8_HMM
d;SSSSSMSC8VRH;S
SSCSSMH8RVS;
SCSSMb8RsCFO#
#;-------------------------------------------------------------
-SSDEF8h_q7<.R=LROH4052MRN8FRED
8;
RRRSQ--M0bkRXvzRSRR
CS0lSb4<E=SF_D8q.h7RO&RL5H0j
2;
MSH_Xvz__McHSS:bOsFCS##5l0CbR4,80Fk_Rj,8_HMs_Cojb,RNM8H2R
RRSSSSoLCHRM
RSRSSOSSNS#C0bCl4#RH
RRRSSSSSCIEMjS"j="S>R
RRSSSSHSSMz_vXc_MRR<=8_HMs_CojR;
RSRSSISSESCM""j4S
=>RSRRSSSSS_HMv_zXM<cR=NRb8;HM
RRRSSSSSCIEM4S"j="S>R
RRSSSSHSSMz_vXc_MRR<=80Fk_
j;RSRRSSSSIMECS4"4">S=
RRRSSSSSMSH_Xvz_RMc<8=RF_k0jR;
RSRSSISSERCMFC0EsS#R=R>
RSRSSSSSHvM_zMX_c=R<R''j;R
RRSSSSMSC8NRO#
C;RSRRSCSSMb8RsCFO#
#;
------------------------k8F0ojRCsMCN-0C-----------------------------8
SF_k0jS_H:sSbF#OC#lS5F,8CRM8H_osC_R4,HvM_zMX_cS2
SCSLo
HMSSSSH5VSlCF8=''42ES0CSM
SSSS80Fk_<jS=HS8MC_so;_4
SSSS#CDCS
SS8SSF_k0j=S<S_HMv_zXM
c;SSSSCRM8H
V;SCSSMb8RsCFO#
#;S8
SFjk0SS<=80Fk_
j;--------------------------------------------------------------------S-
S-0mkbRk0)HCo#s0C
SS
80Fk_osC_Hj_Sb:SsCFO#5#SFOk0DM	_4R.,sH#0FS2
SLSSCMoH
SSSSVSHS#5s0=HF'24'SC0EMS
SSSSS80Fk_osC_<jS=jS''S;
SSSSCHD#VFS5kD0O	4_M.CR'P0CMR8NMR0FkO_D	M=4.'24'RC0EMS
SSSSS80Fk_osC_<jS=8S8sMj_4
4;SSSSS8CMR;HV
SSSS8CMRFbsO#C#;S

-k-vGRC#VRFsmbk0ks0RC#oH0#Cs
SS
80Fk_osC_Mj_R=S<R0MFRk8F0C_so;_j
4SMgSRSSR<=MRF050FkO_D	MR4.FOsRL5H0.;22
SS
)_CoFWs_H_sCh_4(HSS:bOsFCS##5HOL025.,FR8ks0_Cjo__RM,8j8s2S
SSLSSCMoH
SSSSHSSVOS5L5H0.'2=4S'20MEC
SSSSSSS)_CoFWs_H_sChS4(<8=SF_k0s_Coj;_M
SSSSCSSD
#CSSSSS)SSCFo_sH_WshC_4<(S=8S8s
j;SSSSSMSC8VRH;S
SSCSSMb8RsCFO#
#;SM
S4HU_SSSS:sSbF#OC#MS54Rg,80Fk_osC_R4,80Fk_osC_
j2SSSSSoLCHSM
SSSSSSHV5gM4=''42ES0CSM
SSSSS4SMU=S<Sk8F0C_so;_4
SSSSCSSD
#CSSSSSMSS4<US=FS8ks0_Cjo_;S
SSSSSCRM8H
V;SSSSS8CMRFbsO#C#;S

M_4cHSSSSb:SsCFO#5#SO0LH5,d2Ro)C__FsWCHs_(h4,4RMU
2SSSSSSoLCHSM
SSSSSSHV5HOL025d=''42ES0CSM
SSSSS4SMc=S<So)C__FsWCHs_(h4;S
SSSSSCCD#
SSSSSSSMS4c<M=S4
U;SSSSSMSC8VRH;S
SSCSSMb8RsCFO#
#;SSSSSb
SNk8F0S_HSSS:bOsFCS##58lFC8,RF_k0s_Co4M,R4
c2SSSSSoLCHSM
SSSSSSHV58lFC4=''02SE
CMSSSSSbSSNk8F0=S<Sk8F0C_so;_4
SSSSCSSD
#CSSSSSbSSNk8F0=S<ScM4;S
SSSSSCRM8H
V;SSSSS8CMRFbsO#C#;S

-a-KqqtR#o#HMS#

8S8sMj_4H4_SSS:bOsFCS##5H#EVR0,0#sH0CN0_RJ,8j8s2S
SSLSSCMoH
SSSSHSSV#S5E0HV=''42ES0CSM
SSSSS8S8sMj_4<4S=sS0HN#00JC_;S
SSSSSCCD#
SSSSSSS8j8s_4M4SS<=8j8s;S
SSSSSCRM8H
V;SSSSS8CMRFbsO#C#;S

FOk0DM	_4H._SSS:bOsFCS##5_L#CRM,0	OD,kRF0	OD2S
SSLSSCMoH
SSSSHSSVLS5#M_C=''42ES0CSM
SSSSSkSF0	OD_.M4SS<=0	OD;S
SSSSSCCD#
SSSSSSSFOk0DM	_4<.S=kSF0	OD;S
SSSSSCRM8H
V;SSSSS8CMRFbsO#C#;S
SS
SSSs8844_MdS_HSb:SsCFO#5#SLC#_M8,RF_k0s_Coj8,R82s4
SSSSCSLo
HMSSSSSVSHS#5L_=CM'24'SC0EMS
SSSSSSs8844_Md=S<Sk8F0C_so;_j
SSSSCSSD
#CSSSSS8SS8_s4MS4d<8=S8;s4
SSSSCSSMH8RVS;
SSSSCRM8bOsFC;##
-
S-qKatCRso0H#C
sRSk8F0C_so__4H:SSSFbsO#C#Sk5F0	OD_.M4,#Rs02HF
SSSSCSLo
HMSSSSSVSHS#5s0=HF'24'SC0EMS
SSSSSSk8F0C_soS_4<'=Sj
';SSSSSDSC#SHV50FkO_D	MR4.'CCPMN0RMF8RkD0O	4_M.j=''02RE
CMSSSSS8SSF_k0s_Co4=S<Ss8844_MdS;
SSSSS8CMR;HV
SSSSMSC8sRbF#OC#S;
SSSS
-----------------------------------------------------------------------------
-
S--mbk0k 0RMDNLCFRpo
HO---
----------------------------------------------------------------------------
-S-ma Rs0H#NR0C)HCo#s0C
sS0HN#00HC_Sb:SsCFO#5#S#VEH0#,R8RH,FHCbMS2
SLSSCMoH
SSSSVSHSE5#H=V0'24'SC0EMS
SSSSS0#sH0CN0SS<=#;8H
SSSSDSC#SC
SSSSSH0s#00NC=S<SbFCH
M;SSSSS8CMR;HV
SSSS8CMRFbsO#C#;S

0#sH0CN0_HJ_Sb:SsCFO#5#SFOk0DM	_.R.,sH#0FS2
SLSSCMoH
SSSSVSHS#5s0=HF'24'SC0EMS
SSSSS0#sH0CN0_<JS=jS''S;
SSSSCHD#VFS5kD0O	._M.CR'P0CMR8NMR0FkO_D	MR..=4R''02RE
CMSSSSSsS0HN#00JC_SS<=0#sH0CN0;S
SSCSSMH8RVS;
SCSSMb8RsCFO#
#;SSSS
-S-KtaqRosCHC#0sF
SkD0O	._M.S_H:sSbF#OC#LS5#M_C,OR0DR	,FOk0D
	2SSSSLHCoMS
SSHSSVLS5#M_C=''42ES0CSM
SSSSS0FkO_D	MS..<0=SO;D	
SSSSDSC#SC
SSSSS0FkO_D	MS..<F=SkD0O	S;
SSSSCRM8H
V;SSSSCRM8bOsFC;##
SS
[o0N__FCs_CoHSS:bOsFCS##50FkO_D	M,..R0s#H
F2SSSSLHCoMS
SSHSSVsS5#F0H=''42ES0CSM
SSSSSN[0oC_F_osCSS<=';j'
SSSSDSC#SHV50FkO_D	MR..'CCPMN0RMF8RkD0O	._M.'R=jR'20MEC
SSSSHSSV[S50_NokNb80MC_d'j=4S'20MEC
SSSSSSS[o0N__FCsSCo<b=SNM8H_;Md
SSSSCSSMH8RVS;
SSSSCRM8H
V;SSSSCRM8bOsFC;##
RS
R0RSC.lbSS<=O0LH5R62&LROHc052
;RR-RS-CSFM__MM_.cHSS:bOsFCS##5HOL0256,HOL025c,CRFb,HMRH0s#00NC2_JRR
RSMFC_MM_.Hc_Sb:SsCFO#5#S0bCl.F,RCMbH,sR0HN#00JC_2RR
RSSSSCSLoRHM
SRRSSSSSO--NS#CO0LH5R62&LROHc052#RHRR
RSSSSSNSO#0CSC.lbRRH#
SRRSSSSSESIC"MSjSj"=
>RRSRSSSSSSMFC_MM_.<cS=jS''
;RRSRSSSSSSCIEMjS"4="S>RR
RSSSSSSSF_CMM._Mc=S<S''4;RR
RSSSSSSSIMECSj"4">S=RR
RSSSSSFSSCMM__cM.SS<=FHCbM
;RRSRSSSSSSCIEM4S"4="S>R
RRSSSSSSSF_CMM._Mc=S<SH0s#00NC;_JRR
RRSSSSSSSIMECREF0CSs#SR=>
RRRSSSSSFSSCMM__cM.SS<=';j'RR
RRSSSSCSSMO8RN;#CRR
RRSSSSMSC8sRbF#OC#S;

.SMnS_HSSS:bOsFCS##58lFC[,R0_NoFsC_CRo,F_CMM._McS2
SLSSCMoH
SSSSVSHSF5l8'C=4S'20MEC
SSSSMSS.<nS=0S[NFo_CC_soS;
SSSSCCD#
SSSSMSS.<nS=CSFM__MM;.c
SSSSMSC8VRH;S
SSMSC8sRbF#OC#
;
S8bNFRCM<M=RF50RE_HxLMRN8.RMn
2;SM
C8sRbCF_H_
P;
-------------------------------------------------------------------------
-SSSSS_1AQ-m
---------------------------------------------------------------------
--
LDHs$NsRCHCCk;
#HCRC3CC#_08DHFoO4_4nNc3D
D;kR#CHCCC38#0_oDFHNO_sEH03DND;#
kCCRHC#C30D8_FOoH_#kMHCoM8D3ND-;
-LDHs$NsSsIF	k;
#ICSF3s	#_08DHFoOA_1aD3ND
;
CHM001$SAm_QR
H#
CSoMHCsO
R5ShSS at_)tQt :)RR0LHSSSSS=S:S''j;S
SShuQ_uaY RS:L_H0P0COF5sR6FR8IFM0RSj2:"=Sjjjjj;j"
SSSupzpzSuS:HRL0SSSS:SS=jS''S;
SmSQ_q1ah)7q7RS:#H0sMSoSS:SS=1S"Ae_pB1vm"S
SS
2;SsbF0SR
SS5
Sm7_z4a_RRSSR:RRRRHM#_08DHFoOS;
Sm7_zja_RRSSR:RRRRHM#_08DHFoOS;
SmBpB i_hpqA :SSRRHM#_08DHFoOS;
SapqBQ]_hauz_peqz: SRRHM#_08DHFoOS;
SuQhzBa_pSiSSH:RM0R#8F_Do;HO

SSS_S7Q4h_SSSS:kRF00R#8F_Do;HO
7SS__QhjSSSSF:Rk#0R0D8_FOoH;S
Smuzaz a_hpqA :SSRRHM#_08DHFoO=S:';]'
mSSzzauap_BiSSS:MRHR8#0_oDFH
O;SqSuBtiq Q_uhSSS:MRHFSk0#_08koDFHSO
SR2;

SSCRM81QA_m
R;Ns00H0LkC$R#MD_LN_O	LRFGF1VRAm_QRO:RFFlbM0CMRRH#0Csk;N

sHOE00COkRsC1QA_mR_eF1VRAm_QR
H#
FSOlMbFCSM0b_sCHSF
b0FsSS5
SFSED:8SSRHMS8#0_oDFH
O;SsSS#F0HSH:SM0S#8F_Do;HO
SSSLC#_MSS:H#MS0D8_FOoH;S
SSH#EV:0SSSHM#_08DHFoOS;
SOS0D:	SSSHM#_08DHFoOS;
SMSHOSD	:MSHS8#0_oDFH
O;SFSSkD0O	SS:H#MS0D8_FOoH;S
SS8kbNS0C:MSHS8#0_oDFH
O;SFSSCMbHSH:SM0S#8F_Do;HO
SSS#S8HSH:SM0S#8F_Do;HO
SSSlCF8SH:SM0S#8F_Do;HO
SSSE_HxLSS:H#MS0D8_FOoH;S
SSF#8SSS:FSk0#_08DHFoOS;
SFS8kS04:kSF00S#8F_Do;HO
SSS80FkjSS:FSk0#_08DHFoOS;
S8S8s:4SSSHM#_08DHFoOS;
S8S8s:jSSSHM#_08DHFoOS;
SNSb8SHM:MSHS8#0_oDFH
O;SbSSNk8F0SS:FSk0#_08DHFoOS;
SNSb8MFCSF:Sk#0S0D8_FOoH;S
SSHOL0SS:H#MS0D8_FOoH_OPC0SFs586RF0IMF2Rj
SSS2S;
CRM8ObFlFMMC0
;
So#HMSNDHDMO	,_MR0FkO_D	MH,RM	OD,kRF0	OD,F#8S#:S0D8_FOoH;

SSo#HMSNDLC#_MSS:#_08DHFoO=S:';j'SA--F8kMNRs$#MONRNCMLRDCRRRRRRRRRSR
#MHoN#DSE0HVS#:S0D8_FOoHS':=jS';-F-AkNM8s#$RORNM#VEH0RRRRRRRRRRRR#
SHNoMDOS0D:	SS8#0_oDFH:OS=''j;-S-AMFk8$NsRN#OMDROFRO	RRRRRRRRR
RRSo#HMSNDkNb80:CSS8#0_oDFH:OS=''j;-S-AMFk8$NsRN#OMbRk8CN0RRRRRRRRR
RRSo#HMSND#S8HS#:S0D8_FOoHS':=jS';-F-AkNM8s#$RORNM#HCsN8DRNR0NHRMRR#
SHNoMDFSl8:CSS8#0_oDFH:OS=''j;-S-AMFk8$NsRN#OMFRl8RCRRRRRRRRRR
RRSo#HMSNDE_HxLSS:#_08DHFoO=S:';4'SA--F8kMNRs$#MONRHas#00NCFROMF0sDSR

HS#oDMNSMbH_HOL0#:S0D8_FOoH_OPC05Fs6FR8IFM0R;j2
HS#oDMNSoMC_H0so#:S0D8_FOoH;#
SHNoMDkSbDkD_bSS:#_08DHFoOS;
#MHoNEDSF,D8FHCbMN,b8MFC,8bNF,k0bHN8MSS:#_08DHFoOL;
CMoH
SS
b_HMO0LHSS<=a1m_am7pteQB mBa)uS5Qah_Y2u ;M
SC0o_sSHo<a=Sma_17tpmQ5BSh_ tat)Qt2 );b
Sk_DDkSbS<a=Sma_17tpmQ5BSupzpz;u2
H
SM	OD_<MS=QRShauz_iBpRsGFRoMC_H0soS;
FOk0DM	_<m=Szzauap_BiFRGsCRMos_0H
o;SOHMD<	S=MSHO_D	MMRN8pRBm_Bi Ahqp
 ;S0FkOSD	<F=SkD0O	R_MNRM8BBpmih_ q Ap;

SSDEF8=S<SapqBQ]_hauz_peqz
 ;SbFCH<MS=zSmaauz_q hA;p 
SS
uiqBq_t u_QhHSS:bOsFCS##58bNF,CMR8bNF,k0RBuqi qt_huQ2L
SCMoH
bSSNM8HSS<=uiqBq_t u;Qh
HSSVbS5NC8FM4=''02RE
CMSuSSqqBitu _Q<hS=ZS''S;
S#CDCS
SSBuqi qt_huQSS<=bFN8k
0;SMSC8VRH;C
SMb8RsCFO#
#;-----------------------------------------------------------------SS
b_sCHHF_Sb:SsHC_Fb
SFRs0lSNb5S
SSFSED=8S>FSED
8,SSSSsH#0F>S=S''j,S
SS#SL_SCM=L>S#M_C,S
SSES#HSV0=#>SE0HV,S
SSOS0D=	S>OS0D
	,SSSSHDMO	>S=SOHMD
	,SSSSFOk0D=	S>kSF0	OD,S
SSbSk8CN0SS=>kNb80
C,SSSSFHCbM>S=SbFCH
M,SSSS#S8HSS=>#,8H
SSSS8lFC>S=S8lFCS,
SESSHLx_SS=>E_HxLS,
S#SS8SFS=#>S8
F,SSSS80Fk4>S=SQ7_h,_4
SSSSk8F0=jS>_S7Qjh_,S
SS8S8s=4S>_S7m_za4S,
S8SS8Ssj=7>S_amz_
j,SSSSbHN8M>S=S8bNH
M,SSSSbFN8k=0S>NSb80Fk,S
SSNSb8MFCSS=>bFN8C
M,SSSSO0LHSS=>b_HMO0LH
SSSS
2;CSM81QA_m;_e
-
---------------------------------------------------------------------
S--SSSS1tA_Am_Q
--------------------------------------------------------------------
--
LDHs$NsRCHCCk;
#HCRC3CC#_08DHFoO4_4nNc3D
D;kR#CHCCC38#0_oDFHNO_sEH03DND;#
kCCRHC#C30D8_FOoH_#kMHCoM8D3ND-;
-LDHs$NsSsIF	k;
#ICSF3s	#_08DHFoOA_1aD3ND
;
CHM001$SAA_t_RQmHS#
oCCMsSHO5S
SSth _Qa)t)t RL:RHS0SSSSS:'=Sj
';SuSSQah_YSu :HRL0C_POs0FRR568MFI0jFR2=S:Sj"jjjjj"S;
SzSupupzSRS:LSH0SSSSSS:=';j'
SSSQ1m_a7qhqS)7:0R#soHMSSSSSS:="_1ApveBm
1"S2SS;S
SSb
SFSs05S
SSBuqi qt_huQS:SSSFHMk#0S0k8_DHFoOS;
SqSpa_B]Qzhuaq_epSz :MSHS0S#8F_Do;HO
SSSBBpmih_ q ApRRRRRRRR:MSHS0S#8F_Do;HO
SSSQzhuap_BiRRRRRRRRRRR:MSHS0S#8F_Do;HO
SSSmuzazBa_pRiRRRRRRRRR:MSHS0S#8F_Do;HO
SSSmuzaz a_hpqA :SSRRHM#_08DHFoO=S:';]'
SSS7z_maR_4RRRRRRRRRRRR:MSHS0S#8F_Do;HO
SSS7z_maR_jRRRRRRRRRRRR:MSHS0S#8F_Do;HO
SSS7h_Q_R4RRRRRRRRRRRRR:kSF0#SS0D8_FOoH;S
SSQ7_hR_jRRRRRRRRRRRRRF:SkS0S#_08DHFoOS;
SpStmpAq_wAzw_ )muzazSa:FSk0S8#0_oDFHSO
S;S2
8CMR_1AtQA_mN;
0H0sLCk0RM#$_NLDOL	_FFGRVAR1__tAQ:mRRlOFbCFMMH0R#sR0k
C;
ONsECH0Os0kCAR1__tAQem_RRFV1tA_Am_QR
H#
FSOlMbFCSM0b_sCHSF
b0FsSS5
SFSED:8SSRHMS8#0_oDFH
O;SsSS#F0HSH:SM0S#8F_Do;HO
SSSLC#_MSS:H#MS0D8_FOoH;S
SSH#EV:0SSSHM#_08DHFoOS;
SOS0D:	SSSHM#_08DHFoOS;
SMSHOSD	:MSHS8#0_oDFH
O;SFSSkD0O	SS:H#MS0D8_FOoH;S
SS8kbNS0C:MSHS8#0_oDFH
O;SFSSCMbHSH:SM0S#8F_Do;HO
SSS#S8HSH:SM0S#8F_Do;HO
SSSlCF8SH:SM0S#8F_Do;HO
SSSE_HxLSS:H#MS0D8_FOoH;S
SSF#8SSS:FSk0#_08DHFoOS;
SFS8kS04:kSF00S#8F_Do;HO
SSS80FkjSS:FSk0#_08DHFoOS;
S8S8s:4SSSHM#_08DHFoOS;
S8S8s:jSSSHM#_08DHFoOS;
SNSb8SHM:MSHS8#0_oDFH
O;SbSSNk8F0SS:FSk0#_08DHFoOS;
SNSb8MFCSF:Sk#0S0D8_FOoH;S
SSHOL0SS:H#MS0D8_FOoH_OPC0SFs586RF0IMF2Rj
SSS2S;
CRM8ObFlFMMC0S;

HS#oDMNSOHMDM	_,0FkO_D	MM,HO,D	FOk0D#	,8:FSS8#0_oDFH
O;S#
SHNoMD#SL_SCM:0S#8F_DoSHO:j=''-;S-kAFMs8N$OR#NCMRMDNLCRRRRRRRRRRR
HS#oDMNSH#EV:0SS8#0_oDFH:OS=''j;-S-AMFk8$NsRN#OMER#HRV0RRRRRRRRR
RRSo#HMSND0	ODS#:S0D8_FOoHS':=jS';-F-AkNM8s#$RORNMOODF	RRRRRRRRRRRR#
SHNoMDbSk8CN0S#:S0D8_FOoHS':=jS';-F-AkNM8s#$RORNMkNb80RCRRRRRRRRRR#
SHNoMD8S#H:SSS8#0_oDFH:OS=''j;-S-AMFk8$NsRN#OMCR#sDHNR08NNMRHR
RRSo#HMSNDlCF8S#:S0D8_FOoHS':=jS';-F-AkNM8s#$RORNMlCF8RRRRRRRRRRRRR#
SHNoMDHSExS_L:0S#8F_DoSHO:4=''-;S-kAFMs8N$OR#NaMRs0H#NR0CO0FMsRFD
SS
#MHoNEDSF,D8FHCbMN,b8MFC,8bNF,k0bHN8MSS:#_08DHFoOS;

HS#oDMNSoMC_H0so#:S0D8_FOoH;#
SHNoMDkSbDkD_bSS:#_08DHFoOS;
#MHoNbDSHOM_L:H0S8#0_oDFHPO_CFO0sR568MFI0jFR2S;

oLCHSM

CSMos_0H<oS=mSa_71apQmtBhS5 at_)tQt ;)2
HSbML_OH<0S=mSa_71apQmtBBe aSm)5huQ_uaY 
2;SDbkDb_kS=S<S_am1pa7mBtQSz5upupz2
;
SOHMDM	_SR<=SuQhzBa_pGiRFMsRC0o_s;Ho
kSF0	OD_<MS=zSmaauz_iBpRsGFRoMC_H0soS;
HDMO	=S<SOHMDM	_R8NMRmBpB i_hpqA S;
FOk0D<	S=kSF0	OD_NMRMB8RpimB_q hA;p 
SS
E8FDSS<=pBqa]h_Qu_zaezqp S;
FHCbM=S<Samzu_za Ahqp
 ;Su
SqqBitu _QHh_Sb:SsCFO#5#SbFN8CRM,bFN8kR0,uiqBq_t u2Qh
CSLo
HMSNSb8SHM<u=SqqBitu _Q
h;SVSHSN5b8MFC=''42ER0CSM
SqSuBtiq Q_uh=S<S''Z;S
SCCD#
SSSuiqBq_t uSQh<b=SNk8F0S;
S8CMR;HV
MSC8sRbF#OC#S;

pStmpAq_wAzw_ )muzaz<aS=NSb8;HM
----------------------------------------------------------------
-S
sSbCF_H_:HSSCbs_
HFSsbF0NRlb
S5SSSSE8FDSS=>E8FD,S
SS#Ss0SHF='>Sj
',SSSSLC#_M>S=S_L#C
M,SSSS#VEH0>S=SH#EV
0,SSSS0	ODSS=>0	OD,S
SSMSHOSD	=H>SM	OD,S
SSkSF0	ODSS=>FOk0D
	,SSSSkNb80=CS>bSk8CN0,S
SSCSFbSHM=F>SCMbH,S
SS8S#H=SS>8S#HS,
SlSSFS8C=l>SF,8C
SSSSxEH_=LS>HSEx,_L
SSSSF#8S>S=SF#8,S
SSFS8kS04=7>S__Qh4S,
S8SSFjk0SS=>7h_Q_
j,SSSS848sSS=>7z_ma,_4
SSSSs88j>S=Sm7_zja_,S
SSNSb8SHM=b>SNM8H,S
SSNSb80FkSS=>bFN8k
0,SSSSbFN8C=MS>NSb8MFC,S
SSLSOH=0S>HSbML_OHS0
S2SS;M
C8AS1__tAQem_;-

----------------------------------------------------------------
S--SSSS1tA_A-
--------------------------------------------------------------
--
LDHs$NsRCHCCk;
#HCRC3CC#_08DHFoO4_4nNc3D
D;kR#CHCCC38#0_oDFHNO_sEH03DND;#
kCCRHC#C30D8_FOoH_#kMHCoM8D3ND-;
-LDHs$NsSsIF	k;
#ICSF3s	#_08DHFoOA_1aD3ND
;
CHM001$SAA_tS
H#
sbF0
S5SpStmpAq_wAzw_ )muzazSaSSF:Sk#0S0D8_FOoH;S
Sz)1 _t1Qh_qpatm_pqmApz_Aw)w SH:SM0S#8F_Do
HOS;S2
M
C8AS1_;tA
0N0skHL0#CR$LM_D	NO_GLFRRFV1tA_ARR:ObFlFMMC0#RHRk0sC
;
NEsOHO0C0CksS_1AteA_RRFV1tA_A#RH
oLCHSM
tApmqAp_z ww)z_maauzSS<=z)1 _t1Qh_qpatm_pqmApz_Aw)w ;M
C8AR1__tAe
;

D

HNLssH$RC;CC
Ck#RCHCC03#8F_Do_HO4c4n3DND;#
kCCRHC#C30D8_FOoH_HNs0NE3D
D;kR#CHCCC38#0_oDFHkO_Mo#HM3C8N;DD
M
C0$H0S_1AWvq)AammS
H#b0FsSS5
SmAmaSS:H#MS0D8_FOoH;S
S1S4S:MSHS8#0_oDFH
O;SjS1SSS:H#MS0D8_FOoH;S
S2
;
CRM81WA_qA)vm;ma
0N0skHL0#CR$LM_D	NO_GLFRRFV1WA_qA)vmRma:FROlMbFCRM0H0#Rs;kC
0N0skHL0#CR$MM_FkbsMFCRVAR1_)WqvmAmaRR:ObFlFMMC0#RHRk0sC
;
---------------------------------------------------------
---S-SSAS1__Qm7-1
---------------------------------------------------------
--
LDHs$NsRCHCCk;
#HCRC3CC#_08DHFoO4_4nNc3D
D;kR#CHCCC38#0_oDFHNO_sEH03DND;#
kCCRHC#C30D8_FOoH_#kMHCoM8D3ND-;
-LDHs$NsSsIF	k;
#ICSF3s	#_08DHFoOA_1aD3ND
;
S7--HCVVs0CMHRND#MHoNMDHomRQ
0CMHS0$1QA_m1_7S
H#SMoCCOsHSS5
S Sht)_aQ tt)RR:LSH0SSSSSS:=';j'
SSSu_Qha YuSL:RHP0_CFO0s6R5RI8FMR0Fj:2S=jS"jjjjj
";SQSSma_1qqh7):7SRs#0HSMoSSSS:"=S1pA_e_71muzaz
a"S2SS;S

b0FsSS5
S_S7m_za4SSS:MSHS8#0_oDFHSO;-Q-RM0bkR0FkbRk04SR
S_S7m_zajSSS:MSHS8#0_oDFHSO;-Q-RM0bkR0FkbRk0jSR
SpSBm_Bi Ahqp: SSSHM#_08DHFoO-;S-DRBFRO	CLMNDRC#hR W-FROlMlFRR0FHFM/kO0RD	FO#SR
S_S7Q4h_S:SSS0FkS8#0_oDFHSO;-m-Rkk0b0MRHbRk04S
SSQ7_hS_jSSS:FSk0#_08DHFoO-;S-kRm00bkRbHMkj0R
SSSmuzaz a_hpqA :SSRRHM#_08DHFoO=S:';]'SR--mkkb0M- NCLDRS
SSapqBQ]_hauz_peqz: SSSHM#_08DHFoO-;S-MRQbRk0O0FMsRFD
SSSQzhuap_Bi:SSSSHM#_08DHFoO-;S-MRQbRk0OODF	SR
SzSmaauz_iBpSSS:H#MS0D8_FOoH;-RR-kRm00bkRFODOS	
SqSuBtiq Q_uh:SSSFHMk#0S0k8_DHFoO-;S-#RzC#s'RObN	CNoRMbHR'-Ru'q7R0FkbRk0RS
SSBuqi qt_huQ_:ASSFHMk#0S0k8_DHFoO-S-RCz#sR'#b	NONRoCbRHM-uR'qR7'Fbk0kR0R
SSS2
;
CRM81QA_m1_7;0
N0LsHkR0C#_$MLODN	F_LGVRFR_1AQ7m_1RR:ObFlFMMC0#RHRk0sC
;
NEsOHO0C0CksR_1AQ7m_1R_eF1VRAm_Q_R71HS#
-#-SHNoMD-#
--------------------
HS#oDMNSOHMDM	_,0FkO_D	MM,HO,D	FOk0D#	,8:FSS8#0_oDFH
O;S#
SHNoMD#SL_SCM:0S#8F_DoSHO:j=''-;S-kAFMs8N$OR#NCMRMDNLCRRRRRRRRRRR
HS#oDMNSH#EV:0SS8#0_oDFH:OS=''j;-S-AMFk8$NsRN#OMER#HRV0RRRRRRRRR
RRSo#HMSND0	ODS#:S0D8_FOoHS':=jS';-F-AkNM8s#$RORNMOODF	RRRRRRRRRRRR#
SHNoMDbSk8CN0S#:S0D8_FOoHS':=jS';-F-AkNM8s#$RORNMkNb80RCRRRRRRRRRR#
SHNoMD8S#H:SSS8#0_oDFH:OS=''j;-S-AMFk8$NsRN#OMCR#sDHNR08NNMRHR
RRSo#HMSNDlCF8S#:S0D8_FOoHS':=jS';-F-AkNM8s#$RORNMlCF8RRRRRRRRRRRRR#
SHNoMDHSExS_L:0S#8F_DoSHO:4=''-;S-kAFMs8N$OR#NaMRs0H#NR0CO0FMsRFD
SS
#MHoNEDSF,D8FHCbMSS:#_08DHFoO-;S-CaERJsCkCHs8NRbOo	NCHRbM$R0blCRkR#0L#CRCI0RERCMHlF_NFOsRRH#H0M#NHM0N80C3#
SHNoMDNSb8MFC,NRb80Fk,NRb8SHM:0S#8F_Do;HO
SS
#MHoNbDSHOM_L:H0S8#0_oDFHPO_CFO0sR568MFI0jFR2S;
#MHoNMDSC0o_s:HoS8#0_oDFH
O;S-
S-FSOlMbFCRM0b_sCHSF
ObFlFMMC0sSbCF_H
FSbs50S
SSSE8FDSH:SM#RS0D8_FOoH;S
SS0s#H:FSSSHM#_08DHFoOS;
S#SL_SCM:MSHS8#0_oDFH
O;S#SSE0HVSH:SM0S#8F_Do;HO
SSS0	ODSH:SM0S#8F_Do;HO
SSSHDMO	SS:H#MS0D8_FOoH;S
SS0FkOSD	:MSHS8#0_oDFH
O;SkSSb08NCSS:H#MS0D8_FOoH;S
SSbFCH:MSSSHM#_08DHFoOS;
S8S#H:SSSSHM#_08DHFoOS;
SFSl8:CSSSHM#_08DHFoOS;
SHSExS_L:MSHS8#0_oDFH
O;S#SS8SFS:kSF00S#8F_Do;HO
SSS80Fk4SS:FSk0#_08DHFoOS;
SFS8kS0j:kSF00S#8F_Do;HO
SSS848sSH:SM0S#8F_Do;HO
SSS8j8sSH:SM0S#8F_Do;HO
SSSbHN8MSS:H#MS0D8_FOoH;S
SS8bNFSk0:kSF00S#8F_Do;HO
SSSbFN8C:MSS0FkS8#0_oDFH
O;SOSSLSH0:MSHS8#0_oDFHPO_CFO0s6S5RI8FMR0FjS2
S;S2
MSC8FROlMbFC;M0
C
Lo
HMSoMC_H0so=S<S_am1pa7mBtQS 5ht)_aQ tt)
2;SMbH_HOL0=S<S_am1pa7mBtQea Bm5)Su_Qha Yu2S;

H
SM	OD_<MS=QRShauz_iBpRsGFRoMC_H0soS;
FOk0DM	_SS<=muzazBa_pGiRFMsRC0o_s;Ho
MSHOSD	<H=SM	OD_NMRMB8RpimB_q hA;p 
kSF0	ODSS<=FOk0DM	_R8NMRmBpB i_hpqA S;

FSED<8S=qSpa_B]Qzhuaq_ep;z 
CSFbSHM<m=Szzauah_ q Ap;

SSBuqi qt_huQ_:HSSFbsO#C#SN5b8MFC,NRb80Fk2L
SCMoH
HSSVbS5NC8FM4=''02RE
CMSuSSqqBitu _Q<hS=ZS''S;
S#CDCS
SSBuqi qt_huQSS<=bFN8k
0;SMSC8VRH;C
SMb8RsCFO#
#;Sb
SNM8HRR<=uiqBq_t uRQh;

SSBuqi qt_huQ_HA_Sb:SsCFO#5#SbFN8CRM,bFN8k
02SoLCHSM
SSHV58bNF=CM'24'RC0EMS
SSBuqi qt_huQ_<AS=ZS''S;
S#CDCS
SSBuqi qt_huQ_<AS=FSM0NRb80Fk;S
SCRM8H
V;S8CMRFbsO#C#;S

E8FDSR<=pBqa]h_Qu_zaezqp S;
FHCbM<RS=zRmaauz_q hA;p 
-
-SCbs__HFHb
SsHC_FS_H:sSbCF_H
FSbsl0RN5bS
SSSSDEF8>S=SDEF8S,
SsSS#F0HSS=>',j'
SSSS_L#C=MS>#SL_,CM
SSSSH#EV=0S>ES#H,V0
SSSSD0O	>S=SD0O	S,
SHSSM	ODSS=>HDMO	S,
SFSSkD0O	>S=S0FkO,D	
SSSS8kbNS0C=k>Sb08NCS,
SFSSCMbHSS=>FHCbMS,
S#SS8SHS=#>S8
H,SSSSlCF8SS=>lCF8,S
SSHSExS_L=E>SHLx_,S
SS8S#F=SS>8S#FS,
S8SSF4k0SS=>7h_Q_
4,SSSS80Fkj>S=SQ7_h,_j
SSSSs884>S=Sm7_z4a_,S
SS8S8s=jS>_S7m_zajS,
SbSSNM8HSS=>bHN8MS,
SbSSNk8F0>S=S8bNF,k0
SSSS8bNFSCM=b>SNC8FMS,
SOSSLSH0=b>SHOM_L
H0SSSS2
;
CRM81QA_m1_7_
e;
--------------------------------------------------------------
-SSSShSt7-
----------------------------------------------------------
--
LDHs$NsRCHCCk;
#HCRC3CC#_08DHFoO4_4nNc3D
D;kR#CHCCC38#0_oDFHNO_sEH03DND;#
kCCRHC#C30D8_FOoH_#kMHCoM8D3ND
;
CHM00t$ShH7S#F
bs50S
YSSSF:Sk#0S0D8_FOoH
2SS;C

Mt8Rh
7;Ns00H0LkC$R#MD_LN_O	LRFGFtVRh:7RRlOFbCFMMH0R#sR0k
C;
ONsECH0Os0kChRt7R_eFtVRhH7R#C
Lo
HMS<YS=jS''C;
Mt8Rhe7_;-

------------------------------------------------------------
S--SSSSe
BB-------------------------------------------------------------D

HNLssH$RC;CC
Ck#RCHCC03#8F_Do_HO4c4n3DND;#
kCCRHC#C30D8_FOoH_HNs0NE3D
D;kR#CHCCC38#0_oDFHkO_Mo#HM3C8N;DD
M
C0$H0SBeBS
H#b0FsSS5
S:YSS0FkS8#0_oDFHSO
S
2;
8CMRBeB;0
N0LsHkR0C#_$MLODN	F_LGVRFRBeBRO:RFFlbM0CMRRH#0Csk;N

sHOE00COkRsCe_BBeVRFRBeBR
H#LHCoMY
SSS<=';4'
8CMRBeB_
e;
-
----------------------------------------------------------
---S-SSRSRu_ppB m)S-
----------------------------------------------------------
--DsHLNRs$Q   ;#
kC RQ 1 3ap7_mBtQ_n44cD3NDk;
#QCR 3  1_a7pQmtBh_z1hQt N73D
D;kR#CQ   38#0_oDFHNO_sEH03DND;1
z  RQ M 3kslCH#O_0q83p
p;
0CMHR0$#bL_DOD_FRsCH
#
RCRoMHCsO
R5SSRR)  w)B h p_Bi)_w  TzhRBYSH:RMo0CCSsR:j=R;SR
Spupm_zawT) zB hYSRS:MRH0CCos:RS=jR4jS;
S w 7BAqiq_uaR]SS:SSRs#0HRMoR=S:RH"#lCbD"
;SS S7p_qYqz7K1 avhva_mR7 SRS:#H0sMRoRSR:="M8$NOlH"
;RSQSwX_ 77q pY7_qKaz1va hR:SSR0HMCsoCR:RS=;RjRS
S AhqpQ _Bq taS RS:SSR0LHR:SS=jR''S;
Spupm_zau1]q SSSS#:R0MsHo:RS=MS"F"MC;S
S7wQeSSSSSRS:L_H0P0COF6s5RI8FMR0Fj
2;SQS7eS)SSSSS:HRL0C_POs0F58dRF0IMF2Rj;S
S7TQeSSSSSRS:L_H0P0COF.s5RI8FMR0Fj
2;SQSwp)a _h)qtS SSSSS:HRL0C_POs0F58.RF0IMF2RjRSR
S8--Cs0ClCHMRV8CN0kDRDPNk
C#S-S-7)QeSSSSSRS:L_H0P0COFds5RI8FMR0Fj:2R=jR"j"jj2R;
RRRRR;R2
bRRFRs05RR
RRRRR)RR )w   hBBSpiSH:RM0R#8F_Do;HO
RRRRRRRRpupmBzamS) SRS:FRk0#_08DHFoOR;
RRRRRuRRpzpmamtpASqpSF:Rk#0R0D8_FOoH;R
RRRRRRXR a w 7BAqiSSS:MRHR8#0_oDFH
O;SRSR7qYhv7QB YpqSRS:H#MR0D8_FOoH_OPC0RFs58dRF0IMF2RjRR;
RRRRRARRY1uq1SSSSH:RM0R#8F_Do;HO
RRRRRRRR1)  SaSSRS:H#MR0D8_FOoH;R
RRRRRR7R1mSSSSF:Rk#0R0D8_FOoH;R
RRRRRR7R1QSSSSH:RM0R#8F_Do;HO
RRRRRRRRp1BiSSSSH:RM0R#8F_Do;HO
RRRRRRRRBpmiSSSSH:RM0R#8F_Do;HO
RRRRRRRRapqBh]Quezaq pzSRS:H#MR0D8_FOoH
RRRRRRR2R;
RM
C8LR#_DbD_sOFC
;
NEsOHO0C0CksR_#Lb_DDOCFs_ONsEVRFR_#Lb_DDOCFsR
H#LHCoMCR
M#8RLD_bDF_OsNC_s;OE
0N0skHL0#CR$LM_D	NO_GLFRRFV#bL_DOD_FRsC:FROlMbFCRM0H0#Rs;kC
-
----------------------------------------------------------
---S-SSuSSpup_q-7
------------------------------------------------------------
LDHs$NsR Q  k;
#QCR 3  1_a7pQmtB4_4nNc3D
D;kR#CQ   371a_tpmQzB_ht1Qh3 7N;DD
Ck#R Q  03#8F_Do_HON0sHED3NDz;
1Q R 3  MCkls_HO#308q;pp
M
C0$H0R_#Lb_DDbRN8H
#
RCRoMHCsO
R5SSRR)  w)B h p_Bi)_w  TzhRBYSH:RMo0CC:sR=;RjR-
S-)RR )w   hB_iBp_e7QQ_7 ASYR:MRH0CCos=R:R
4;SR--Rw)  h) BB _pvi_zQpau_pYASYR:MRH0CCos=R:RR4;SSS
Spupm_zawT) zB hYSRS:MRH0CCos=R:Rj4j;S
Sw7  AiqB_auq]SRSSRS:#H0sMRoR:"=R#bHlD;C"SS
S7q pY7_qKaz1va h_7vm SRS:0R#soHMR=R:R$"8MHNlOR";
wSSQ7X _p7 qqY_71Kzahv aSRS:MRH0CCos:RR=;RjRS
S AhqpQ _Bq taS RS:SSR0LHR:SS=jR''S;
Spupm_zau1]q SSSS#:R0MsHo:RS=MS"F"MC;S
S7wQeSSSSSRS:L_H0P0COF6s5RI8FMR0Fj
2;SQS7eS)SSSSS:HRL0C_POs0F58dRF0IMF2Rj;S
S7TQeSSSSSRS:L_H0P0COF.s5RI8FMR0Fj
2;SQSwp)a _h)qtS SS:SSR0LH_OPC05Fs.FR8IFM0RRj2RS
S-C-80lCsHRMC8NCVkRD0PkNDCR#
RRRRR;R2
bRRFRs05RR
RRRRRuRRqqBitQ uh:SSRRHM#_08DHFoOR;
RRRRRuRRpzpma)Bm SSS:kRF00R#8F_Do;HO
RRRRRRRRpupmtzapqmAp:SSR0FkR8#0_oDFH
O;RRRRRRRR wXa A 7qSBiSRS:H#MR0D8_FOoH;S
SRYR7hQqvBp7 qSYS:MRHR8#0_oDFHPO_CFO0sdR5RI8FMR0Fj;2R
RRRRRRRRuAYqS11S:SSRRHM#_08DHFoOR;
RRRRR)RR a1 SSSS:MRHR8#0_oDFH
O;RRRRRRRR1S7mS:SSR0FkR8#0_oDFH
O;RRRRRRRR1S7QS:SSRRHM#_08DHFoOR;
RRRRR1RRBSpiS:SSRRHM#_08DHFoOR;
RRRRRpRRmSBiS:SSRRHM#_08DHFoOR;
RRRRRpRRq]aBQzhuapeqzS S:MRHR8#0_oDFHRO
RRRRR;R2

RRCRM8#bL_DbD_N
8;Ns00H0LkC$R#MD_LN_O	LRFGF#VRLD_bDN_b8RR:ObFlFMMC0#RHRk0sC
;
NEsOHO0C0CksR_#Lb_DDb_N8NEsORRFV#bL_DbD_NH8R#C
LoRHM
8CMR_#Lb_DDb_N8NEsO;0
N0LsHkR0C#_$MLODN	F_LGVRFR_#Lb_DDb_N8NEsORO:RFFlbM0CMRRH#0Csk;-

------------------------------------------------------------
S--SSSSu_pp.q_u7-
----------------------------------------------------------
--DsHLNRs$Q   ;#
kC RQ 1 3ap7_mBtQ_n44cD3NDk;
#QCR 3  1_a7pQmtBh_z1hQt N73D
D;kR#CQ   38#0_oDFHNO_sEH03DND;1
z  RQ M 3kslCH#O_0q83p
p;
0CMHR0$#bL_D.D__8bNR
H#
oRRCsMCH5OR
RSRSw)  h) BB _pwi_)z T YhBRRS:HCM0oRCs:j=R;SR
-)-S )w   hB_iBp_e7QQ_7 ASYR:MRH0CCos=R:R
4;SS--)  w)B h p_Biz_vpuaQpAY_Y:RSR0HMCsoCRR:=4S;RS-
S-pSupamz_)umawq_)z T YhBRRH#NNDI$=#RRw) BRpiVJsCkOCM$S
Sumppzua_mA)a_ w)Thz BSYRSH:RMo0CC:sR=jR4jS;
S w 7BAqiq_uaS]RS:SSRs#0HRMoRR:="l#Hb"DC;SS
Sp7 qqY_71Kzahv am_v7S RS#:R0MsHo:RR=8R"$lMNH;O"RS
Sw QX7 _7p_qYqz7K1 avhSaRSH:RMo0CCRsR:j=R;SR
Sq hA_p QtB qRa SSSS:HRL0=R:R''j;S
Sumppzua_] q1SSSSR:RRRs#0HRMoSS:="MMFC
";SQS7eSwSSSSS:HRL0C_POs0F586RF0IMF2Rj;S
S7)QeSSSSSRS:L_H0P0COFds5RI8FMR0Fj
2;SQS7eSTSSSSS:HRL0C_POs0F58.RF0IMF2Rj;S
SwaQp ))_q htRRRRRRRRRSRSSL:RHP0_CFO0sR5.8MFI0jFR2
RRS-S-8CC0sMlHCCR8VDNk0NRPD#kC
RRRRRRR2R;
RsbF0RR5
RRRRRRRRBuqi qtuSQhSRS:H#MR0D8_FOoH;R
RRRRRRpRupamzB m)qSSS:kRF00R#8F_Do;HO
RRRRRRRRpupmtzapqmApSqS:kRF00R#8F_Do;HO
RRRRRRRRpupmBzamA) S:SSR0FkR8#0_oDFH
O;RRRRRRRRumppzpatmpAqA:SSR0FkR8#0_oDFH
O;RRRRRRRR wXa A 7qSBiSRS:H#MR0D8_FOoH;S
SRYR7hQqvBp7 qSYS:MRHR8#0_oDFHPO_CFO0sdR5RI8FMR0Fj;2R
RRRRRRRRuAYqS11S:SSRRHM#_08DHFoOR;
RRRRR)RR a1 SSSS:MRHR8#0_oDFH
O;RRRRRRRR1S7mS:SSR0FkR8#0_oDFH
O;RRRRRRRR1S7QS:SSRRHM#_08DHFoOR;
RRRRR1RRBSpiS:SSRRHM#_08DHFoOR;
RRRRRpRRmSBiS:SSRRHM#_08DHFoOR;
RRRRRpRRq]aBQzhuapeqzS S:MRHR8#0_oDFHRO
RRRRR;R2

RRCRM8#bL_D.D__8bN;0
N0LsHkR0C#_$MLODN	F_LGVRFR_#Lb_DD.N_b8RR:ObFlFMMC0#RHRk0sC
;
NEsOHO0C0CksR_#Lb_DD.N_b8s_NOFERVLR#_DbD_b._NH8R#C
LoRHM
8CMR_#Lb_DD.N_b8s_NO
E;
