// pll.v

// Generated using ACDS version 13.0 156 at 2020.03.31.04:13:02

`timescale 1 ps / 1 ps
module pll (
		input  wire  clki,    //  clki.clk
		output wire  clko,    //  clko.clk
		output wire  clkop    //  clko.clk
	);
	assign clko = clki;
	pll_altpll_0 altpll_0 (
		.clk       (clki),    //       inclk_interface.clk
		.reset     (1'b0), // inclk_interface_reset.reset
		.read      (),            //             pll_slave.read
		.write     (),            //                      .write
		.address   (),            //                      .address
		.readdata  (),            //                      .readdata
		.writedata (),            //                      .writedata
		.c0        (clkop),    //                    c0.clk
		.areset    (),            //        areset_conduit.export
		.locked    (),            //        locked_conduit.export
		.phasedone ()             //     phasedone_conduit.export
	);

endmodule
