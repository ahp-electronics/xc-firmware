--
@ER--B$FbsEHo0OR52gR4g-cRRj.jd$R1MHbDO$H0ROQM
R--fN]C8:CsR#//$DMbH0OH$N/lb0DN.Uj4J4.b/blNb#Cs/DGHH/MGD/HLoCCMs/HOo_CMoCCMs/HOs_NlssI_38PEyf4R

--
----B-R RppXv)qd4.X7-R--
--DsHLNRs$HCCC;#
kCCRHC#C30D8_FOoH_n44cD3NDk;
#HCRC3CC#_08DHFoOH_#o8MC3DND;H
DLssN$MRkHl#H;#
kCMRkHl#H3FPOlMbFC#M03DND;C

M00H$)RXq.vdXR47HR#
RsbF0
R5RRRRRRRR7RumRRR:FRk0#_08koDFHRO;RRRRR
RRRRRRRRRR1RumRRR:FRk0#_08koDFH
O;
RRRRRRRRRqjR:RRRRHM#_08koDFH
O;RRRRRRRRqR4RRRR:H#MR0k8_DHFoOR;
RRRRRqRR.RRRRH:RM0R#8D_kFOoH;R
RRRRRRdRqRRRR:MRHR8#0_FkDo;HO
RRRRRRRRRqcR:RRRRHM#_08koDFH
O;RRRRRRRR7RRRRRR:H#MR0k8_DHFoOR;
RRRRR7RRuj)qRH:RM0R#8D_kFOoH;R
RRRRRRuR7)Rq4:MRHR8#0_FkDo;HO
RRRRRRRR)7uq:.RRRHM#_08koDFH
O;RRRRRRRR7qu)dRR:H#MR0k8_DHFoOR;
RRRRR7RRuc)qRH:RM0R#8D_kFOoH;R
RRRRRRBRWpRiR:MRHR8#0_FkDo;HORRRRRRRR
RRRRRRRRRW R:RRRRHM#_08koDFHRO
RRRRR;R2RCR
MX8R)dqv.7X4;s
NO0EHCkO0sXCR)dqv.7X4_FeRV)RXq.vdXR47HR#
RHS#oDMNRjIC,CRI4#,RFRj,#,F4Rj8F,FR84#:R0D8_FOoH;C
Lo
HMSm7uRR<=8RFjIMECRu57)Rqc=jR''C2RDR#C8;F4
uS1m=R<Rj#FRCIEMqR5cRR='2j'R#CDCFR#4S;
IRCj<W=R MRN8MR5Fq0Rc
2;S4ICRR<=WN RMq8RcR;
SRzj:qR)vX4n4
7RRRRRRRRRRRRRRRRRb0FsRblNRR57=7>R,jRqRR=>qRj,q=4R>4Rq,.RqRR=>qR.,q=dR>dRq,S
RSuS7)Rqj=7>Ruj)q,uR7)Rq4=7>Ru4)q,uR7)Rq.=7>Ru.)q,uR7)Rqd=7>Rud)q,SR
S SWRR=>I,CjRpWBi>R=RpWBi7,Ru=mR>FR8j1,Ru=mR>FR#j
2;R4SzR):Rqnv4XR47
RRRRRRRRRRRRRRRRsbF0NRlb7R5RR=>7q,Rj>R=R,qjRRq4=q>R4q,R.>R=R,q.RRqd=q>RdR,
S7SSuj)qRR=>7qu)j7,Ru4)qRR=>7qu)47,Ru.)qRR=>7qu).7,Rud)qRR=>7qu)d
,RSWSS >R=R4IC,BRWp=iR>BRWpRi,7Rum=8>RFR4,1Rum=#>RF;42
8CMRqX)vXd.4e7_;-

----RpB p)RXqcvnXR47-----H
DLssN$CRHC
C;kR#CHCCC38#0_oDFH4O_43ncN;DD
Ck#RCHCC03#8F_Do_HO#MHoCN83D
D;DsHLNRs$k#MHH
l;kR#Ck#MHHPl3ObFlFMMC0N#3D
D;
0CMHR0$Xv)qn4cX7#RH
bRRFRs05R
RRRRRRuR7mRRR:kRF00R#8D_kFOoH;RRRRRRRRR
RRRRRRuR1mRRR:kRF00R#8D_kFOoH;R

RRRRRqRRjRRRRH:RM0R#8D_kFOoH;R
RRRRRR4RqRRRR:MRHR8#0_FkDo;HO
RRRRRRRRRq.R:RRRRHM#_08koDFH
O;RRRRRRRRqRdRRRR:H#MR0k8_DHFoOR;
RRRRRqRRcRRRRH:RM0R#8D_kFOoH;R
RRRRRR6RqRRRR:MRHR8#0_FkDo;HO
RRRRRRRRR7RR:RRRRHM#_08koDFH
O;RRRRRRRR7qu)jRR:H#MR0k8_DHFoOR;
RRRRR7RRu4)qRH:RM0R#8D_kFOoH;R
RRRRRRuR7)Rq.:MRHR8#0_FkDo;HO
RRRRRRRR)7uq:dRRRHM#_08koDFH
O;RRRRRRRR7qu)cRR:H#MR0k8_DHFoOR;
RRRRR7RRu6)qRH:RM0R#8D_kFOoH;R
RRRRRRBRWpRiR:MRHR8#0_FkDo;HORRRRRRRR
RRRRRRRRRW R:RRRRHM#_08koDFHRO
RRRRR;R2RCR
MX8R)nqvc7X4;s
NO0EHCkO0sXCR)nqvc7X4_FeRV)RXqcvnXR47HR#
RHS#oDMNRjIC,CRI4I,RCR.,I,CdRj#F,FR#4#,RFR.,#,FdRj8F,FR848,RFR.,8:FdR8#0_oDFH
O;LHCoM7
Su<mR=8RRFIjRERCM5)7uq=6RR''jR8NMR)7uq=cRR''j2DRC#
CRSFS84ERIC5MR7qu)6RR='Rj'NRM87qu)cRR='24'R#CDCSR
S.8FRCIEM7R5u6)qR'=R4N'RM78Ruc)qR'=RjR'2CCD#RS
S8;Fd
uS1m=R<RFR#jERIC5MRq=6RR''jR8NMRRqc=jR''C2RDR#C
#SSFI4RERCM5Rq6=jR''MRN8cRqR'=R4R'2CCD#RS
S#RF.IMECR65qR'=R4N'RMq8RcRR='2j'R#CDCSR
Sd#F;I
SC<jR= RWR8NMRF5M06Rq2MRN8MR5Fq0Rc
2;S4ICRR<=WN RM58RMRF0qR62NRM8q
c;S.ICRR<=WN RMq8R6MRN8MR5Fq0Rc
2;SdICRR<=WN RMq8R6MRN8cRq;S
Rz:jRRv)q44nX7RR
RRRRRRRRRRRRRbRRFRs0lRNb5=7R>,R7RRqj=q>Rjq,R4>R=R,q4RRq.=q>R.q,Rd>R=R,qd
SRSS)7uq=jR>uR7),qjR)7uq=4R>uR7),q4R)7uq=.R>uR7),q.R)7uq=dR>uR7),qdRS
SSRW =I>RCRj,WiBpRR=>WiBp,uR7m>R=Rj8F,uR1m>R=Rj#F2R;
SRz4:qR)vX4n4
7RRRRRRRRRRRRRRRRRb0FsRblNRR57=7>R,jRqRR=>qRj,q=4R>4Rq,.RqRR=>qR.,q=dR>dRq,S
RSuS7)Rqj=7>Ruj)q,uR7)Rq4=7>Ru4)q,uR7)Rq.=7>Ru.)q,uR7)Rqd=7>Rud)q,SR
S SWRR=>I,C4RpWBi>R=RpWBi7,Ru=mR>FR841,Ru=mR>FR#4
2;R.SzR):Rqnv4XR47
RRRRRRRRRRRRRRRRsbF0NRlb7R5RR=>7q,Rj>R=R,qjRRq4=q>R4q,R.>R=R,q.RRqd=q>RdR,
S7SSuj)qRR=>7qu)j7,Ru4)qRR=>7qu)47,Ru.)qRR=>7qu).7,Rud)qRR=>7qu)d
,RSWSS >R=R.IC,BRWp=iR>BRWpRi,7Rum=8>RFR.,1Rum=#>RF;.2
zRSdRR:)4qvn7X4RR
RRRRRRRRRRRRRRFRbsl0RN5bR7>R=RR7,q=jR>jRq,4RqRR=>qR4,q=.R>.Rq,dRqRR=>q
d,RSSS7qu)j>R=R)7uqRj,7qu)4>R=R)7uqR4,7qu).>R=R)7uqR.,7qu)d>R=R)7uqRd,
SSSW= R>CRIdW,RBRpi=W>RB,piRm7uRR=>8,FdRm1uRR=>#2Fd;M
C8)RXqcvnX_47e
;
---
-HR1lCbDRv)qR0IHECR#bNNs0qCR7 7)1V1RFssRCRN8NRM8I0sHC-
-RsaNoRC0:HRXDGHM

--
LDHs$NsRCHCCk;
#HCRC3CC#_08DHFoO4_4nNc3D
D;kR#CHCCC38#0_oDFH#O_HCoM8D3NDD;
HNLssk$RMHH#lk;
#kCRMHH#lO3PFFlbM0CM#D3NDC;
M00H$qR)vW_)_H)R#R
RRCRoMHCsO
R5RRRRRRRRVHNlD:$RRs#0HRMo:"=RMCFM"R;
RRRRRIRRHE80RH:RMo0CC:sR=;R4RR
RRRRRR8RN8HsI8R0E:MRH0CCos=R:RRn;RRRRRRRRRR--LRHoCkMFoVERF8sRCEb0
RRRRRRRRb8C0:ERR0HMCsoCRR:=c
j;RRRRRRRRsk8F0C_soRR:LDFFCRNM:0=Rs;kCRRRRR-R-R#ENR0FkbRk0s
CoRRRRRRRRIk8F0C_soRR:LDFFCRNM:0=Rs;kCRRRRR-R-R#ENR0FkbRk0s
CoRRRRRRRR8_HMsRCo:FRLFNDCM=R:RDVN#RC;RRRRR-RR-NRE#NR80HNRM0bkRosC
RRRRRRRR8sN8ss_C:oRRFLFDMCNRR:=V#NDCR;RRRRR-E-RNs#RCRN8Ns88CR##s
CoRRRRRRRRI8N8sC_soRR:LDFFCRNMRR:=V#NDCRRRR-RR-NRE#sRIHR0CNs88CR##s
CoRRRRRRRR2R;
RbRRFRs05R
RRRRRR_R)7amzRF:Rk#0R0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2R;
RRRRRWRR_z7maRR:FRk0#_08DHFoOC_POs0F58IH04E-RI8FMR0Fj
2;RRRRRRRR)7q7)RR:H#MR0D8_FOoH_OPC05FsNs88I0H8ER-48MFI0jFR2R;
RRRRR7RRQRhR:MRHR8#0_oDFHPO_CFO0sH5I8-0E4FR8IFM0R;j2
RRRRRRRR7Wq7:)RRRHM#_08DHFoOC_POs0F58N8s8IH04E-RI8FMR0Fj
2;RRRRRRRRWR R:MRHR8#0_oDFHRO;RRRRR-R-RHIs0CCRMDNLCFRVsNRslR
RRRRRRpRBiRR:H#MR0D8_FOoH;RRRRRRR-O-RD	FORsVFRlsN,8RN8Rs,8
HMRRRRRRRR)B_mp:iRRRHM#_08DHFoOR;RR-R-R0FbRFODOV	RFssR_k8F0R
RRRRRR_RWmiBpRH:RM0R#8F_DoRHORRRR-F-RbO0RD	FORsVFR8I_F
k0RRRRRRRR2C;
MC8RM00H$qR)vW_)_
);
R--LODF	NRslsRNONE
sHOE00COkRsCLODF	N_slVRFRv)q__)W)#RH
0N0skHL0oCRCsMCNs0F_bsCFRs0:0R#soHM;0
N0LsHkR0CoCCMsFN0sC_sb0FsRRFVLODF	N_slRR:NEsOHO0C0CksRRH#"N7kDFRbsA0RD	FORv)qR0MFRb#kb0FsC$8RCR0,HCMVsMsHoCR1D0CORv)q"O;
FFlbM0CMRqX)vXd.4R7RRsbF0
R5RRRRRRRR7RumRRR:FRk0#_08koDFHRO;RRRRR
RRRRRRRRRR1RumRRR:FRk0#_08koDFH
O;
RRRRRRRRRqjR:RRRRHM#_08koDFH
O;RRRRRRRRqR4RRRR:H#MR0k8_DHFoOR;
RRRRRqRR.RRRRH:RM0R#8D_kFOoH;R
RRRRRRdRqRRRR:MRHR8#0_FkDo;HO
RRRRRRRRRqcR:RRRRHM#_08koDFH
O;RRRRRRRR7RRRRRR:H#MR0k8_DHFoOR;
RRRRR7RRuj)qRH:RM0R#8D_kFOoH;R
RRRRRRuR7)Rq4:MRHR8#0_FkDo;HO
RRRRRRRR)7uq:.RRRHM#_08koDFH
O;RRRRRRRR7qu)dRR:H#MR0k8_DHFoOR;
RRRRR7RRuc)qRH:RM0R#8D_kFOoH;R
RRRRRRBRWpRiR:MRHR8#0_FkDo;HORRRRRRRR
RRRRRRRRRW R:RRRRHM#_08koDFHRO
RRRRR;R2RCR
MO8RFFlbM0CM;F
OlMbFCRM0Xv)qn4cX7RRRb0FsRR5
RRRRR7RRuRmRRF:Rk#0R0k8_DHFoOR;RRRRRRRR
RRRRR1RRuRmRRF:Rk#0R0k8_DHFoO
;
RRRRRRRRqRjRRRR:H#MR0k8_DHFoOR;
RRRRRqRR4RRRRH:RM0R#8D_kFOoH;R
RRRRRR.RqRRRR:MRHR8#0_FkDo;HO
RRRRRRRRRqdR:RRRRHM#_08koDFH
O;RRRRRRRRqRcRRRR:H#MR0k8_DHFoOR;
RRRRRqRR6RRRRH:RM0R#8D_kFOoH;R
RRRRRRRR7RRRR:MRHR8#0_FkDo;HO
RRRRRRRR)7uq:jRRRHM#_08koDFH
O;RRRRRRRR7qu)4RR:H#MR0k8_DHFoOR;
RRRRR7RRu.)qRH:RM0R#8D_kFOoH;R
RRRRRRuR7)Rqd:MRHR8#0_FkDo;HO
RRRRRRRR)7uq:cRRRHM#_08koDFH
O;RRRRRRRR7qu)6RR:H#MR0k8_DHFoOR;
RRRRRWRRBRpiRH:RM0R#8D_kFOoH;RRRRRRRRR
RRRRRR RWRRRR:MRHR8#0_FkDo
HORRRRR2RR;
RRCRM8ObFlFMMC0V;
k0MOHRFMo_C0M_kln8c5CEb0:MRH0CCoss2RCs0kMMRH0CCos#RH
sPNHDNLCNRPDRR:HCM0oRCs:j=R;C
Lo
HMRNRPD=R:Rb8C0nE/cR;
RRHV5C58bR0ElRF8nRc2>URc2ER0CRM
RPRRN:DR=NRPDRR+4R;
R8CMR;HV
sRRCs0kMNRPDC;
Mo8RCM0_knl_cV;
k0MOHRFMo_C0D0CVFsPC_5d.80CbERR:HCM0o2CsR0sCkRsMHCM0oRCsHL#
CMoH
sRRCs0kMC58bR0ElRF8n;c2
8CMR0oC_VDC0CFPs._d;k
VMHO0FoMRCD0_CFV0P5Cs80CbERR:HCM0o;CsRGlNRH:RMo0CCRs2skC0sHMRMo0CCHsR#N
PsLHNDPCRN:DRR0HMCsoCRR:=jL;
CMoH
HRRV8R5CEb0Rl-RN>GR=2RjRC0EMR
RRNRPD=R:Rb8C0-ERRGlN;R
RCCD#
RRRRDPNRR:=80CbER;
R8CMR;HV
sRRCs0kMN5PD
2;CRM8o_C0D0CVFsPC;k
VMHO0FoMRCM0_kdl_.C58bR0E:MRH0CCoss2RCs0kMMRH0CCos#RH
sPNHDNLCNRPDRR:HCM0oRCs:j=R;C
Lo
HMRVRHRC58bR0E<c=RUMRN8CR8bR0E>nR42ER0CRM
RRRRPRND:4=R;R
RCRM8H
V;RCRs0MksRDPN;M
C8CRo0k_Ml._d;k
VMHO0FoMRCM0_k4l_nC58bR0E:MRH0CCoss2RCs0kMMRH0CCos#RH
sPNHDNLCNRPDRR:HCM0oRCs:j=R;C
Lo
HMRVRHRC58bR0E<4=RnMRN8CR8bR0E>2RjRC0EMR
RRPRRN:DR=;R4
CRRMH8RVR;
R0sCkRsMP;ND
8CMR0oC_lMk_;4n
MVkOF0HMCRo0M_C8C_8b50E#CHxRH:RMo0CC;sRRb8C0:ERR0HMCsoC2CRs0MksR0HMCsoCR
H#PHNsNCLDRMlH_x#HCRR:HCM0oRCs:j=R;C
Lo
HMRHRlMH_#x:CR=CR8b;0E
HRRV#R5HRxC<CR8b20ERC0EMR
RRHRlMH_#x:CR=HR#x
C;RMRC8VRH;R
RskC0slMRH#M_H;xC
8CMR0oC_8CM_b8C0
E;O#FM00NMRlMk_DOCDc_nRH:RMo0CC:sR=CRo0k_Mlc_n5b8C0;E2
MOF#M0N0CRDVP0FCds_.RR:HCM0oRCs:o=RCD0_CFV0P_Csd8.5CEb02O;
F0M#NRM0M_klODCD_Rd.:MRH0CCos=R:R0oC_lMk_5d.D0CVFsPC_2d.;F
OMN#0MD0RCFV0P_Cs4:nRR0HMCsoCRR:=o_C0D0CVFsPC5VDC0CFPs._d,.Rd2O;
F0M#NRM0M_klODCD_R4n:MRH0CCos=R:R0oC_lMk_54nD0CVFsPC_24n;0

$RbCF_k0L_k#0C$b_RncHN#Rs$sNRk5MlC_ODnD_cFR8IFM0RRj,I0H8ER-48MFI0jFR2VRFR8#0_oDFH
O;0C$bR0Fk_#Lk_b0$C._dRRH#NNss$MR5kOl_C_DDd8.RF0IMF,RjR8IH04E-RI8FMR0FjF2RV0R#8F_Do;HO
b0$CkRF0k_L#$_0b4C_n#RHRsNsN5$RM_klODCD_R4n8MFI0jFR,HRI8-0E4FR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNRksF0k_L#c_nRF:RkL0_k0#_$_bCnRc;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RVFR8k50RHkMb0FR0RH0s-N#002C#
o#HMRNDs0Fk_#Lk_Rd.:kRF0k_L#$_0bdC_.R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFRk8F0HR5M0bkRR0F0-sH#00NC
#2#MHoNsDRF_k0L_k#4:nRR0Fk_#Lk_b0$Cn_4;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFV80FkRM5HbRk000FRs#H-0CN0##2
HNoMDFRskC0_MRR:#_08DHFoOC_POs0F5lMk_DOCDc_nRI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-C-RMDNLCV#RF0sRs#H-0CN0#H
#oDMNRkIF0k_L#c_nRF:RkL0_k0#_$_bCnRc;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RVFR8k50RHkMb0FR0RH0s-N#002C#
o#HMRNDI0Fk_#Lk_Rd.:kRF0k_L#$_0bdC_.R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFRk8F0HR5M0bkRR0F0-sH#00NC
#2#MHoNIDRF_k0L_k#4:nRR0Fk_#Lk_b0$Cn_4;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFV80FkRM5HbRk000FRs#H-0CN0##2
HNoMDFRIkC0_MRR:#_08DHFoOC_POs0F5lMk_DOCDc_nRI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-C-RMDNLCV#RF0sRs#H-0CN0#H
#oDMNRksF0M_C_Rd.:0R#8F_Do;HO
o#HMRNDs0Fk__CM4:nRR8#0_oDFH
O;#MHoNIDRF_k0CdM_.RR:#_08DHFoO#;
HNoMDFRIkC0_Mn_4R#:R0D8_FOoH;H
#oDMNR0Is_RCM:0R#8F_Do_HOP0COFMs5kOl_C_DDn8cRF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RHIs0CCRMDNLCV#RFCsRNROEsRFIF)VRqOvRC#DD
o#HMRNDI_s0CdM_.RR:#_08DHFoO#;
HNoMDsRI0M_C_R4n:0R#8F_Do;HO
o#HMRNDHsM_C:oRR8#0_oDFHPO_CFO0sH5I8-0E4FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-#RkC08RFCRso0H#C7sRQ
hR#MHoNsDRF_k0sRCo:0R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-#RkC08RFCRso0H#C7sRm
za#MHoNIDRF_k0sRCo:0R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-#RkC08RFCRso0H#C7sRm
za#MHoNsDRNs8_C:oRR8#0_oDFHPO_CFO0s85N8HsI8-0E4FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-#RkC08RFCRso0H#CqsR7
7)#MHoNIDRNs8_C:oRR8#0_oDFHPO_CFO0s85N8HsI8-0E4FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-#RkC08RFCRso0H#CqsR7
7)#MHoNDDRFsI_Ns88R#:R0D8_FOoH_OPC05Fs6FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-8RN8LsRHR0#HkMb0FR0Rv)qRDOCD5#RcHRL0s#RCHJks2C8
o#HMRNDD_FII8N8sRR:#_08DHFoOC_POs0F586RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-N-R8R8sL#H0RbHMk00RFqR)vCRODRD#5LcRHR0#skCJH8sC20
N0LsHkR0C\N3slV_FV0#C\RR:#H0sM
o;
oLCH
M
RRRR-Q-RV8RN8HsI8R0E<RR6NH##o'MRj0'RFMRkk8#CR0LH#R
RRjRzRRR:H5VRNs88I0H8ERR=4o2RCsMCN
0CRRRRRRRRD_FIs8N8s=R<Rj"jj"jjRs&RNs8_Cjo52R;
RRRRRDRRFII_Ns88RR<="jjjjRj"&NRI8C_so25j;R
RRMRC8CRoMNCs0zCRjR;
RzRR4:RRRRHV58N8s8IH0=ERRR.2oCCMsCN0
RRRRRRRRIDF_8sN8<sR=jR"j"jjRs&RNs8_C4o5RI8FMR0Fj
2;RRRRRRRRD_FII8N8s=R<Rj"jjRj"&NRI8C_soR548MFI0jFR2R;
RCRRMo8RCsMCNR0Cz
4;RRRRzR.R:VRHR85N8HsI8R0E=2RdRMoCC0sNCR
RRRRRRFRDIN_s8R8s<"=Rj"jjRs&RNs8_C.o5RI8FMR0Fj
2;RRRRRRRRD_FII8N8s=R<Rj"jj&"RR8IN_osC58.RF0IMF2Rj;R
RRMRC8CRoMNCs0zCR.R;
RzRRd:RRRRHV58N8s8IH0=ERRRc2oCCMsCN0
RRRRRRRRIDF_8sN8<sR=jR"j&"RR8sN_osC58dRF0IMF2Rj;R
RRRRRRFRDIN_I8R8s<"=RjRj"&NRI8C_soR5d8MFI0jFR2R;
RCRRMo8RCsMCNR0Cz
d;SSzc:VRHR85N8HsI8R0E=2R6RMoCC0sNCS
SD_FIs8N8s=R<R''jRs&RNs8_Cco5RI8FMR0Fj
2;SFSDIN_I8R8s<'=Rj&'RR8IN_osC58cRF0IMF2Rj;C
SMo8RCsMCNR0Cz
c;RRRRzR6R:VRHR85N8HsI8R0E>2R6RMoCC0sNCR
RRRRRRFRDIN_s8R8s<s=RNs8_C6o5RI8FMR0Fj
2;RRRRRRRRD_FII8N8s=R<R8IN_osC586RF0IMF2Rj;R
RRMRC8CRoMNCs0zCR6
;
RRRR-Q-RV8R5HsM_CRo2sHCo#s0CRh7QRHk#MBoRpRi
RzRRn:RRRRHV5M8H_osC2CRoMNCs0RC
RRRRRbRRsCFO#5#RB,piRh7Q2CRLo
HMRRRRRRRRRRRRH5VRBRpi=4R''MRN8pRBiP'CC2M0RC0EMR
RRRRRRRRRRRRRRMRH_osCRR<=7;Qh
RRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMRFbsO#C#;R
RRMRC8CRoMNCs0zCRnR;
RzRR(:RRRRHV50MFRM8H_osC2CRoMNCs0RC
RRRRRRRRRHRRMC_so=R<Rh7Q;R
RRMRC8CRoMNCs0zCR(
;
RRRR-Q-RV8R5F_k0s2CoRosCHC#0smR7zkaR#oHMRpmBiR
RRURzs:RRRRHV5Fs8ks0_CRo2oCCMsCN0
RRRRRRRRFbsO#C#R_5)miBp,FRsks0_CRo2LHCoMR
RRRRRRRRRRVRHR_5)miBpR'=R4N'RM)8R_pmBiP'CC2M0RC0EMR
RRRRRRRRRRRRRR_R)7amzRR<=s0Fk_osC;R
RRRRRRRRRRMRC8VRH;R
RRRRRRMRC8sRbF#OC#R;
RCRRMo8RCsMCNR0Cz;Us
RRRRszgRRR:H5VRMRF0sk8F0C_soo2RCsMCN
0CRRRRRRRRRRRR)m_7z<aR=FRsks0_C
o;RRRRCRM8oCCMsCN0Rszg;R

R-RR-VRQRF58ks0_CRo2sHCo#s0CRz7ma#RkHRMomiBp
RRRRIzURRR:H5VRIk8F0C_soo2RCsMCN
0CRRRRRRRRbOsFCR##5mW_B,piRkIF0C_soL2RCMoH
RRRRRRRRRRRRRHV5mW_BRpi=4R''MRN8_RWmiBp'CCPMR020MEC
RRRRRRRRRRRRRRRR7W_mRza<I=RF_k0s;Co
RRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMRFbsO#C#;R
RRMRC8CRoMNCs0zCRU
I;RRRRzRgIRH:RVMR5FI0R80Fk_osC2CRoMNCs0RC
RRRRRRRRRWRR_z7ma=R<RkIF0C_soR;
RCRRMo8RCsMCNR0Cz;gI
R
RR-R-RRQV58N8sC_sos2RC#oH0RCsq)77RHk#MBoRpRi
RzRR4RjR:VRHRN5s8_8ss2CoRMoCC0sNCR
RRRRRRsRbF#OC#)R5_pmBi),Rq)772CRLo
HMRRRRRRRRRRRRH5VR)B_mp=iRR''4R8NMRm)_B'piCMPC002RE
CMRRRRRRRRRRRRRRRRs_N8sRCo<)=Rq)7758N8s8IH04E-RI8FMR0Fj
2;RRRRRRRRRRRRCRM8H
V;RRRRRRRRCRM8bOsFC;##
RRRR8CMRMoCC0sNC4RzjR;
RzRR4:4RRRHV50MFR8sN8ss_CRo2oCCMsCN0
RRRRRRRRRRRR8sN_osCRR<=)7q7)R;
RCRRMo8RCsMCNR0Cz;44
R
RR-R-RRQV58N8sC_sos2RC#oH0RCsq)77RHk#MBoRpRi
RzRR4R.R:VRHRN5I8_8ss2CoRMoCC0sNCR
RRRRRRsRbF#OC#BR5pRi,W7q7)L2RCMoH
RRRRRRRRRRRRRHV5iBpR'=R4N'RMB8RpCi'P0CM2ER0CRM
RRRRRRRRRRRRRIRRNs8_C<oR=qRW757)Ns88I0H8ER-48MFI0jFR2R;
RRRRRRRRRCRRMH8RVR;
RRRRRCRRMb8RsCFO#
#;RRRRCRM8oCCMsCN0R.z4;R
RR4RzdRR:H5VRMRF0I8N8sC_soo2RCsMCN
0CRRRRRRRRRRRRI_N8sRCo<W=Rq)77;R
RRMRC8CRoMNCs0zCR4
d;RRRRRRRR
RRRRR--tCCMsCN0RC0ERv)qRDOCDN#RM#8RCODC0FRDo
HORRRRzR4c:FRVsRRHH5MRM_klODCD_Rnc-2R4RI8FMR0FjCRoMNCs0RC
R-RR-VRQR85N8HsI8R0E>2R6RCMC8FR0RCOsNR0CI0sHCMRCNCLDR8NMR0FkbRk0CLMND#CRCODC0FRDo
HORRRRRRRRzR46:VRHR85N8HsI8R0E>2RnRMoCC0sNCR
RRRRRRRRRRRRRRFRskC0_M25HRR<='R4'IMECRN5s8C_so85N8HsI8-0E4FR8IFM0RRn2=2RHR#CDCjR''R;
RRRRRRRRRRRRRIRRF_k0CHM52=R<R''4RCIEMIR5Ns8_CNo58I8sHE80-84RF0IMF2RnRH=R2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0CHM52=R<RRW IMECRN5I8C_so85N8HsI8-0E4FR8IFM0RRn2=2RHR#CDCjR''R;
RRRRRCRRMo8RCsMCNR0Cz;46
RRRRR--Q5VRNs88I0H8E=R<RR62MIFRsCH0RNCMLRDCFFsRkk0b0MRCNCLDRD#CCRO0DHFoOCRMC88C
RRRRRRRRnz4RH:RVNR58I8sHE80RR<=no2RCsMCN
0CRRRRRRRRRRRRRRRRs0Fk_5CMH<2R=4R''R;
RRRRRRRRRRRRRIRRF_k0CHM52=R<R''4;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R R;
RRRRRCRRMo8RCsMCNR0Cz;4n
RRRRR--tCCMsCN0RC0ERv)qRDOCDN#RM08Rs#H-0CN0#R
RRRRRR4Rz(RR:VRFs[MRHRH5I8R0E-2R4RI8FMR0FjCRoMNCs0RC
RRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)RzqcvnRD:RNDLCRRH#"a17"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloHC5*2ncR"&RW&"RR0HMCsoC'NHlo[C52RR&"R "&MRH0CCosl'HN5oCo_C0C_M880CbEH55+*42nRc,80CbER22&XR""RR&HCM0o'CsHolNC+5[4
2;RRRRRRRRRRRRLHCoMR
RRRRRRRRRR)RzqcvnRX:R)nqvc7X4RR
RRRRRRRRRRRRRRFRbsl0RN5bR7>R=R_HMs5Co[R2,q=jR>FRDIN_I858sjR2,q=4R>FRDIN_I858s4R2,q=.R>FRDIN_I858s.
2,RRRRRRRRRRRRRRRRRRRRRRRRRdRqRR=>D_FII8N8s25d,cRqRR=>D_FII8N8s25c,6RqRR=>D_FII8N8s256,SR
SSSSS7RRuj)qRR=>D_FIs8N8s25j,uR7)Rq4=D>RFsI_Ns885,42R)7uq=.R>FRDIN_s858s.
2,SSSSSRSR7qu)d>R=RIDF_8sN8ds527,Ruc)qRR=>D_FIs8N8s25c,uR7)Rq6=D>RFsI_Ns885,62RS
SSSSSR RWRR=>I_s0CHM52W,RBRpi=B>RpRi,7Rum=s>RF_k0L_k#nHc5,,[2Rm1uRR=>I0Fk_#Lk_5ncH2,[2R;
RRRRRRRRRRRRRsRRF_k0s5Co[<2R=FRskL0_kn#_c,5H[I2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRkIF0C_so25[RR<=I0Fk_#Lk_5ncH2,[RCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRCRRMo8RCsMCNR0Cz;4(
RRRRMRC8CRoMNCs0zCR4Rc;RRRRRRRRR
RRRRRRRRR
R-RR-CRtMNCs0NCRRRd.I8FsRC8CbqR)vCRODHDRVbRNbbsFs0HNCRRRRRRRRRRRRRRR
RRRRUz4RH:RVMR5kOl_C_DDd=.RRR42oCCMsCN0
RRRRR--Q5VRNs88I0H8ERR>(M2RCRC80OFRs0CNCsRIHR0CCLMNDNCRMF8Rkk0b0MRCNCLDRD#CCRO0DHFoOR
RRRRRR4Rzg:NRRRHV58N8s8IH0>ERRRn2oCCMsCN0
RRRRRRRRRRRRRRRRksF0M_C_Rd.<'=R4I'RERCM5N5s8C_so85N8HsI8-0E4FR8IFM0RRn2=kRMlC_ODnD_cN2RM58Rs_N8s5Co6=2RR''j2C2RDR#C';j'
RRRRRRRRRRRRRRRRkIF0M_C_Rd.<'=R4I'RERCM5N5I8C_so85N8HsI8-0E4FR8IFM0RRn2=kRMlC_ODnD_cN2RM58RI_N8s5Co6=2RR''j2C2RDR#C';j'
RRRRRRRRRRRRRRRR0Is__CMd<.R= RWRCIEM5R5I_N8s5CoNs88I0H8ER-48MFI0nFR2RR=M_klODCD_2ncR8NMRN5I8C_so256R'=Rj2'2R#CDCjR''R;
RRRRRCRRMo8RCsMCNR0CzN4g;R
RRRRRR4Rzg:LRRRHV58N8s8IH0=ERRNnRMM8RkOl_C_DDn=cRRRj2oCCMsCN0
RRRRRRRRRRRRRRRRksF0M_C_Rd.<'=R4I'RERCM5N5s8C_so256R'=Rj2'2R#CDCjR''R;
RRRRRRRRRRRRRIRRF_k0CdM_.=R<R''4RCIEM5R5I_N8s5Co6=2RR''j2C2RDR#C';j'
RRRRRRRRRRRRRRRR0Is__CMd<.R= RWRCIEM5R5I_N8s5Co6=2RR''j2C2RDR#C';j'
RRRRRRRR8CMRMoCC0sNC4RzgRL;R-RR-VRQR85N8HsI8R0E<6=R2FRMRHIs0CCRMDNLCsRFR0FkbRk0CLMND#CRCODC0FRDoRHOM8CCCR8
RRRRRzRR.:jRRRHV58N8s8IH0<ER=2R6RMoCC0sNCR
RRRRRRRRRRRRRRFRskC0_M._dRR<=';4'
RRRRRRRRRRRRRRRRkIF0M_C_Rd.<'=R4
';RRRRRRRRRRRRRRRRI_s0CdM_.=R<R;W 
RRRRRRRR8CMRMoCC0sNC.RzjR;
R-RR-CRtMNCs00CRE)CRqOvRCRDDNRM80-sH#00NCR
RRRRRR.Rz4RR:VRFs[MRHRH5I8R0E-2R4RI8FMR0FjCRoMNCs0RC
RRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)Rzq.vdRD:RNDLCRRH#"a17"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloMC5kOl_C_DDnnc*c&2RR""WRH&RMo0CCHs'lCNo5R[2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50EM_klODCD_*ncn+cRR,d.Rb8C02E2R"&RX&"RR0HMCsoC'NHlo[C5+;42
RRRRRRRRRRRRoLCHRM
RRRRRRRRRzRR)dqv.RR:Xv)qd4.X7RR
RRRRRRRRRRRRRbRRFRs0lRNb5=7R>MRH_osC5,[2RRqj=D>RFII_Ns885,j2RRq4=D>RFII_Ns885,42RRq.=D>RFII_Ns885,.2
RRRRRRRRRRRRRRRRRRRRRRRRqRRd>R=RIDF_8IN8ds52q,Rc>R=RIDF_8IN8cs52
,RSSSSSRSR7qu)j>R=RIDF_8sN8js527,Ru4)qRR=>D_FIs8N8s254,uR7)Rq.=D>RFsI_Ns885,.2
SSSSRSSR)7uq=dR>FRDIN_s858sdR2,7qu)c>R=RIDF_8sN8cs52
,RSSSSSRSRW= R>sRI0M_C_,d.RpWBi>R=RiBp,uR7m>R=RksF0k_L#._d5lMk_DOCD._d,,[2Rm1uRR=>I0Fk_#Lk_5d.M_klODCD_,d.R2[2;R
RRRRRRRRRRRRRRFRsks0_C[o52=R<RksF0k_L#._d5lMk_DOCD._d,R[2IMECRF5skC0_M._dR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRIks0_C[o52=R<RkIF0k_L#._d5lMk_DOCD._d,R[2IMECRF5IkC0_M._dR'=R4R'2CCD#R''Z;R
RRRRRRCRRMo8RCsMCNR0Cz;.4
RRRRMRC8CRoMNCs0zCR4RU;RRRRRRRRRR

R-RR-CRtMNCs0NCRRR4nI8FsRC8CbqR)vCRODHDRVbRNbbsFs0HNCRRRRRRRRRRRRRRR
RRRR.z.RH:RVMR5kOl_C_DD4=nRRR42oCCMsCN0
RRRRR--Q5VRNs88I0H8ERR>6M2RCRC80OFRs0CNCsRIHR0CCLMNDNCRMF8Rkk0b0MRCNCLDRD#CCRO0DHFoOR
RRRRRR.Rzd:NRRRHV58N8s8IH0>ERRNnRMM8RkOl_C_DDd=.RRR42oCCMsCN0
RRRRRRRRRRRRRRRRksF0M_C_R4n<'=R4I'RERCM5N5s8C_so85N8HsI8-0E4FR8IFM0RRn2=kRMlC_ODnD_cN2RM58Rs_N8s5Co6=2RR''42MRN8sR5Ns8_Cco52RR='2j'2DRC#'CRj
';RRRRRRRRRRRRRRRRI0Fk__CM4<nR=4R''ERIC5MR58IN_osC58N8s8IH04E-RI8FMR0Fn=2RRlMk_DOCDc_n2MRN8IR5Ns8_C6o52RR='24'R8NMRN5I8C_so25cR'=Rj2'2R#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_Mn_4RR<=WI RERCM5N5I8C_so85N8HsI8-0E4FR8IFM0RRn2=kRMlC_ODnD_cN2RM58RI_N8s5Co6=2RR''42MRN8IR5Ns8_Cco52RR='2j'2DRC#'CRj
';RRRRRRRRCRM8oCCMsCN0Rdz.NR;
RRRRRzRR.RdL:VRHR85N8HsI8R0E>RRnNRM8M_klODCD_Rd./4=R2CRoMNCs0RC
RRRRRRRRRRRRRsRRF_k0C4M_n=R<R''4RCIEM5R5s_N8s5CoNs88I0H8ER-48MFI0nFR2RR=M_klODCD_2ncR8NMRN5s8C_so256R'=RjR'2NRM858sN_osC5Rc2=jR''R22CCD#R''j;R
RRRRRRRRRRRRRRFRIkC0_Mn_4RR<='R4'IMECRI55Ns8_CNo58I8sHE80-84RF0IMF2RnRM=RkOl_C_DDnRc2NRM858IN_osC5R62=jR''N2RM58RI_N8s5Coc=2RR''j2C2RDR#C';j'
RRRRRRRRRRRRRRRR0Is__CM4<nR= RWRCIEM5R5I_N8s5CoNs88I0H8ER-48MFI0nFR2RR=M_klODCD_2ncR8NMRN5I8C_so256R'=RjR'2NRM858IN_osC5Rc2=jR''R22CCD#R''j;R
RRRRRRMRC8CRoMNCs0zCR.;dL
RRRRRRRRdz.ORR:H5VRNs88I0H8ERR=nMRN8kRMlC_ODdD_.RR=4o2RCsMCN
0CRRRRRRRRRRRRRRRRs0Fk__CM4<nR=4R''ERIC5MR58sN_osC5R62=4R''N2RM58Rs_N8s5Coc=2RR''j2C2RDR#C';j'
RRRRRRRRRRRRRRRRkIF0M_C_R4n<'=R4I'RERCM5N5I8C_so256R'=R4R'2NRM858IN_osC5Rc2=jR''R22CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C_R4n<W=R ERIC5MR58IN_osC5R62=4R''N2RM58RI_N8s5Coc=2RR''j2C2RDR#C';j'
RRRRRRRR8CMRMoCC0sNC.Rzd
O;RRRRRRRRzL.dRH:RVNR58I8sHE80R6=RR8NMRlMk_DOCD._dRR/=4o2RCsMCN
0CRRRRRRRRRRRRRRRRs0Fk__CM4<nR=4R''ERIC5MR58sN_osC58N8s8IH04E-RI8FMR0Fn=2RRlMk_DOCD._d2C2RDR#C';j'
RRRRRRRRRRRRRRRRkIF0M_C_R4n<'=R4I'RERCM5N5I8C_so85N8HsI8-0E4FR8IFM0RRn2=kRMlC_ODdD_.R22CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C_R4n<W=R ERIC5MR58IN_osC58N8s8IH04E-RI8FMR0Fn=2RRlMk_DOCD._d2C2RDR#C';j'
RRRRRRRR8CMRMoCC0sNC.RzdRL;R-RR-VRQR85N8HsI8R0E<6=R2FRMRHIs0CCRMDNLCsRFR0FkbRk0CLMND#CRCODC0FRDoRHOM8CCCR8
RRRRRzRR.:cRRRHV58N8s8IH0<ER=2RcRMoCC0sNCR
RRRRRRRRRRRRRRFRskC0_Mn_4RR<=';4'
RRRRRRRRRRRRRRRRkIF0M_C_R4n<'=R4
';RRRRRRRRRRRRRRRRI_s0C4M_n=R<R;W 
RRRRRRRR8CMRMoCC0sNC.RzcR;
R-RR-CRtMNCs00CRE)CRqOvRCRDDNRM80-sH#00NCR
RRRRRR.Rz6RR:VRFs[MRHRH5I8R0E-2R4RI8FMR0FjCRoMNCs0RC
RRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)Rzqnv4RD:RNDLCRRH#"a17"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloMC5kOl_C_DDnnc*cRR+M_klODCD_*d.dR.2&WR""RR&HCM0o'CsHolNC25[R"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05lMk_DOCDc_n*Rnc+kRMlC_ODdD_..*dR4+Rn8,RCEb02&2RR""XRH&RMo0CCHs'lCNo54[+2R;
RRRRRRRRRLRRCMoH
RRRRRRRRRRRRqz)vR4n:qR)vX4n4
7RRRRRRRRRRRRRRRRRb0FsRblNRR57=H>RMC_so25[,jRqRR=>D_FII8N8s25j,4RqRR=>D_FII8N8s254,.RqRR=>D_FII8N8s25.,R
RRRRRRRRRRRRRRRRRRRRRRRRRq=dR>FRDIN_I858sdR2,7qu)j>R=RIDF_8sN8js527,Ru4)qRR=>D_FIs8N8s254,uR7)Rq.=D>RFsI_Ns885,.2
SSSSRSSR)7uq=dR>FRDIN_s858sdR2,W= R>sRI0M_C_,4nRpWBi>R=RiBp,uR7m>R=RksF0k_L#n_45lMk_DOCDn_4,,[2Rm1uRR=>I0Fk_#Lk_54nM_klODCD_,4nR2[2;R
RRRRRRRRRRRRRRFRsks0_C[o52=R<RksF0k_L#n_45lMk_DOCDn_4,R[2IMECRF5skC0_Mn_4R'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRIks0_C[o52=R<RkIF0k_L#n_45lMk_DOCDn_4,R[2IMECRF5IkC0_Mn_4R'=R4R'2CCD#R''Z;R
RRRRRRMRC8CRoMNCs0zCR.
6;RRRRCRM8oCCMsCN0R.z.;R
RRRRRRR
RRRRRRRRRRRRRRRRRRRRRRRRRRM
C8sRNO0EHCkO0sLCRD	FO_lsN;-

-FRM__sIOOEC	sRNONE
sHOE00COkRsCMsF_IE_OCRO	F)VRq)v_WR_)HN#
0H0sLCk0RMoCC0sNFss_CsbF0RR:#H0sM
o;Ns00H0LkCCRoMNCs0_FssFCbsF0RVFRM__sIOOEC	RR:NEsOHO0C0CksRRH#"N7kDFRbsA0RD	FORv)qR0MFRb#kb0FsC$8RCR0,HCMVsMsHoCR1D0CORv)q"O;
FFlbM0CMRqX)vXd.4R7RRsbF0
R5RRRRRRRR7RumRRR:FRk0#_08koDFHRO;RRRRR
RRRRRRRRRR1RumRRR:FRk0#_08koDFH
O;
RRRRRRRRRqjR:RRRRHM#_08koDFH
O;RRRRRRRRqR4RRRR:H#MR0k8_DHFoOR;
RRRRRqRR.RRRRH:RM0R#8D_kFOoH;R
RRRRRRdRqRRRR:MRHR8#0_FkDo;HO
RRRRRRRRRqcR:RRRRHM#_08koDFH
O;RRRRRRRR7RRRRRR:H#MR0k8_DHFoOR;
RRRRR7RRuj)qRH:RM0R#8D_kFOoH;R
RRRRRRuR7)Rq4:MRHR8#0_FkDo;HO
RRRRRRRR)7uq:.RRRHM#_08koDFH
O;RRRRRRRR7qu)dRR:H#MR0k8_DHFoOR;
RRRRR7RRuc)qRH:RM0R#8D_kFOoH;R
RRRRRRBRWpRiR:MRHR8#0_FkDo;HORRRRRRRR
RRRRRRRRRW R:RRRRHM#_08koDFHRO
RRRRR;R2RCR
MO8RFFlbM0CM;F
OlMbFCRM0Xv)qn4cX7RRRb0FsRR5
RRRRR7RRuRmRRF:Rk#0R0k8_DHFoOR;RRRRRRRR
RRRRR1RRuRmRRF:Rk#0R0k8_DHFoO
;
RRRRRRRRqRjRRRR:H#MR0k8_DHFoOR;
RRRRRqRR4RRRRH:RM0R#8D_kFOoH;R
RRRRRR.RqRRRR:MRHR8#0_FkDo;HO
RRRRRRRRRqdR:RRRRHM#_08koDFH
O;RRRRRRRRqRcRRRR:H#MR0k8_DHFoOR;
RRRRRqRR6RRRRH:RM0R#8D_kFOoH;R
RRRRRRRR7RRRR:MRHR8#0_FkDo;HO
RRRRRRRR)7uq:jRRRHM#_08koDFH
O;RRRRRRRR7qu)4RR:H#MR0k8_DHFoOR;
RRRRR7RRu.)qRH:RM0R#8D_kFOoH;R
RRRRRRuR7)Rqd:MRHR8#0_FkDo;HO
RRRRRRRR)7uq:cRRRHM#_08koDFH
O;RRRRRRRR7qu)6RR:H#MR0k8_DHFoOR;
RRRRRWRRBRpiRH:RM0R#8D_kFOoH;RRRRRRRRR
RRRRRR RWRRRR:MRHR8#0_FkDo
HORRRRR2RR;
RRCRM8ObFlFMMC0V;
k0MOHRFMo_C0M_kln8c5CEb0:MRH0CCoss2RCs0kMMRH0CCos#RH
sPNHDNLCNRPDRR:HCM0oRCs:j=R;C
Lo
HMRNRPD=R:Rb8C0nE/cR;
RRHV5C58bR0ElRF8nRc2>URc2ER0CRM
RPRRN:DR=NRPDRR+4R;
R8CMR;HV
sRRCs0kMNRPDC;
Mo8RCM0_knl_cV;
k0MOHRFMo_C0D0CVFsPC_5d.80CbERR:HCM0o2CsR0sCkRsMHCM0oRCsHL#
CMoH
sRRCs0kMC58bR0ElRF8n;c2
8CMR0oC_VDC0CFPs._d;k
VMHO0FoMRCD0_CFV0P5Cs80CbERR:HCM0o;CsRGlNRH:RMo0CCRs2skC0sHMRMo0CCHsR#N
PsLHNDPCRN:DRR0HMCsoCRR:=jL;
CMoH
HRRV8R5CEb0Rl-RN>GR=2RjRC0EMR
RRNRPD=R:Rb8C0-ERRGlN;R
RCCD#
RRRRDPNRR:=80CbER;
R8CMR;HV
sRRCs0kMN5PD
2;CRM8o_C0D0CVFsPC;k
VMHO0FoMRCM0_kdl_.C58bR0E:MRH0CCoss2RCs0kMMRH0CCos#RH
sPNHDNLCNRPDRR:HCM0oRCs:j=R;C
Lo
HMRVRHRC58bR0E<c=RUMRN8CR8bR0E>nR42ER0CRM
RRRRPRND:4=R;R
RCRM8H
V;RCRs0MksRDPN;M
C8CRo0k_Ml._d;k
VMHO0FoMRCM0_k4l_nC58bR0E:MRH0CCoss2RCs0kMMRH0CCos#RH
sPNHDNLCNRPDRR:HCM0oRCs:j=R;C
Lo
HMRVRHRC58bR0E<4=RnMRN8CR8bR0E>2RjRC0EMR
RRPRRN:DR=;R4
CRRMH8RVR;
R0sCkRsMP;ND
8CMR0oC_lMk_;4n
MVkOF0HMCRo0M_C8C_8b50E#CHxRH:RMo0CC;sRRb8C0:ERR0HMCsoC2CRs0MksR0HMCsoCR
H#PHNsNCLDRMlH_x#HCRR:HCM0oRCs:j=R;C
Lo
HMRHRlMH_#x:CR=CR8b;0E
HRRV#R5HRxC<CR8b20ERC0EMR
RRHRlMH_#x:CR=HR#x
C;RMRC8VRH;R
RskC0slMRH#M_H;xC
8CMR0oC_8CM_b8C0
E;O#FM00NMRlMk_DOCDc_nRH:RMo0CC:sR=CRo0k_Mlc_n5b8C0;E2
MOF#M0N0CRDVP0FCds_.RR:HCM0oRCs:o=RCD0_CFV0P_Csd8.5CEb02O;
F0M#NRM0M_klODCD_Rd.:MRH0CCos=R:R0oC_lMk_5d.D0CVFsPC_2d.;F
OMN#0MD0RCFV0P_Cs4:nRR0HMCsoCRR:=o_C0D0CVFsPC5VDC0CFPs._d,.Rd2O;
F0M#NRM0M_klODCD_R4n:MRH0CCos=R:R0oC_lMk_54nD0CVFsPC_24n;0

$RbCF_k0L_k#0C$b_RncHN#Rs$sNRk5MlC_ODnD_cFR8IFM0RRj,I0H8ER-48MFI0jFR2VRFR8#0_oDFH
O;0C$bR0Fk_#Lk_b0$C._dRRH#NNss$MR5kOl_C_DDd8.RF0IMF,RjR8IH04E-RI8FMR0FjF2RV0R#8F_Do;HO
b0$CkRF0k_L#$_0b4C_n#RHRsNsN5$RM_klODCD_R4n8MFI0jFR,HRI8-0E4FR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNRksF0k_L#c_nRF:RkL0_k0#_$_bCnRc;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RVFR8k50RHkMb0FR0RH0s-N#002C#
o#HMRNDs0Fk_#Lk_Rd.:kRF0k_L#$_0bdC_.R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFRk8F0HR5M0bkRR0F0-sH#00NC
#2#MHoNsDRF_k0L_k#4:nRR0Fk_#Lk_b0$Cn_4;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFV80FkRM5HbRk000FRs#H-0CN0##2
HNoMDFRskC0_MRR:#_08DHFoOC_POs0F5lMk_DOCDc_nRI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-C-RMDNLCV#RF0sRs#H-0CN0#H
#oDMNRkIF0k_L#c_nRF:RkL0_k0#_$_bCnRc;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RVFR8k50RHkMb0FR0RH0s-N#002C#
o#HMRNDI0Fk_#Lk_Rd.:kRF0k_L#$_0bdC_.R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFRk8F0HR5M0bkRR0F0-sH#00NC
#2#MHoNIDRF_k0L_k#4:nRR0Fk_#Lk_b0$Cn_4;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFV80FkRM5HbRk000FRs#H-0CN0##2
HNoMDFRIkC0_MRR:#_08DHFoOC_POs0F5lMk_DOCDc_nRI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-C-RMDNLCV#RF0sRs#H-0CN0#H
#oDMNRksF0M_C_Rd.:0R#8F_Do;HO
o#HMRNDs0Fk__CM4:nRR8#0_oDFH
O;#MHoNIDRF_k0CdM_.RR:#_08DHFoO#;
HNoMDFRIkC0_Mn_4R#:R0D8_FOoH;H
#oDMNR0Is_RCM:0R#8F_Do_HOP0COFMs5kOl_C_DDn8cRF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RHIs0CCRMDNLCV#RFCsRNROEsRFIF)VRqOvRC#DD
o#HMRNDI_s0CdM_.RR:#_08DHFoO#;
HNoMDsRI0M_C_R4n:0R#8F_Do;HO
o#HMRNDHsM_C:oRR8#0_oDFHPO_CFO0sH5I8-0E4FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-#RkC08RFCRso0H#C7sRQ
hR#MHoNsDRF_k0sRCo:0R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-#RkC08RFCRso0H#C7sRm
za#MHoNIDRF_k0sRCo:0R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-#RkC08RFCRso0H#C7sRm
za#MHoNsDRNs8_C:oRR8#0_oDFHPO_CFO0s85N8HsI8-0E4FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-#RkC08RFCRso0H#CqsR7
7)#MHoNIDRNs8_C:oRR8#0_oDFHPO_CFO0s85N8HsI8-0E4FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-#RkC08RFCRso0H#CqsR7
7)#MHoNDDRFsI_Ns88R#:R0D8_FOoH_OPC05Fs6FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-8RN8LsRHR0#HkMb0FR0Rv)qRDOCD5#RcHRL0s#RCHJks2C8
o#HMRNDD_FII8N8sRR:#_08DHFoOC_POs0F586RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-N-R8R8sL#H0RbHMk00RFqR)vCRODRD#5LcRHR0#skCJH8sC20
N0LsHkR0C\N3slV_FV0#C\RR:#H0sM
o;
oLCH
M
RRRR-Q-RV8RN8HsI8R0E<RR6NH##o'MRj0'RFMRkk8#CR0LH#R
RRjRzRRR:H5VRNs88I0H8ERR=4o2RCsMCN
0CRRRRRRRRD_FIs8N8s=R<Rj"jj"jjRs&RNs8_Cjo52R;
RRRRRDRRFII_Ns88RR<="jjjjRj"&NRI8C_so25j;R
RRMRC8CRoMNCs0zCRjR;
RzRR4:RRRRHV58N8s8IH0=ERRR.2oCCMsCN0
RRRRRRRRIDF_8sN8<sR=jR"j"jjRs&RNs8_C4o5RI8FMR0Fj
2;RRRRRRRRD_FII8N8s=R<Rj"jjRj"&NRI8C_soR548MFI0jFR2R;
RCRRMo8RCsMCNR0Cz
4;RRRRzR.R:VRHR85N8HsI8R0E=2RdRMoCC0sNCR
RRRRRRFRDIN_s8R8s<"=Rj"jjRs&RNs8_C.o5RI8FMR0Fj
2;RRRRRRRRD_FII8N8s=R<Rj"jj&"RR8IN_osC58.RF0IMF2Rj;R
RRMRC8CRoMNCs0zCR.R;
RzRRd:RRRRHV58N8s8IH0=ERRRc2oCCMsCN0
RRRRRRRRIDF_8sN8<sR=jR"j&"RR8sN_osC58dRF0IMF2Rj;R
RRRRRRFRDIN_I8R8s<"=RjRj"&NRI8C_soR5d8MFI0jFR2R;
RCRRMo8RCsMCNR0Cz
d;SSzc:VRHR85N8HsI8R0E=2R6RMoCC0sNCS
SD_FIs8N8s=R<R''jRs&RNs8_Cco5RI8FMR0Fj
2;SFSDIN_I8R8s<'=Rj&'RR8IN_osC58cRF0IMF2Rj;C
SMo8RCsMCNR0Cz
c;RRRRzR6R:VRHR85N8HsI8R0E>2R6RMoCC0sNCR
RRRRRRFRDIN_s8R8s<s=RNs8_C6o5RI8FMR0Fj
2;RRRRRRRRD_FII8N8s=R<R8IN_osC586RF0IMF2Rj;R
RRMRC8CRoMNCs0zCR6
;
RRRR-Q-RV8R5HsM_CRo2sHCo#s0CRh7QRHk#MBoRpRi
RzRRn:RRRRHV5M8H_osC2CRoMNCs0RC
RRRRRbRRsCFO#5#RB,piRh7Q2CRLo
HMRRRRRRRRRRRRH5VRBRpi=4R''MRN8pRBiP'CC2M0RC0EMR
RRRRRRRRRRRRRRMRH_osCRR<=7;Qh
RRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMRFbsO#C#;R
RRMRC8CRoMNCs0zCRnR;
RzRR(:RRRRHV50MFRM8H_osC2CRoMNCs0RC
RRRRRRRRRHRRMC_so=R<Rh7Q;R
RRMRC8CRoMNCs0zCR(
;
RRRR-Q-RV8R5F_k0s2CoRosCHC#0smR7zkaR#oHMRpmBiR
RRURzs:RRRRHV5Fs8ks0_CRo2oCCMsCN0
RRRRRRRRFbsO#C#R_5)miBp,FRsks0_CRo2LHCoMR
RRRRRRRRRRVRHR_5)miBpR'=R4N'RM)8R_pmBiP'CC2M0RC0EMR
RRRRRRRRRRRRRR_R)7amzRR<=s0Fk_osC;R
RRRRRRRRRRMRC8VRH;R
RRRRRRMRC8sRbF#OC#R;
RCRRMo8RCsMCNR0Cz;Us
RRRRszgRRR:H5VRMRF0sk8F0C_soo2RCsMCN
0CRRRRRRRRRRRR)m_7z<aR=FRsks0_C
o;RRRRCRM8oCCMsCN0Rszg;R

R-RR-VRQRF58ks0_CRo2sHCo#s0CRz7ma#RkHRMomiBp
RRRRIzURRR:H5VRIk8F0C_soo2RCsMCN
0CRRRRRRRRbOsFCR##5mW_B,piRkIF0C_soL2RCMoH
RRRRRRRRRRRRRHV5mW_BRpi=4R''MRN8_RWmiBp'CCPMR020MEC
RRRRRRRRRRRRRRRR7W_mRza<I=RF_k0s;Co
RRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMRFbsO#C#;R
RRMRC8CRoMNCs0zCRU
I;RRRRzRgIRH:RVMR5FI0R80Fk_osC2CRoMNCs0RC
RRRRRRRRRWRR_z7ma=R<RkIF0C_soR;
RCRRMo8RCsMCNR0Cz;gI
R
RR-R-RRQV58N8sC_sos2RC#oH0RCsq)77RHk#MBoRpRi
RzRR4RjR:VRHRN5s8_8ss2CoRMoCC0sNCR
RRRRRRsRbF#OC#)R5_pmBi),Rq)772CRLo
HMRRRRRRRRRRRRH5VR)B_mp=iRR''4R8NMRm)_B'piCMPC002RE
CMRRRRRRRRRRRRRRRRs_N8sRCo<)=Rq)7758N8s8IH04E-RI8FMR0Fj
2;RRRRRRRRRRRRCRM8H
V;RRRRRRRRCRM8bOsFC;##
RRRR8CMRMoCC0sNC4RzjR;
RzRR4:4RRRHV50MFR8sN8ss_CRo2oCCMsCN0
RRRRRRRRRRRR8sN_osCRR<=)7q7)R;
RCRRMo8RCsMCNR0Cz;44
R
RR-R-RRQV58N8sC_sos2RC#oH0RCsq)77RHk#MBoRpRi
RzRR4R.R:VRHRN5I8_8ss2CoRMoCC0sNCR
RRRRRRsRbF#OC#BR5pRi,W7q7)L2RCMoH
RRRRRRRRRRRRRHV5iBpR'=R4N'RMB8RpCi'P0CM2ER0CRM
RRRRRRRRRRRRRIRRNs8_C<oR=qRW757)Ns88I0H8ER-48MFI0jFR2R;
RRRRRRRRRCRRMH8RVR;
RRRRRCRRMb8RsCFO#
#;RRRRCRM8oCCMsCN0R.z4;R
RR4RzdRR:H5VRMRF0I8N8sC_soo2RCsMCN
0CRRRRRRRRRRRRI_N8sRCo<W=Rq)77;R
RRMRC8CRoMNCs0zCR4
d;RRRRRRRR
RRRRR--tCCMsCN0RC0ERv)qRDOCDN#RM#8RCODC0FRDo
HORRRRzR4c:FRVsRRHH5MRM_klODCD_Rnc-2R4RI8FMR0FjCRoMNCs0RC
R-RR-VRQR85N8HsI8R0E>2R6RCMC8FR0RCOsNR0CI0sHCMRCNCLDR8NMR0FkbRk0CLMND#CRCODC0FRDo
HORRRRRRRRzR46:VRHR85N8HsI8R0E>2RnRMoCC0sNCR
RRRRRRRRRRRRRRFRskC0_M25HRR<='R4'IMECRN5s8C_so85N8HsI8-0E4FR8IFM0RRn2=2RHR#CDCjR''R;
RRRRRRRRRRRRRIRRF_k0CHM52=R<R''4RCIEMIR5Ns8_CNo58I8sHE80-84RF0IMF2RnRH=R2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0CHM52=R<RRW IMECRN5I8C_so85N8HsI8-0E4FR8IFM0RRn2=2RHR#CDCjR''R;
RRRRRCRRMo8RCsMCNR0Cz;46
RRRRR--Q5VRNs88I0H8E=R<RR62MIFRsCH0RNCMLRDCFFsRkk0b0MRCNCLDRD#CCRO0DHFoOCRMC88C
RRRRRRRRnz4RH:RVNR58I8sHE80RR<=no2RCsMCN
0CRRRRRRRRRRRRRRRRs0Fk_5CMH<2R=4R''R;
RRRRRRRRRRRRRIRRF_k0CHM52=R<R''4;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R R;
RRRRRCRRMo8RCsMCNR0Cz;4n
RRRRR--tCCMsCN0RC0ERv)qRDOCDN#RM08Rs#H-0CN0#R
RRRRRR4Rz(RR:VRFs[MRHRH5I8R0E-2R4RI8FMR0FjCRoMNCs0RC
RRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)RzqcvnRD:RNDLCRRH#"a17"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloHC5*2ncR"&RW&"RR0HMCsoC'NHlo[C52RR&"R "&MRH0CCosl'HN5oCo_C0C_M880CbEH55+*42nRc,80CbER22&XR""RR&HCM0o'CsHolNC+5[4
2;RRRRRRRRRRRRLHCoMR
RRRRRRRRRR)RzqcvnRX:R)nqvc7X4RR
RRRRRRRRRRRRRRFRbsl0RN5bR7>R=R_HMs5Co[R2,q=jR>FRDIN_I858sjR2,q=4R>FRDIN_I858s4R2,q=.R>FRDIN_I858s.
2,RRRRRRRRRRRRRRRRRRRRRRRRRdRqRR=>D_FII8N8s25d,cRqRR=>D_FII8N8s25c,6RqRR=>D_FII8N8s256,SR
SSSSS7RRuj)qRR=>D_FIs8N8s25j,uR7)Rq4=D>RFsI_Ns885,42R)7uq=.R>FRDIN_s858s.
2,SSSSSRSR7qu)d>R=RIDF_8sN8ds527,Ruc)qRR=>D_FIs8N8s25c,uR7)Rq6=D>RFsI_Ns885,62RS
SSSSSR RWRR=>I_s0CHM52W,RBRpi=B>RpRi,7Rum=s>RF_k0L_k#nHc5,,[2Rm1uRR=>I0Fk_#Lk_5ncH2,[2R;
RRRRRRRRRRRRRsRRF_k0s5Co[<2R=FRskL0_kn#_c,5H[I2RERCM5ksF0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRkIF0C_so25[RR<=I0Fk_#Lk_5ncH2,[RCIEMIR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRCRRMo8RCsMCNR0Cz;4(
RRRRMRC8CRoMNCs0zCR4Rc;RRRRRRRRR
RRRRRRRRR
R-RR-CRtMNCs0NCRRRd.I8FsRC8CbqR)vCRODHDRVbRNbbsFs0HNCRRRRRRRRRRRRRRR
RRRRUz4RH:RVMR5kOl_C_DDd=.RRR42oCCMsCN0
RRRRR--Q5VRNs88I0H8ERR>(M2RCRC80OFRs0CNCsRIHR0CCLMNDNCRMF8Rkk0b0MRCNCLDRD#CCRO0DHFoOR
RRRRRR4Rzg:NRRRHV58N8s8IH0>ERRRn2oCCMsCN0
RRRRRRRRRRRRRRRRksF0M_C_Rd.<'=R4I'RERCM5N5s8C_so85N8HsI8-0E4FR8IFM0RRn2=kRMlC_ODnD_cN2RM58Rs_N8s5Co6=2RR''j2C2RDR#C';j'
RRRRRRRRRRRRRRRRkIF0M_C_Rd.<'=R4I'RERCM5N5I8C_so85N8HsI8-0E4FR8IFM0RRn2=kRMlC_ODnD_cN2RM58RI_N8s5Co6=2RR''j2C2RDR#C';j'
RRRRRRRRRRRRRRRR0Is__CMd<.R= RWRCIEM5R5I_N8s5CoNs88I0H8ER-48MFI0nFR2RR=M_klODCD_2ncR8NMRN5I8C_so256R'=Rj2'2R#CDCjR''R;
RRRRRCRRMo8RCsMCNR0CzN4g;R
RRRRRR4Rzg:LRRRHV58N8s8IH0=ERRNnRMM8RkOl_C_DDn=cRRRj2oCCMsCN0
RRRRRRRRRRRRRRRRksF0M_C_Rd.<'=R4I'RERCM5N5s8C_so256R'=Rj2'2R#CDCjR''R;
RRRRRRRRRRRRRIRRF_k0CdM_.=R<R''4RCIEM5R5I_N8s5Co6=2RR''j2C2RDR#C';j'
RRRRRRRRRRRRRRRR0Is__CMd<.R= RWRCIEM5R5I_N8s5Co6=2RR''j2C2RDR#C';j'
RRRRRRRR8CMRMoCC0sNC4RzgRL;R-RR-VRQR85N8HsI8R0E<6=R2FRMRHIs0CCRMDNLCsRFR0FkbRk0CLMND#CRCODC0FRDoRHOM8CCCR8
RRRRRzRR.:jRRRHV58N8s8IH0<ER=2R6RMoCC0sNCR
RRRRRRRRRRRRRRFRskC0_M._dRR<=';4'
RRRRRRRRRRRRRRRRkIF0M_C_Rd.<'=R4
';RRRRRRRRRRRRRRRRI_s0CdM_.=R<R;W 
RRRRRRRR8CMRMoCC0sNC.RzjR;
R-RR-CRtMNCs00CRE)CRqOvRCRDDNRM80-sH#00NCR
RRRRRR.Rz4RR:VRFs[MRHRH5I8R0E-2R4RI8FMR0FjCRoMNCs0RC
RRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)Rzq.vdRD:RNDLCRRH#"a17"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloMC5kOl_C_DDnnc*c&2RR""WRH&RMo0CCHs'lCNo5R[2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50EM_klODCD_*ncn+cRR,d.Rb8C02E2R"&RX&"RR0HMCsoC'NHlo[C5+;42
RRRRRRRRRRRRoLCHRM
RRRRRRRRRzRR)dqv.RR:Xv)qd4.X7RR
RRRRRRRRRRRRRbRRFRs0lRNb5=7R>MRH_osC5,[2RRqj=D>RFII_Ns885,j2RRq4=D>RFII_Ns885,42RRq.=D>RFII_Ns885,.2
RRRRRRRRRRRRRRRRRRRRRRRRqRRd>R=RIDF_8IN8ds52q,Rc>R=RIDF_8IN8cs52
,RSSSSSRSR7qu)j>R=RIDF_8sN8js527,Ru4)qRR=>D_FIs8N8s254,uR7)Rq.=D>RFsI_Ns885,.2
SSSSRSSR)7uq=dR>FRDIN_s858sdR2,7qu)c>R=RIDF_8sN8cs52
,RSSSSSRSRW= R>sRI0M_C_,d.RpWBi>R=RiBp,uR7m>R=RksF0k_L#._d5lMk_DOCD._d,,[2Rm1uRR=>I0Fk_#Lk_5d.M_klODCD_,d.R2[2;R
RRRRRRRRRRRRRRFRsks0_C[o52=R<RksF0k_L#._d5lMk_DOCD._d,R[2IMECRF5skC0_M._dR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRIks0_C[o52=R<RkIF0k_L#._d5lMk_DOCD._d,R[2IMECRF5IkC0_M._dR'=R4R'2CCD#R''Z;R
RRRRRRCRRMo8RCsMCNR0Cz;.4
RRRRMRC8CRoMNCs0zCR4RU;RRRRRRRRRR

R-RR-CRtMNCs0NCRRR4nI8FsRC8CbqR)vCRODHDRVbRNbbsFs0HNCRRRRRRRRRRRRRRR
RRRR.z.RH:RVMR5kOl_C_DD4=nRRR42oCCMsCN0
RRRRR--Q5VRNs88I0H8ERR>6M2RCRC80OFRs0CNCsRIHR0CCLMNDNCRMF8Rkk0b0MRCNCLDRD#CCRO0DHFoOR
RRRRRR.Rzd:NRRRHV58N8s8IH0>ERRNnRMM8RkOl_C_DDd=.RRR42oCCMsCN0
RRRRRRRRRRRRRRRRksF0M_C_R4n<'=R4I'RERCM5N5s8C_so85N8HsI8-0E4FR8IFM0RRn2=kRMlC_ODnD_cN2RM58Rs_N8s5Co6=2RR''42MRN8sR5Ns8_Cco52RR='2j'2DRC#'CRj
';RRRRRRRRRRRRRRRRI0Fk__CM4<nR=4R''ERIC5MR58IN_osC58N8s8IH04E-RI8FMR0Fn=2RRlMk_DOCDc_n2MRN8IR5Ns8_C6o52RR='24'R8NMRN5I8C_so25cR'=Rj2'2R#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_Mn_4RR<=WI RERCM5N5I8C_so85N8HsI8-0E4FR8IFM0RRn2=kRMlC_ODnD_cN2RM58RI_N8s5Co6=2RR''42MRN8IR5Ns8_Cco52RR='2j'2DRC#'CRj
';RRRRRRRRCRM8oCCMsCN0Rdz.NR;
RRRRRzRR.RdL:VRHR85N8HsI8R0E>RRnNRM8M_klODCD_Rd./4=R2CRoMNCs0RC
RRRRRRRRRRRRRsRRF_k0C4M_n=R<R''4RCIEM5R5s_N8s5CoNs88I0H8ER-48MFI0nFR2RR=M_klODCD_2ncR8NMRN5s8C_so256R'=RjR'2NRM858sN_osC5Rc2=jR''R22CCD#R''j;R
RRRRRRRRRRRRRRFRIkC0_Mn_4RR<='R4'IMECRI55Ns8_CNo58I8sHE80-84RF0IMF2RnRM=RkOl_C_DDnRc2NRM858IN_osC5R62=jR''N2RM58RI_N8s5Coc=2RR''j2C2RDR#C';j'
RRRRRRRRRRRRRRRR0Is__CM4<nR= RWRCIEM5R5I_N8s5CoNs88I0H8ER-48MFI0nFR2RR=M_klODCD_2ncR8NMRN5I8C_so256R'=RjR'2NRM858IN_osC5Rc2=jR''R22CCD#R''j;R
RRRRRRMRC8CRoMNCs0zCR.;dL
RRRRRRRRdz.ORR:H5VRNs88I0H8ERR=nMRN8kRMlC_ODdD_.RR=4o2RCsMCN
0CRRRRRRRRRRRRRRRRs0Fk__CM4<nR=4R''ERIC5MR58sN_osC5R62=4R''N2RM58Rs_N8s5Coc=2RR''j2C2RDR#C';j'
RRRRRRRRRRRRRRRRkIF0M_C_R4n<'=R4I'RERCM5N5I8C_so256R'=R4R'2NRM858IN_osC5Rc2=jR''R22CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C_R4n<W=R ERIC5MR58IN_osC5R62=4R''N2RM58RI_N8s5Coc=2RR''j2C2RDR#C';j'
RRRRRRRR8CMRMoCC0sNC.Rzd
O;RRRRRRRRzL.dRH:RVNR58I8sHE80R6=RR8NMRlMk_DOCD._dRR/=4o2RCsMCN
0CRRRRRRRRRRRRRRRRs0Fk__CM4<nR=4R''ERIC5MR58sN_osC58N8s8IH04E-RI8FMR0Fn=2RRlMk_DOCD._d2C2RDR#C';j'
RRRRRRRRRRRRRRRRkIF0M_C_R4n<'=R4I'RERCM5N5I8C_so85N8HsI8-0E4FR8IFM0RRn2=kRMlC_ODdD_.R22CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C_R4n<W=R ERIC5MR58IN_osC58N8s8IH04E-RI8FMR0Fn=2RRlMk_DOCD._d2C2RDR#C';j'
RRRRRRRR8CMRMoCC0sNC.RzdRL;R-RR-VRQR85N8HsI8R0E<6=R2FRMRHIs0CCRMDNLCsRFR0FkbRk0CLMND#CRCODC0FRDoRHOM8CCCR8
RRRRRzRR.:cRRRHV58N8s8IH0<ER=2RcRMoCC0sNCR
RRRRRRRRRRRRRRFRskC0_Mn_4RR<=';4'
RRRRRRRRRRRRRRRRkIF0M_C_R4n<'=R4
';RRRRRRRRRRRRRRRRI_s0C4M_n=R<R;W 
RRRRRRRR8CMRMoCC0sNC.RzcR;
R-RR-CRtMNCs00CRE)CRqOvRCRDDNRM80-sH#00NCR
RRRRRR.Rz6RR:VRFs[MRHRH5I8R0E-2R4RI8FMR0FjCRoMNCs0RC
RRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)Rzqnv4RD:RNDLCRRH#"a17"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloMC5kOl_C_DDnnc*cRR+M_klODCD_*d.dR.2&WR""RR&HCM0o'CsHolNC25[R"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05lMk_DOCDc_n*Rnc+kRMlC_ODdD_..*dR4+Rn8,RCEb02&2RR""XRH&RMo0CCHs'lCNo54[+2R;
RRRRRRRRRLRRCMoH
RRRRRRRRRRRRqz)vR4n:qR)vX4n4
7RRRRRRRRRRRRRRRRRb0FsRblNRR57=H>RMC_so25[,jRqRR=>D_FII8N8s25j,4RqRR=>D_FII8N8s254,.RqRR=>D_FII8N8s25.,R
RRRRRRRRRRRRRRRRRRRRRRRRRq=dR>FRDIN_I858sdR2,7qu)j>R=RIDF_8sN8js527,Ru4)qRR=>D_FIs8N8s254,uR7)Rq.=D>RFsI_Ns885,.2
SSSSRSSR)7uq=dR>FRDIN_s858sdR2,W= R>sRI0M_C_,4nRpWBi>R=RiBp,uR7m>R=RksF0k_L#n_45lMk_DOCDn_4,,[2Rm1uRR=>I0Fk_#Lk_54nM_klODCD_,4nR2[2;R
RRRRRRRRRRRRRRFRsks0_C[o52=R<RksF0k_L#n_45lMk_DOCDn_4,R[2IMECRF5skC0_Mn_4R'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRFRIks0_C[o52=R<RkIF0k_L#n_45lMk_DOCDn_4,R[2IMECRF5IkC0_Mn_4R'=R4R'2CCD#R''Z;R
RRRRRRMRC8CRoMNCs0zCR.
6;RRRRCRM8oCCMsCN0R.z.;R
RRRRRRR
RRRRRRRRRRRRRRRRRRRRRRRRRRM
C8sRNO0EHCkO0sMCRFI_s_COEO
	;RRRRRRRRRRRRRRRRRRRRRRRRR
RR---
--
-R#pN0lRHblDCCNM00MHFRRH#8NCVk
D0-N-
sHOE00COkRsC#CCDOs0_NFlRVqR)vW_)_H)R#k
VMHO0FoMRCC0_M88_CEb05x#HCRR:HCM0oRCs;CR8bR0E:MRH0CCoss2RCs0kMMRH0CCos#RH
sPNHDNLCHRlMH_#x:CRR0HMCsoCRR:=jL;
CMoH
lRRH#M_HRxC:8=RCEb0;R
RH5VR#CHxR8<RCEb02ER0CRM
RlRRH#M_HRxC:#=RH;xC
CRRMH8RVR;
R0sCkRsMl_HM#CHx;M
C8CRo0M_C8C_8b;0E
MOF#M0N0kRMlC_ODRD#:MRH0CCos=R:R855CEb0R4-R2n/42R;RRRRRRRRRR-R-RFyRVqR)vX4n4O7RC#DDRCMC8
C80C$bR0Fk_#Lk_b0$C#RHRsNsN5$RM_klODCD#FR8IFM0RRj,I0H8ER-48MFI0jFR2VRFR8#0_oDFH
O;#MHoNsDRF_k0LRk#:kRF0k_L#$_0bRC;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFVsF_8k50RHkMb0FR0RH0s-N#002C#
o#HMRNDs0Fk_RCM:0R#8F_Do_HOP0COFMs5kOl_C#DDRI8FMR0FjR2;RRRRR-R-RNCML#DCRsVFRH0s-N#00
C##MHoNIDRF_k0LRk#:kRF0k_L#$_0bRC;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFVIF_8k50RHkMb0FR0RH0s-N#002C#
o#HMRNDI0Fk_RCM:0R#8F_Do_HOP0COFMs5kOl_C#DDRI8FMR0FjR2;RRRRR-R-RNCML#DCRsVFRH0s-N#00
C##MHoNIDRsC0_MRR:#_08DHFoOC_POs0F5lMk_DOCD8#RF0IMF2Rj;RRRRRRRRR--I0sHCMRCNCLD#FRVsNRCOsERFFIRVqR)vCROD
D##MHoNHDRMC_soRR:#_08DHFoOC_POs0F58IH04E-RI8FMR0FjR2;RRRRRRRRRR--k8#CRR0FsHCo#s0CRh7QRH
#oDMNRksF0C_soRR:#_08DHFoOC_POs0F58IH04E-RI8FMR0FjR2;RRRRR-RR-#RkC08RFCRso0H#C)sR_z7maH
#oDMNRkIF0C_soRR:#_08DHFoOC_POs0F58IH04E-RI8FMR0FjR2;RRRRR-RR-#RkC08RFCRso0H#CWsR_z7maH
#oDMNR8sN_osCR#:R0D8_FOoH_OPC05FsNs88I0H8ER-48MFI0jFR2R;RR-RR-#RkC08RFCRso0H#C)sRq)77
o#HMRNDI_N8sRCo:0R#8F_Do_HOP0COFNs58I8sHE80-84RF0IMF2Rj;RRRR-R-RCk#8FR0RosCHC#0sqRW7
7)#MHoNDDRFsI_Ns88R#:R0D8_FOoH_OPC05FsdFR8IFM0R;j2RRRRRRRRRRRRRR--s8N8sHRL0H#RM0bkRR0F)RqvODCD#cR5R0LH#CRsJskHC
82#MHoNDDRFII_Ns88R#:R0D8_FOoH_OPC05FsdFR8IFM0R;j2RRRRRRRRRRRRRR--I8N8sHRL0H#RM0bkRR0F)RqvODCD#cR5R0LH#CRsJskHC
82Ns00H0LkC3R\s_NlF#VVCR0\:0R#soHM;L

CMoH
R
RR-R-RRQVNs88I0H8ERR<c#RN#MHoR''jRR0Fk#MkCL8RH
0#RRRRzR4R:VRHR85N8HsI8R0E=2R4RMoCC0sNCR
RRRRRRFRDIN_s8R8s<"=Rj"jjRs&RNs8_Cjo52R;
RRRRRDRRFII_Ns88RR<="jjj"RR&I_N8s5Coj
2;RRRRCRM8oCCMsCN0R;z4
RRRRRz.RH:RVNR58I8sHE80R.=R2CRoMNCs0RC
RRRRRDRRFsI_Ns88RR<=""jjRs&RNs8_C4o5RI8FMR0Fj
2;RRRRRRRRD_FII8N8s=R<Rj"j"RR&I_N8s5Co4FR8IFM0R;j2
RRRR8CMRMoCC0sNC.Rz;R
RRdRzRRR:H5VRNs88I0H8ERR=do2RCsMCN
0CRRRRRRRRD_FIs8N8s=R<R''jRs&RNs8_C.o5RI8FMR0Fj
2;RRRRRRRRD_FII8N8s=R<R''jRI&RNs8_C.o5RI8FMR0Fj
2;RRRRCRM8oCCMsCN0R;zd
RRRRRzcRH:RVNR58I8sHE80Rd>R2CRoMNCs0RC
RRRRRDRRFsI_Ns88RR<=s_N8s5CodFR8IFM0R;j2
RRRRRRRRIDF_8IN8<sR=NRI8C_soR5d8MFI0jFR2R;
RCRRMo8RCsMCNR0Cz
c;
RRRRR--Q5VR8_HMs2CoRosCHC#0sQR7h#RkHRMoB
piRRRRzR6R:VRHRH58MC_soo2RCsMCN
0CRRRRRRRRbOsFCR##5iBp,QR7hL2RCMoH
RRRRRRRRRRRRRHV5iBpR'=R4N'RMB8RpCi'P0CM2ER0CRM
RRRRRRRRRRRRRHRRMC_so=R<Rh7Q;R
RRRRRRRRRRMRC8VRH;R
RRRRRRMRC8sRbF#OC#R;
RCRRMo8RCsMCNR0Cz
6;RRRRzRnR:VRHRF5M0HR8MC_soo2RCsMCN
0CRRRRRRRRRRRRHsM_C<oR=QR7hR;
RCRRMo8RCsMCNR0Cz
n;
RRRRR--Q5VRs0Fk_osC2CRso0H#C7sRmRzakM#HoBRmpRi
RzRR(RsR:VRHR85sF_k0s2CoRMoCC0sNCR
RRRRRRsRbF#OC#)R5_pmBis,RF_k0s2CoRoLCHRM
RRRRRRRRRHRRV)R5_pmBiRR='R4'NRM8)B_mpCi'P0CM2ER0CRM
RRRRRRRRRRRRR)RR_z7ma=R<RksF0C_soR;
RRRRRRRRRCRRMH8RVR;
RRRRRCRRMb8RsCFO#
#;RRRRCRM8oCCMsCN0Rsz(;R
RRURzs:RRRRHV50MFRFs8ks0_CRo2oCCMsCN0
RRRRRRRRRRRR7)_mRza<s=RF_k0s;Co
RRRR8CMRMoCC0sNCURzs
;
RRRR-Q-RVsR5F_k0s2CoRosCHC#0smR7zkaR#oHMRpmBiR
RR(RzI:RRRRHV5FI8ks0_CRo2oCCMsCN0
RRRRRRRRFbsO#C#R_5WmiBp,FRIks0_CRo2LHCoMR
RRRRRRRRRRVRHR_5WmiBpR'=R4N'RMW8R_pmBiP'CC2M0RC0EMR
RRRRRRRRRRRRRR_RW7amzRR<=I0Fk_osC;R
RRRRRRRRRRMRC8VRH;R
RRRRRRMRC8sRbF#OC#R;
RCRRMo8RCsMCNR0Cz;(I
RRRRIzURRR:H5VRMRF0Ik8F0C_soo2RCsMCN
0CRRRRRRRRRRRRWm_7z<aR=FRIks0_C
o;RRRRCRM8oCCMsCN0RIzU;R

R-RR-VRQRN5s8_8ss2CoRosCHC#0sqR)7R7)kM#HoBRmpRi
RzRRg:RRRRHV58sN8ss_CRo2oCCMsCN0
RRRRRRRRFbsO#C#R_5)miBp,qR)727)RoLCHRM
RRRRRRRRRHRRV)R5_pmBiRR='R4'NRM8)B_mpCi'P0CM2ER0CRM
RRRRRRRRRRRRRsRRNs8_C<oR=qR)757)Ns88I0H8ER-48MFI0jFR2R;
RRRRRRRRRCRRMH8RVR;
RRRRRCRRMb8RsCFO#
#;RRRRCRM8oCCMsCN0R;zg
RRRRjz4RH:RVMR5Fs0RNs88_osC2CRoMNCs0RC
RRRRRRRRRsRRNs8_C<oR=qR)7;7)
RRRR8CMRMoCC0sNC4RzjR;
RRRRR
RRRRRR-Q-RVIR5Ns88_osC2CRso0H#CWsRq)77RHk#MBoRpRi
RzRR4R6R:VRHRN5I8_8ss2CoRMoCC0sNCR
RRRRRRsRbF#OC#BR5pRi,W7q7)L2RCMoH
RRRRRRRRRRRRRHV5iBpR'=R4N'RMB8RpCi'P0CM2ER0CRM
RRRRRRRRRRRRRIRRNs8_C<oR=qRW757)Ns88I0H8ER-48MFI0jFR2R;
RRRRRRRRRCRRMH8RVR;
RRRRRCRRMb8RsCFO#
#;RRRRCRM8oCCMsCN0R6z4;R
RR4RznRR:H5VRMRF0I8N8sC_soo2RCsMCN
0CRRRRRRRRRRRRI_N8sRCo<W=Rq)77;R
RRMRC8CRoMNCs0zCR4
n;
RRRRR--tCCMsCN0RC0ERv)qRDOCDN#RM#8RCODC0FRDo
HORRRRzR44:FRVsRRHHMMRkOl_C#DDRI8FMR0FjCRoMNCs0RC
RRRRR-RR-VRQR85N8HsI8R0E>2RcRCMC8FR0RCOsNR0CI0sHCMRCNCLDR8NMR0FkbRk0CLMND#CRCODC0FRDo
HORRRRRRRRzR4.:VRHR85N8HsI8R0E>2RcRMoCC0sNCR
RRRRRRRRRRRRRRFRskC0_M25HRR<='R4'IMECRN5s8C_so85N8HsI8-0E4FR8IFM0RRc2=2RHR#CDCjR''R;
RRRRRRRRRRRRRIRRF_k0CHM52=R<R''4RCIEMIR5Ns8_CNo58I8sHE80-84RF0IMF2RcRH=R2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0CHM52=R<RRW IMECRN5I8C_so85N8HsI8-0E4FR8IFM0RRc2=2RHR#CDCjR''R;
RRRRRCRRMo8RCsMCNR0Cz;4.
RRRRRRRRR--Q5VRNs88I0H8E=R<RRc2MIFRsCH0RNCMLRDCFFsRkk0b0MRCNCLDRD#CCRO0DHFoOCRMC88C
RRRRRRRRdz4RH:RVNR58I8sHE80RR<=co2RCsMCN
0CRRRRRRRRRRRRRRRRs0Fk_5CMH<2R=4R''R;
RRRRRRRRRRRRRIRRF_k0CHM52=R<R''4;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R R;
RRRRRRRRRCRRMo8RCsMCNR0Cz;4d
RRRRR--tsMCNR0C0REC)RqvODCD#MRN8sR0H0-#N#0C
RRRRRRRRcz4RV:RF[sRRRHM58IH0-ERRR428MFI0jFRRMoCC0sNCR
RRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqz)vRR:DCNLD#RHR7"1a&"RR0HMCsoC'NHloIC5HE802RR&"R7"&MRH0CCosl'HN5oCHn*42RR&"RW"&MRH0CCosl'HN5oC[&2RR"" RH&RMo0CCHs'lCNo50oC_8CM_b8C05E5H2+4*,4nRb8C02E2R"&RX&"RR0HMCsoC'NHlo[C5+;42
RRRRRRRRRRRRoLCHRM
RRRRRRRRRzRR):qvRv)q44nX7RR
RRRRRRRRRRRRRbRRFRs0lRNb5=7R>MRH_osC5,[2RRqj=D>RFII_Ns885,j2RRq4=D>RFII_Ns885,42RRq.=D>RFII_Ns885,.2
RRRRRRRRRRRRRRRRRRRRRRRRqRRd>R=RIDF_8IN8ds527,Ruj)qRR=>D_FIs8N8s25j,uR7)Rq4=D>RFsI_Ns885,42RR
RRRRRRRRRRRRRRRRRRRRRRRRR7qu).>R=RIDF_8sN8.s527,Rud)qRR=>D_FIs8N8s25d, RWRR=>I_s0CHM52
,RRRRRRRRRRRRRRRRRRRRRRRRRRBRWp=iR>pRBi7,Ru=mR>FRskL0_kH#5,,[2Rm1uRR=>I0Fk_#Lk5[H,2
2;RRRRRRRRRRRRs0Fk_osC5R[2<s=RF_k0L5k#H2,[RCIEMsR5F_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRIRRF_k0s5Co[<2R=FRIkL0_kH#5,R[2IMECRF5IkC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRMRC8CRoMNCs0zCR4
c;RRRRRRRRCRM8oCCMsCN0R4z4;R
RRRRRRRRRRRRRRRRRRRRRRRRRR
RRCRM8NEsOHO0C0CksRD#CC_O0s;Nl
